module top (x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, y0);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34;
  output y0;
  wire n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84;
  LUT3 #(.INIT(8'hE8)) lut_n37 (.I0(x0), .I1(x1), .I2(x2), .O(n37));
  LUT3 #(.INIT(8'hE8)) lut_n38 (.I0(x6), .I1(x7), .I2(x8), .O(n38));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n39 (.I0(x3), .I1(x4), .I2(x5), .I3(n37), .I4(n38), .O(n39));
  LUT3 #(.INIT(8'hE8)) lut_n40 (.I0(x12), .I1(x13), .I2(x14), .O(n40));
  LUT5 #(.INIT(32'hE81717E8)) lut_n41 (.I0(x3), .I1(x4), .I2(x5), .I3(n37), .I4(n38), .O(n41));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n42 (.I0(x9), .I1(x10), .I2(x11), .I3(n40), .I4(n41), .O(n42));
  LUT3 #(.INIT(8'hE8)) lut_n43 (.I0(x18), .I1(x19), .I2(x20), .O(n43));
  LUT5 #(.INIT(32'hE81717E8)) lut_n44 (.I0(x9), .I1(x10), .I2(x11), .I3(n40), .I4(n41), .O(n44));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n45 (.I0(x15), .I1(x16), .I2(x17), .I3(n43), .I4(n44), .O(n45));
  LUT3 #(.INIT(8'hE8)) lut_n46 (.I0(n39), .I1(n42), .I2(n45), .O(n46));
  LUT3 #(.INIT(8'hE8)) lut_n47 (.I0(x24), .I1(x25), .I2(x26), .O(n47));
  LUT5 #(.INIT(32'hE81717E8)) lut_n48 (.I0(x15), .I1(x16), .I2(x17), .I3(n43), .I4(n44), .O(n48));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n49 (.I0(x21), .I1(x22), .I2(x23), .I3(n47), .I4(n48), .O(n49));
  LUT3 #(.INIT(8'hE8)) lut_n50 (.I0(x27), .I1(x28), .I2(x29), .O(n50));
  LUT5 #(.INIT(32'hE81717E8)) lut_n51 (.I0(x21), .I1(x22), .I2(x23), .I3(n47), .I4(n48), .O(n51));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n52 (.I0(x30), .I1(x31), .I2(x32), .I3(n50), .I4(n51), .O(n52));
  LUT3 #(.INIT(8'h96)) lut_n53 (.I0(n39), .I1(n42), .I2(n45), .O(n53));
  LUT3 #(.INIT(8'hE8)) lut_n54 (.I0(n49), .I1(n52), .I2(n53), .O(n54));
  LUT5 #(.INIT(32'hE81717E8)) lut_n55 (.I0(x30), .I1(x31), .I2(x32), .I3(n50), .I4(n51), .O(n55));
  LUT3 #(.INIT(8'hFE)) lut_n56 (.I0(x33), .I1(x34), .I2(n55), .O(n56));
  LUT3 #(.INIT(8'h96)) lut_n57 (.I0(n49), .I1(n52), .I2(n53), .O(n57));
  LUT2 #(.INIT(4'hE)) lut_n58 (.I0(n56), .I1(n57), .O(n58));
  LUT3 #(.INIT(8'h1E)) lut_n59 (.I0(x33), .I1(x34), .I2(n55), .O(n59));
  LUT2 #(.INIT(4'h6)) lut_n60 (.I0(n56), .I1(n57), .O(n60));
  LUT3 #(.INIT(8'h96)) lut_n61 (.I0(x0), .I1(x1), .I2(x2), .O(n61));
  LUT3 #(.INIT(8'h96)) lut_n62 (.I0(x6), .I1(x7), .I2(x8), .O(n62));
  LUT5 #(.INIT(32'hFF969600)) lut_n63 (.I0(x3), .I1(x4), .I2(x5), .I3(n61), .I4(n62), .O(n63));
  LUT3 #(.INIT(8'h96)) lut_n64 (.I0(x12), .I1(x13), .I2(x14), .O(n64));
  LUT5 #(.INIT(32'h96696996)) lut_n65 (.I0(x3), .I1(x4), .I2(x5), .I3(n61), .I4(n62), .O(n65));
  LUT5 #(.INIT(32'hFF969600)) lut_n66 (.I0(x9), .I1(x10), .I2(x11), .I3(n64), .I4(n65), .O(n66));
  LUT3 #(.INIT(8'hE8)) lut_n67 (.I0(n59), .I1(n63), .I2(n66), .O(n67));
  LUT3 #(.INIT(8'h96)) lut_n68 (.I0(n46), .I1(n54), .I2(n58), .O(n68));
  LUT4 #(.INIT(16'h7100)) lut_n69 (.I0(n59), .I1(n60), .I2(n67), .I3(n68), .O(n69));
  LUT3 #(.INIT(8'h96)) lut_n70 (.I0(x18), .I1(x19), .I2(x20), .O(n70));
  LUT5 #(.INIT(32'h96696996)) lut_n71 (.I0(x9), .I1(x10), .I2(x11), .I3(n64), .I4(n65), .O(n71));
  LUT5 #(.INIT(32'hFF969600)) lut_n72 (.I0(x15), .I1(x16), .I2(x17), .I3(n70), .I4(n71), .O(n72));
  LUT3 #(.INIT(8'h96)) lut_n73 (.I0(x24), .I1(x25), .I2(x26), .O(n73));
  LUT5 #(.INIT(32'h96696996)) lut_n74 (.I0(x15), .I1(x16), .I2(x17), .I3(n70), .I4(n71), .O(n74));
  LUT5 #(.INIT(32'hFF969600)) lut_n75 (.I0(x21), .I1(x22), .I2(x23), .I3(n73), .I4(n74), .O(n75));
  LUT3 #(.INIT(8'h96)) lut_n76 (.I0(n59), .I1(n63), .I2(n66), .O(n76));
  LUT3 #(.INIT(8'hE8)) lut_n77 (.I0(n72), .I1(n75), .I2(n76), .O(n77));
  LUT3 #(.INIT(8'h96)) lut_n78 (.I0(x30), .I1(x31), .I2(x32), .O(n78));
  LUT3 #(.INIT(8'h96)) lut_n79 (.I0(x27), .I1(x28), .I2(x29), .O(n79));
  LUT5 #(.INIT(32'h96696996)) lut_n80 (.I0(x21), .I1(x22), .I2(x23), .I3(n73), .I4(n74), .O(n80));
  LUT3 #(.INIT(8'h96)) lut_n81 (.I0(n72), .I1(n75), .I2(n76), .O(n81));
  LUT6 #(.INIT(64'hFFFFFFF9F9909000)) lut_n82 (.I0(x33), .I1(x34), .I2(n78), .I3(n79), .I4(n80), .I5(n81), .O(n82));
  LUT6 #(.INIT(64'h9EF78E718E718610)) lut_n83 (.I0(n59), .I1(n60), .I2(n67), .I3(n68), .I4(n77), .I5(n82), .O(n83));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n84 (.I0(n46), .I1(n54), .I2(n58), .I3(n69), .I4(n83), .O(n84));
  assign y0 = n84;
endmodule
