module top (x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, y0);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20;
  output y0;
  wire n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45;
  LUT3 #(.INIT(8'hE8)) lut_n23 (.I0(x0), .I1(x1), .I2(x2), .O(n23));
  LUT3 #(.INIT(8'hE8)) lut_n24 (.I0(x6), .I1(x7), .I2(x8), .O(n24));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n25 (.I0(x3), .I1(x4), .I2(x5), .I3(n23), .I4(n24), .O(n25));
  LUT3 #(.INIT(8'hE8)) lut_n26 (.I0(x12), .I1(x13), .I2(x14), .O(n26));
  LUT5 #(.INIT(32'hE81717E8)) lut_n27 (.I0(x3), .I1(x4), .I2(x5), .I3(n23), .I4(n24), .O(n27));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n28 (.I0(x9), .I1(x10), .I2(x11), .I3(n26), .I4(n27), .O(n28));
  LUT3 #(.INIT(8'hE8)) lut_n29 (.I0(x18), .I1(x19), .I2(x20), .O(n29));
  LUT5 #(.INIT(32'hE81717E8)) lut_n30 (.I0(x9), .I1(x10), .I2(x11), .I3(n26), .I4(n27), .O(n30));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n31 (.I0(x15), .I1(x16), .I2(x17), .I3(n29), .I4(n30), .O(n31));
  LUT3 #(.INIT(8'h96)) lut_n32 (.I0(x0), .I1(x1), .I2(x2), .O(n32));
  LUT3 #(.INIT(8'h96)) lut_n33 (.I0(x6), .I1(x7), .I2(x8), .O(n33));
  LUT5 #(.INIT(32'hFF969600)) lut_n34 (.I0(x3), .I1(x4), .I2(x5), .I3(n32), .I4(n33), .O(n34));
  LUT5 #(.INIT(32'hE81717E8)) lut_n35 (.I0(x15), .I1(x16), .I2(x17), .I3(n29), .I4(n30), .O(n35));
  LUT3 #(.INIT(8'h96)) lut_n36 (.I0(n25), .I1(n28), .I2(n31), .O(n36));
  LUT3 #(.INIT(8'h96)) lut_n37 (.I0(x12), .I1(x13), .I2(x14), .O(n37));
  LUT5 #(.INIT(32'h96696996)) lut_n38 (.I0(x3), .I1(x4), .I2(x5), .I3(n32), .I4(n33), .O(n38));
  LUT5 #(.INIT(32'hFF969600)) lut_n39 (.I0(x9), .I1(x10), .I2(x11), .I3(n37), .I4(n38), .O(n39));
  LUT3 #(.INIT(8'h96)) lut_n40 (.I0(x15), .I1(x16), .I2(x17), .O(n40));
  LUT5 #(.INIT(32'h96696996)) lut_n41 (.I0(x9), .I1(x10), .I2(x11), .I3(n37), .I4(n38), .O(n41));
  LUT5 #(.INIT(32'hFF969600)) lut_n42 (.I0(x18), .I1(x19), .I2(x20), .I3(n40), .I4(n41), .O(n42));
  LUT5 #(.INIT(32'h96696996)) lut_n43 (.I0(x18), .I1(x19), .I2(x20), .I3(n40), .I4(n41), .O(n43));
  LUT6 #(.INIT(64'hE787870687060600)) lut_n44 (.I0(n34), .I1(n35), .I2(n36), .I3(n39), .I4(n42), .I5(n43), .O(n44));
  LUT6 #(.INIT(64'hFFFEFEFEE8808080)) lut_n45 (.I0(n25), .I1(n28), .I2(n31), .I3(n34), .I4(n35), .I5(n44), .O(n45));
  assign y0 = n45;
endmodule
