module top (x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, y0);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22;
  output y0;
  wire n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53;
  LUT3 #(.INIT(8'hE8)) lut_n25 (.I0(x0), .I1(x1), .I2(x2), .O(n25));
  LUT3 #(.INIT(8'hE8)) lut_n26 (.I0(x6), .I1(x7), .I2(x8), .O(n26));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n27 (.I0(x3), .I1(x4), .I2(x5), .I3(n25), .I4(n26), .O(n27));
  LUT3 #(.INIT(8'hE8)) lut_n28 (.I0(x12), .I1(x13), .I2(x14), .O(n28));
  LUT5 #(.INIT(32'hE81717E8)) lut_n29 (.I0(x3), .I1(x4), .I2(x5), .I3(n25), .I4(n26), .O(n29));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n30 (.I0(x9), .I1(x10), .I2(x11), .I3(n28), .I4(n29), .O(n30));
  LUT3 #(.INIT(8'hE8)) lut_n31 (.I0(x18), .I1(x19), .I2(x20), .O(n31));
  LUT5 #(.INIT(32'hE81717E8)) lut_n32 (.I0(x9), .I1(x10), .I2(x11), .I3(n28), .I4(n29), .O(n32));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n33 (.I0(x15), .I1(x16), .I2(x17), .I3(n31), .I4(n32), .O(n33));
  LUT3 #(.INIT(8'hE8)) lut_n34 (.I0(n27), .I1(n30), .I2(n33), .O(n34));
  LUT5 #(.INIT(32'hE81717E8)) lut_n35 (.I0(x15), .I1(x16), .I2(x17), .I3(n31), .I4(n32), .O(n35));
  LUT3 #(.INIT(8'hFE)) lut_n36 (.I0(x21), .I1(x22), .I2(n35), .O(n36));
  LUT3 #(.INIT(8'h96)) lut_n37 (.I0(x0), .I1(x1), .I2(x2), .O(n37));
  LUT3 #(.INIT(8'h96)) lut_n38 (.I0(x6), .I1(x7), .I2(x8), .O(n38));
  LUT5 #(.INIT(32'hFF969600)) lut_n39 (.I0(x3), .I1(x4), .I2(x5), .I3(n37), .I4(n38), .O(n39));
  LUT3 #(.INIT(8'h1E)) lut_n40 (.I0(x21), .I1(x22), .I2(n35), .O(n40));
  LUT2 #(.INIT(4'h2)) lut_n41 (.I0(n39), .I1(n40), .O(n41));
  LUT3 #(.INIT(8'h96)) lut_n42 (.I0(n27), .I1(n30), .I2(n33), .O(n42));
  LUT3 #(.INIT(8'h96)) lut_n43 (.I0(x12), .I1(x13), .I2(x14), .O(n43));
  LUT5 #(.INIT(32'h96696996)) lut_n44 (.I0(x3), .I1(x4), .I2(x5), .I3(n37), .I4(n38), .O(n44));
  LUT5 #(.INIT(32'hFF969600)) lut_n45 (.I0(x9), .I1(x10), .I2(x11), .I3(n43), .I4(n44), .O(n45));
  LUT3 #(.INIT(8'h96)) lut_n46 (.I0(x15), .I1(x16), .I2(x17), .O(n46));
  LUT3 #(.INIT(8'h96)) lut_n47 (.I0(x18), .I1(x19), .I2(x20), .O(n47));
  LUT5 #(.INIT(32'h96696996)) lut_n48 (.I0(x9), .I1(x10), .I2(x11), .I3(n43), .I4(n44), .O(n48));
  LUT2 #(.INIT(4'h6)) lut_n49 (.I0(n39), .I1(n40), .O(n49));
  LUT5 #(.INIT(32'hA880FEEA)) lut_n50 (.I0(n45), .I1(n46), .I2(n47), .I3(n48), .I4(n49), .O(n50));
  LUT2 #(.INIT(4'h6)) lut_n51 (.I0(x21), .I1(x22), .O(n51));
  LUT6 #(.INIT(64'hBDD77EEBA995566A)) lut_n52 (.I0(n45), .I1(n46), .I2(n47), .I3(n48), .I4(n49), .I5(n51), .O(n52));
  LUT6 #(.INIT(64'hEAA8A880FEEAEAA8)) lut_n53 (.I0(n34), .I1(n36), .I2(n41), .I3(n42), .I4(n50), .I5(n52), .O(n53));
  assign y0 = n53;
endmodule
