module top (x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255, x256, x257, x258, x259, x260, x261, x262, x263, x264, x265, x266, x267, x268, x269, x270, x271, x272, x273, x274, x275, x276, x277, x278, x279, x280, x281, x282, x283, x284, x285, x286, x287, x288, x289, x290, x291, x292, x293, x294, x295, x296, x297, x298, x299, x300, x301, x302, x303, x304, x305, x306, x307, x308, x309, x310, x311, x312, x313, x314, x315, x316, x317, x318, x319, x320, x321, x322, x323, x324, x325, x326, x327, x328, x329, x330, x331, x332, x333, x334, x335, x336, x337, x338, x339, x340, x341, x342, x343, x344, x345, x346, x347, x348, x349, x350, x351, x352, x353, x354, x355, x356, x357, x358, x359, x360, x361, x362, x363, x364, x365, x366, x367, x368, x369, x370, x371, x372, x373, x374, x375, x376, x377, x378, x379, x380, x381, x382, x383, x384, x385, x386, x387, x388, x389, x390, x391, x392, x393, x394, x395, x396, x397, x398, x399, x400, x401, x402, x403, x404, x405, x406, x407, x408, x409, x410, x411, x412, x413, x414, x415, x416, x417, x418, x419, x420, x421, x422, x423, x424, x425, x426, x427, x428, x429, x430, x431, x432, x433, x434, x435, x436, x437, x438, x439, x440, x441, x442, x443, x444, x445, x446, x447, x448, x449, x450, x451, x452, x453, x454, x455, x456, x457, x458, x459, x460, x461, x462, x463, x464, x465, x466, x467, x468, x469, x470, x471, x472, x473, x474, x475, x476, x477, x478, x479, x480, x481, x482, x483, x484, x485, x486, x487, x488, x489, x490, x491, x492, x493, x494, x495, x496, x497, x498, x499, x500, x501, x502, x503, x504, x505, x506, x507, x508, x509, x510, x511, x512, x513, x514, x515, x516, x517, x518, x519, x520, x521, x522, x523, x524, x525, x526, x527, x528, x529, x530, x531, x532, x533, x534, x535, x536, x537, x538, x539, x540, x541, x542, x543, x544, x545, x546, x547, x548, x549, x550, x551, x552, x553, x554, x555, x556, x557, x558, x559, x560, x561, x562, x563, x564, x565, x566, x567, x568, x569, x570, x571, x572, x573, x574, x575, x576, x577, x578, x579, x580, x581, x582, x583, x584, x585, x586, x587, x588, x589, x590, x591, x592, x593, x594, x595, x596, x597, x598, x599, x600, x601, x602, x603, x604, x605, x606, x607, x608, x609, x610, x611, x612, x613, x614, x615, x616, x617, x618, x619, x620, x621, x622, x623, x624, x625, x626, x627, x628, x629, x630, x631, x632, x633, x634, x635, x636, x637, x638, x639, x640, x641, x642, x643, x644, x645, x646, x647, x648, x649, x650, x651, x652, x653, x654, x655, x656, x657, x658, x659, x660, x661, x662, x663, x664, x665, x666, x667, x668, x669, x670, x671, x672, x673, x674, x675, x676, x677, x678, x679, x680, x681, x682, x683, x684, x685, x686, x687, x688, x689, x690, x691, x692, x693, x694, x695, x696, x697, x698, x699, x700, x701, x702, x703, x704, x705, x706, x707, x708, x709, x710, x711, x712, x713, x714, x715, x716, x717, x718, x719, x720, x721, x722, x723, x724, x725, x726, x727, x728, x729, x730, x731, x732, x733, x734, x735, x736, x737, x738, x739, x740, x741, x742, x743, x744, x745, x746, x747, x748, x749, x750, x751, x752, x753, x754, x755, x756, x757, x758, x759, x760, x761, x762, x763, x764, x765, x766, x767, x768, x769, x770, x771, x772, x773, x774, x775, x776, x777, x778, x779, x780, x781, x782, x783, x784, x785, x786, x787, x788, x789, x790, x791, x792, x793, x794, x795, x796, x797, x798, x799, x800, x801, x802, x803, x804, x805, x806, x807, x808, x809, x810, x811, x812, x813, x814, x815, x816, x817, x818, x819, x820, x821, x822, x823, x824, x825, x826, x827, x828, x829, x830, x831, x832, x833, x834, x835, x836, x837, x838, x839, x840, x841, x842, x843, x844, x845, x846, x847, x848, x849, x850, x851, x852, x853, x854, x855, x856, x857, x858, x859, x860, x861, x862, x863, x864, x865, x866, x867, x868, x869, x870, x871, x872, x873, x874, x875, x876, x877, x878, x879, x880, x881, x882, x883, x884, x885, x886, x887, x888, x889, x890, x891, x892, x893, x894, x895, x896, x897, x898, x899, x900, x901, x902, x903, x904, x905, x906, x907, x908, x909, x910, x911, x912, x913, x914, x915, x916, x917, x918, x919, x920, x921, x922, x923, x924, x925, x926, x927, x928, x929, x930, x931, x932, x933, x934, x935, x936, x937, x938, x939, x940, x941, x942, x943, x944, x945, x946, x947, x948, x949, x950, x951, x952, x953, x954, x955, x956, x957, x958, x959, x960, x961, x962, x963, x964, x965, x966, x967, x968, x969, x970, x971, x972, x973, x974, x975, x976, x977, x978, x979, x980, x981, x982, x983, x984, x985, x986, x987, x988, x989, x990, x991, x992, x993, x994, x995, x996, x997, x998, x999, x1000, x1001, x1002, x1003, x1004, x1005, x1006, x1007, x1008, x1009, x1010, x1011, x1012, x1013, x1014, x1015, x1016, x1017, x1018, x1019, x1020, x1021, x1022, x1023, x1024, x1025, x1026, x1027, x1028, x1029, x1030, x1031, x1032, x1033, x1034, x1035, x1036, x1037, x1038, x1039, x1040, x1041, x1042, x1043, x1044, x1045, x1046, x1047, x1048, x1049, x1050, x1051, x1052, x1053, x1054, x1055, x1056, x1057, x1058, x1059, x1060, x1061, x1062, x1063, x1064, x1065, x1066, x1067, x1068, x1069, x1070, x1071, x1072, x1073, x1074, x1075, x1076, x1077, x1078, x1079, x1080, x1081, x1082, x1083, x1084, x1085, x1086, x1087, x1088, x1089, x1090, x1091, x1092, x1093, x1094, x1095, x1096, x1097, x1098, x1099, x1100, x1101, x1102, x1103, x1104, x1105, x1106, x1107, x1108, x1109, x1110, x1111, x1112, x1113, x1114, x1115, x1116, x1117, x1118, x1119, x1120, x1121, x1122, x1123, x1124, x1125, x1126, x1127, x1128, x1129, x1130, x1131, x1132, x1133, x1134, x1135, x1136, x1137, x1138, x1139, x1140, x1141, x1142, x1143, x1144, x1145, x1146, x1147, x1148, x1149, x1150, x1151, x1152, x1153, x1154, x1155, x1156, x1157, x1158, x1159, x1160, x1161, x1162, x1163, x1164, x1165, x1166, x1167, x1168, x1169, x1170, x1171, x1172, x1173, x1174, x1175, x1176, x1177, x1178, x1179, x1180, x1181, x1182, x1183, x1184, x1185, x1186, x1187, x1188, x1189, x1190, x1191, x1192, x1193, x1194, x1195, x1196, x1197, x1198, x1199, x1200, x1201, x1202, x1203, x1204, x1205, x1206, x1207, x1208, x1209, x1210, x1211, x1212, x1213, x1214, x1215, x1216, x1217, x1218, x1219, x1220, x1221, x1222, x1223, x1224, x1225, x1226, x1227, x1228, x1229, x1230, x1231, x1232, x1233, x1234, x1235, x1236, x1237, x1238, x1239, x1240, x1241, x1242, x1243, x1244, x1245, x1246, x1247, x1248, x1249, x1250, x1251, x1252, x1253, x1254, x1255, x1256, x1257, x1258, x1259, x1260, x1261, x1262, x1263, x1264, x1265, x1266, x1267, x1268, x1269, x1270, x1271, x1272, x1273, x1274, x1275, x1276, x1277, x1278, x1279, x1280, x1281, x1282, x1283, x1284, x1285, x1286, x1287, x1288, x1289, x1290, x1291, x1292, x1293, x1294, x1295, x1296, x1297, x1298, x1299, x1300, x1301, x1302, x1303, x1304, x1305, x1306, x1307, x1308, x1309, x1310, x1311, x1312, x1313, x1314, x1315, x1316, x1317, x1318, x1319, x1320, x1321, x1322, x1323, x1324, x1325, x1326, x1327, x1328, x1329, x1330, x1331, x1332, x1333, x1334, x1335, x1336, x1337, x1338, x1339, x1340, x1341, x1342, x1343, x1344, x1345, x1346, x1347, x1348, x1349, x1350, x1351, x1352, x1353, x1354, x1355, x1356, x1357, x1358, x1359, x1360, x1361, x1362, x1363, x1364, x1365, x1366, x1367, x1368, x1369, x1370, x1371, x1372, x1373, x1374, x1375, x1376, x1377, x1378, x1379, x1380, x1381, x1382, x1383, x1384, x1385, x1386, x1387, x1388, x1389, x1390, x1391, x1392, x1393, x1394, x1395, x1396, x1397, x1398, x1399, x1400, x1401, x1402, x1403, x1404, x1405, x1406, x1407, x1408, x1409, x1410, x1411, x1412, x1413, x1414, x1415, x1416, x1417, x1418, x1419, x1420, x1421, x1422, x1423, x1424, x1425, x1426, x1427, x1428, x1429, x1430, x1431, x1432, x1433, x1434, x1435, x1436, x1437, x1438, x1439, x1440, x1441, x1442, x1443, x1444, x1445, x1446, x1447, x1448, x1449, x1450, x1451, x1452, x1453, x1454, x1455, x1456, x1457, x1458, x1459, x1460, x1461, x1462, x1463, x1464, x1465, x1466, x1467, x1468, x1469, x1470, x1471, x1472, x1473, x1474, x1475, x1476, x1477, x1478, x1479, x1480, x1481, x1482, x1483, x1484, x1485, x1486, x1487, x1488, x1489, x1490, x1491, x1492, x1493, x1494, x1495, x1496, x1497, x1498, x1499, x1500, x1501, x1502, x1503, x1504, x1505, x1506, x1507, x1508, x1509, x1510, x1511, x1512, x1513, x1514, x1515, x1516, x1517, x1518, x1519, x1520, x1521, x1522, x1523, x1524, x1525, x1526, x1527, x1528, x1529, x1530, x1531, x1532, x1533, x1534, x1535, x1536, x1537, x1538, x1539, x1540, x1541, x1542, x1543, x1544, x1545, x1546, x1547, x1548, x1549, x1550, x1551, x1552, x1553, x1554, x1555, x1556, x1557, x1558, x1559, x1560, x1561, x1562, x1563, x1564, x1565, x1566, x1567, x1568, x1569, x1570, x1571, x1572, x1573, x1574, x1575, x1576, x1577, x1578, x1579, x1580, x1581, x1582, x1583, x1584, x1585, x1586, x1587, x1588, x1589, x1590, x1591, x1592, x1593, x1594, x1595, x1596, x1597, x1598, x1599, x1600, x1601, x1602, x1603, x1604, x1605, x1606, x1607, x1608, x1609, x1610, x1611, x1612, x1613, x1614, x1615, x1616, x1617, x1618, x1619, x1620, x1621, x1622, x1623, x1624, x1625, x1626, x1627, x1628, x1629, x1630, x1631, x1632, x1633, x1634, x1635, x1636, x1637, x1638, x1639, x1640, x1641, x1642, x1643, x1644, x1645, x1646, x1647, x1648, x1649, x1650, x1651, x1652, x1653, x1654, x1655, x1656, x1657, x1658, x1659, x1660, x1661, x1662, x1663, x1664, x1665, x1666, x1667, x1668, x1669, x1670, x1671, x1672, x1673, x1674, x1675, x1676, x1677, x1678, x1679, x1680, x1681, x1682, x1683, x1684, x1685, x1686, x1687, x1688, x1689, x1690, x1691, x1692, x1693, x1694, x1695, x1696, x1697, x1698, x1699, x1700, x1701, x1702, x1703, x1704, x1705, x1706, x1707, x1708, x1709, x1710, x1711, x1712, x1713, x1714, x1715, x1716, x1717, x1718, x1719, x1720, x1721, x1722, x1723, x1724, x1725, x1726, x1727, x1728, x1729, x1730, x1731, x1732, x1733, x1734, x1735, x1736, x1737, x1738, x1739, x1740, x1741, x1742, x1743, x1744, x1745, x1746, x1747, x1748, x1749, x1750, x1751, x1752, x1753, x1754, x1755, x1756, x1757, x1758, x1759, x1760, x1761, x1762, x1763, x1764, x1765, x1766, x1767, x1768, x1769, x1770, x1771, x1772, x1773, x1774, x1775, x1776, x1777, x1778, x1779, x1780, x1781, x1782, x1783, x1784, x1785, x1786, x1787, x1788, x1789, x1790, x1791, x1792, x1793, x1794, x1795, x1796, x1797, x1798, x1799, x1800, x1801, x1802, x1803, x1804, x1805, x1806, x1807, x1808, x1809, x1810, x1811, x1812, x1813, x1814, x1815, x1816, x1817, x1818, x1819, x1820, x1821, x1822, x1823, x1824, x1825, x1826, x1827, x1828, x1829, x1830, x1831, x1832, x1833, x1834, x1835, x1836, x1837, x1838, x1839, x1840, x1841, x1842, x1843, x1844, x1845, x1846, x1847, x1848, x1849, x1850, x1851, x1852, x1853, x1854, x1855, x1856, x1857, x1858, x1859, x1860, x1861, x1862, x1863, x1864, x1865, x1866, x1867, x1868, x1869, x1870, x1871, x1872, x1873, x1874, x1875, x1876, x1877, x1878, x1879, x1880, x1881, x1882, x1883, x1884, x1885, x1886, x1887, x1888, x1889, x1890, x1891, x1892, x1893, x1894, x1895, x1896, x1897, x1898, x1899, x1900, x1901, x1902, x1903, x1904, x1905, x1906, x1907, x1908, x1909, x1910, x1911, x1912, x1913, x1914, x1915, x1916, x1917, x1918, x1919, x1920, x1921, x1922, x1923, x1924, x1925, x1926, x1927, x1928, x1929, x1930, x1931, x1932, x1933, x1934, x1935, x1936, x1937, x1938, x1939, x1940, x1941, x1942, x1943, x1944, x1945, x1946, x1947, x1948, x1949, x1950, x1951, x1952, x1953, x1954, x1955, x1956, x1957, x1958, x1959, x1960, x1961, x1962, x1963, x1964, x1965, x1966, x1967, x1968, x1969, x1970, x1971, x1972, x1973, x1974, x1975, x1976, x1977, x1978, x1979, x1980, x1981, x1982, x1983, x1984, x1985, x1986, x1987, x1988, x1989, x1990, x1991, x1992, x1993, x1994, x1995, x1996, x1997, x1998, x1999, x2000, x2001, x2002, x2003, x2004, x2005, x2006, x2007, x2008, x2009, x2010, x2011, x2012, x2013, x2014, x2015, x2016, x2017, x2018, x2019, x2020, x2021, x2022, x2023, x2024, x2025, x2026, x2027, x2028, x2029, x2030, x2031, x2032, x2033, x2034, x2035, x2036, x2037, x2038, x2039, x2040, x2041, x2042, x2043, x2044, x2045, x2046, x2047, x2048, x2049, x2050, x2051, x2052, x2053, x2054, x2055, x2056, x2057, x2058, x2059, x2060, x2061, x2062, x2063, x2064, x2065, x2066, x2067, x2068, x2069, x2070, x2071, x2072, x2073, x2074, x2075, x2076, x2077, x2078, x2079, x2080, x2081, x2082, x2083, x2084, x2085, x2086, x2087, x2088, x2089, x2090, x2091, x2092, x2093, x2094, x2095, x2096, x2097, x2098, x2099, x2100, x2101, x2102, x2103, x2104, x2105, x2106, x2107, x2108, x2109, x2110, x2111, x2112, x2113, x2114, x2115, x2116, x2117, x2118, x2119, x2120, x2121, x2122, x2123, x2124, x2125, x2126, x2127, x2128, x2129, x2130, x2131, x2132, x2133, x2134, x2135, x2136, x2137, x2138, x2139, x2140, x2141, x2142, x2143, x2144, x2145, x2146, x2147, x2148, x2149, x2150, x2151, x2152, x2153, x2154, x2155, x2156, x2157, x2158, x2159, x2160, x2161, x2162, x2163, x2164, x2165, x2166, x2167, x2168, x2169, x2170, x2171, x2172, x2173, x2174, x2175, x2176, x2177, x2178, x2179, x2180, x2181, x2182, x2183, x2184, x2185, x2186, x2187, x2188, x2189, x2190, x2191, x2192, x2193, x2194, x2195, x2196, x2197, x2198, x2199, x2200, x2201, x2202, x2203, x2204, x2205, x2206, x2207, x2208, x2209, x2210, x2211, x2212, x2213, x2214, x2215, x2216, x2217, x2218, x2219, x2220, x2221, x2222, x2223, x2224, x2225, x2226, x2227, x2228, x2229, x2230, x2231, x2232, x2233, x2234, x2235, x2236, x2237, x2238, x2239, x2240, x2241, x2242, x2243, x2244, x2245, x2246, x2247, x2248, x2249, x2250, x2251, x2252, x2253, x2254, x2255, x2256, x2257, x2258, x2259, x2260, x2261, x2262, x2263, x2264, x2265, x2266, x2267, x2268, x2269, x2270, x2271, x2272, x2273, x2274, x2275, x2276, x2277, x2278, x2279, x2280, x2281, x2282, x2283, x2284, x2285, x2286, x2287, x2288, x2289, x2290, x2291, x2292, x2293, x2294, x2295, x2296, x2297, x2298, x2299, x2300, x2301, x2302, x2303, x2304, x2305, x2306, x2307, x2308, x2309, x2310, x2311, x2312, x2313, x2314, x2315, x2316, x2317, x2318, x2319, x2320, x2321, x2322, x2323, x2324, x2325, x2326, x2327, x2328, x2329, x2330, x2331, x2332, x2333, x2334, x2335, x2336, x2337, x2338, x2339, x2340, x2341, x2342, x2343, x2344, x2345, x2346, x2347, x2348, x2349, x2350, x2351, x2352, x2353, x2354, x2355, x2356, x2357, x2358, x2359, x2360, x2361, x2362, x2363, x2364, x2365, x2366, x2367, x2368, x2369, x2370, x2371, x2372, x2373, x2374, x2375, x2376, x2377, x2378, x2379, x2380, x2381, x2382, x2383, x2384, x2385, x2386, x2387, x2388, x2389, x2390, x2391, x2392, x2393, x2394, x2395, x2396, x2397, x2398, x2399, x2400, x2401, x2402, x2403, x2404, x2405, x2406, x2407, x2408, x2409, x2410, x2411, x2412, x2413, x2414, x2415, x2416, x2417, x2418, x2419, x2420, x2421, x2422, x2423, x2424, x2425, x2426, x2427, x2428, x2429, x2430, x2431, x2432, x2433, x2434, x2435, x2436, x2437, x2438, x2439, x2440, x2441, x2442, x2443, x2444, x2445, x2446, x2447, x2448, x2449, x2450, x2451, x2452, x2453, x2454, x2455, x2456, x2457, x2458, x2459, x2460, x2461, x2462, x2463, x2464, x2465, x2466, x2467, x2468, x2469, x2470, x2471, x2472, x2473, x2474, x2475, x2476, x2477, x2478, x2479, x2480, x2481, x2482, x2483, x2484, x2485, x2486, x2487, x2488, x2489, x2490, x2491, x2492, x2493, x2494, x2495, x2496, x2497, x2498, x2499, x2500, x2501, x2502, x2503, x2504, x2505, x2506, x2507, x2508, x2509, x2510, x2511, x2512, x2513, x2514, x2515, x2516, x2517, x2518, x2519, x2520, x2521, x2522, x2523, x2524, x2525, x2526, x2527, x2528, x2529, x2530, x2531, x2532, x2533, x2534, x2535, x2536, x2537, x2538, x2539, x2540, x2541, x2542, x2543, x2544, x2545, x2546, x2547, x2548, x2549, x2550, x2551, x2552, x2553, x2554, x2555, x2556, x2557, x2558, x2559, x2560, x2561, x2562, x2563, x2564, x2565, x2566, x2567, x2568, x2569, x2570, x2571, x2572, x2573, x2574, x2575, x2576, x2577, x2578, x2579, x2580, x2581, x2582, x2583, x2584, x2585, x2586, x2587, x2588, x2589, x2590, x2591, x2592, x2593, x2594, x2595, x2596, x2597, x2598, x2599, x2600, x2601, x2602, x2603, x2604, x2605, x2606, x2607, x2608, x2609, x2610, x2611, x2612, x2613, x2614, x2615, x2616, x2617, x2618, x2619, x2620, x2621, x2622, x2623, x2624, x2625, x2626, x2627, x2628, x2629, x2630, x2631, x2632, x2633, x2634, x2635, x2636, x2637, x2638, x2639, x2640, x2641, x2642, x2643, x2644, x2645, x2646, x2647, x2648, x2649, x2650, x2651, x2652, x2653, x2654, x2655, x2656, x2657, x2658, x2659, x2660, x2661, x2662, x2663, x2664, x2665, x2666, x2667, x2668, x2669, x2670, x2671, x2672, x2673, x2674, x2675, x2676, x2677, x2678, x2679, x2680, x2681, x2682, x2683, x2684, x2685, x2686, x2687, x2688, x2689, x2690, x2691, x2692, x2693, x2694, x2695, x2696, x2697, x2698, x2699, x2700, x2701, x2702, x2703, x2704, x2705, x2706, x2707, x2708, x2709, x2710, x2711, x2712, x2713, x2714, x2715, x2716, x2717, x2718, x2719, x2720, x2721, x2722, x2723, x2724, x2725, x2726, x2727, x2728, x2729, x2730, x2731, x2732, x2733, x2734, x2735, x2736, x2737, x2738, x2739, x2740, x2741, x2742, x2743, x2744, x2745, x2746, x2747, x2748, x2749, x2750, x2751, x2752, x2753, x2754, x2755, x2756, x2757, x2758, x2759, x2760, x2761, x2762, x2763, x2764, x2765, x2766, x2767, x2768, x2769, x2770, x2771, x2772, x2773, x2774, x2775, x2776, x2777, x2778, x2779, x2780, x2781, x2782, x2783, x2784, x2785, x2786, x2787, x2788, x2789, x2790, x2791, x2792, x2793, x2794, x2795, x2796, x2797, x2798, x2799, x2800, x2801, x2802, x2803, x2804, x2805, x2806, x2807, x2808, x2809, x2810, x2811, x2812, x2813, x2814, x2815, x2816, x2817, x2818, x2819, x2820, x2821, x2822, x2823, x2824, x2825, x2826, x2827, x2828, x2829, x2830, x2831, x2832, x2833, x2834, x2835, x2836, x2837, x2838, x2839, x2840, x2841, x2842, x2843, x2844, x2845, x2846, x2847, x2848, x2849, x2850, x2851, x2852, x2853, x2854, x2855, x2856, x2857, x2858, x2859, x2860, x2861, x2862, x2863, x2864, x2865, x2866, x2867, x2868, x2869, x2870, x2871, x2872, x2873, x2874, x2875, x2876, x2877, x2878, x2879, x2880, x2881, x2882, x2883, x2884, x2885, x2886, x2887, x2888, x2889, x2890, x2891, x2892, x2893, x2894, x2895, x2896, x2897, x2898, x2899, x2900, x2901, x2902, x2903, x2904, x2905, x2906, x2907, x2908, x2909, x2910, x2911, x2912, x2913, x2914, x2915, x2916, x2917, x2918, x2919, x2920, x2921, x2922, x2923, x2924, x2925, x2926, x2927, x2928, x2929, x2930, x2931, x2932, x2933, x2934, x2935, x2936, x2937, x2938, x2939, x2940, x2941, x2942, x2943, x2944, x2945, x2946, x2947, x2948, x2949, x2950, x2951, x2952, x2953, x2954, x2955, x2956, x2957, x2958, x2959, x2960, x2961, x2962, x2963, x2964, x2965, x2966, x2967, x2968, x2969, x2970, x2971, x2972, x2973, x2974, x2975, x2976, x2977, x2978, x2979, x2980, x2981, x2982, x2983, x2984, x2985, x2986, x2987, x2988, x2989, x2990, x2991, x2992, x2993, x2994, x2995, x2996, x2997, x2998, x2999, x3000, y0);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255, x256, x257, x258, x259, x260, x261, x262, x263, x264, x265, x266, x267, x268, x269, x270, x271, x272, x273, x274, x275, x276, x277, x278, x279, x280, x281, x282, x283, x284, x285, x286, x287, x288, x289, x290, x291, x292, x293, x294, x295, x296, x297, x298, x299, x300, x301, x302, x303, x304, x305, x306, x307, x308, x309, x310, x311, x312, x313, x314, x315, x316, x317, x318, x319, x320, x321, x322, x323, x324, x325, x326, x327, x328, x329, x330, x331, x332, x333, x334, x335, x336, x337, x338, x339, x340, x341, x342, x343, x344, x345, x346, x347, x348, x349, x350, x351, x352, x353, x354, x355, x356, x357, x358, x359, x360, x361, x362, x363, x364, x365, x366, x367, x368, x369, x370, x371, x372, x373, x374, x375, x376, x377, x378, x379, x380, x381, x382, x383, x384, x385, x386, x387, x388, x389, x390, x391, x392, x393, x394, x395, x396, x397, x398, x399, x400, x401, x402, x403, x404, x405, x406, x407, x408, x409, x410, x411, x412, x413, x414, x415, x416, x417, x418, x419, x420, x421, x422, x423, x424, x425, x426, x427, x428, x429, x430, x431, x432, x433, x434, x435, x436, x437, x438, x439, x440, x441, x442, x443, x444, x445, x446, x447, x448, x449, x450, x451, x452, x453, x454, x455, x456, x457, x458, x459, x460, x461, x462, x463, x464, x465, x466, x467, x468, x469, x470, x471, x472, x473, x474, x475, x476, x477, x478, x479, x480, x481, x482, x483, x484, x485, x486, x487, x488, x489, x490, x491, x492, x493, x494, x495, x496, x497, x498, x499, x500, x501, x502, x503, x504, x505, x506, x507, x508, x509, x510, x511, x512, x513, x514, x515, x516, x517, x518, x519, x520, x521, x522, x523, x524, x525, x526, x527, x528, x529, x530, x531, x532, x533, x534, x535, x536, x537, x538, x539, x540, x541, x542, x543, x544, x545, x546, x547, x548, x549, x550, x551, x552, x553, x554, x555, x556, x557, x558, x559, x560, x561, x562, x563, x564, x565, x566, x567, x568, x569, x570, x571, x572, x573, x574, x575, x576, x577, x578, x579, x580, x581, x582, x583, x584, x585, x586, x587, x588, x589, x590, x591, x592, x593, x594, x595, x596, x597, x598, x599, x600, x601, x602, x603, x604, x605, x606, x607, x608, x609, x610, x611, x612, x613, x614, x615, x616, x617, x618, x619, x620, x621, x622, x623, x624, x625, x626, x627, x628, x629, x630, x631, x632, x633, x634, x635, x636, x637, x638, x639, x640, x641, x642, x643, x644, x645, x646, x647, x648, x649, x650, x651, x652, x653, x654, x655, x656, x657, x658, x659, x660, x661, x662, x663, x664, x665, x666, x667, x668, x669, x670, x671, x672, x673, x674, x675, x676, x677, x678, x679, x680, x681, x682, x683, x684, x685, x686, x687, x688, x689, x690, x691, x692, x693, x694, x695, x696, x697, x698, x699, x700, x701, x702, x703, x704, x705, x706, x707, x708, x709, x710, x711, x712, x713, x714, x715, x716, x717, x718, x719, x720, x721, x722, x723, x724, x725, x726, x727, x728, x729, x730, x731, x732, x733, x734, x735, x736, x737, x738, x739, x740, x741, x742, x743, x744, x745, x746, x747, x748, x749, x750, x751, x752, x753, x754, x755, x756, x757, x758, x759, x760, x761, x762, x763, x764, x765, x766, x767, x768, x769, x770, x771, x772, x773, x774, x775, x776, x777, x778, x779, x780, x781, x782, x783, x784, x785, x786, x787, x788, x789, x790, x791, x792, x793, x794, x795, x796, x797, x798, x799, x800, x801, x802, x803, x804, x805, x806, x807, x808, x809, x810, x811, x812, x813, x814, x815, x816, x817, x818, x819, x820, x821, x822, x823, x824, x825, x826, x827, x828, x829, x830, x831, x832, x833, x834, x835, x836, x837, x838, x839, x840, x841, x842, x843, x844, x845, x846, x847, x848, x849, x850, x851, x852, x853, x854, x855, x856, x857, x858, x859, x860, x861, x862, x863, x864, x865, x866, x867, x868, x869, x870, x871, x872, x873, x874, x875, x876, x877, x878, x879, x880, x881, x882, x883, x884, x885, x886, x887, x888, x889, x890, x891, x892, x893, x894, x895, x896, x897, x898, x899, x900, x901, x902, x903, x904, x905, x906, x907, x908, x909, x910, x911, x912, x913, x914, x915, x916, x917, x918, x919, x920, x921, x922, x923, x924, x925, x926, x927, x928, x929, x930, x931, x932, x933, x934, x935, x936, x937, x938, x939, x940, x941, x942, x943, x944, x945, x946, x947, x948, x949, x950, x951, x952, x953, x954, x955, x956, x957, x958, x959, x960, x961, x962, x963, x964, x965, x966, x967, x968, x969, x970, x971, x972, x973, x974, x975, x976, x977, x978, x979, x980, x981, x982, x983, x984, x985, x986, x987, x988, x989, x990, x991, x992, x993, x994, x995, x996, x997, x998, x999, x1000, x1001, x1002, x1003, x1004, x1005, x1006, x1007, x1008, x1009, x1010, x1011, x1012, x1013, x1014, x1015, x1016, x1017, x1018, x1019, x1020, x1021, x1022, x1023, x1024, x1025, x1026, x1027, x1028, x1029, x1030, x1031, x1032, x1033, x1034, x1035, x1036, x1037, x1038, x1039, x1040, x1041, x1042, x1043, x1044, x1045, x1046, x1047, x1048, x1049, x1050, x1051, x1052, x1053, x1054, x1055, x1056, x1057, x1058, x1059, x1060, x1061, x1062, x1063, x1064, x1065, x1066, x1067, x1068, x1069, x1070, x1071, x1072, x1073, x1074, x1075, x1076, x1077, x1078, x1079, x1080, x1081, x1082, x1083, x1084, x1085, x1086, x1087, x1088, x1089, x1090, x1091, x1092, x1093, x1094, x1095, x1096, x1097, x1098, x1099, x1100, x1101, x1102, x1103, x1104, x1105, x1106, x1107, x1108, x1109, x1110, x1111, x1112, x1113, x1114, x1115, x1116, x1117, x1118, x1119, x1120, x1121, x1122, x1123, x1124, x1125, x1126, x1127, x1128, x1129, x1130, x1131, x1132, x1133, x1134, x1135, x1136, x1137, x1138, x1139, x1140, x1141, x1142, x1143, x1144, x1145, x1146, x1147, x1148, x1149, x1150, x1151, x1152, x1153, x1154, x1155, x1156, x1157, x1158, x1159, x1160, x1161, x1162, x1163, x1164, x1165, x1166, x1167, x1168, x1169, x1170, x1171, x1172, x1173, x1174, x1175, x1176, x1177, x1178, x1179, x1180, x1181, x1182, x1183, x1184, x1185, x1186, x1187, x1188, x1189, x1190, x1191, x1192, x1193, x1194, x1195, x1196, x1197, x1198, x1199, x1200, x1201, x1202, x1203, x1204, x1205, x1206, x1207, x1208, x1209, x1210, x1211, x1212, x1213, x1214, x1215, x1216, x1217, x1218, x1219, x1220, x1221, x1222, x1223, x1224, x1225, x1226, x1227, x1228, x1229, x1230, x1231, x1232, x1233, x1234, x1235, x1236, x1237, x1238, x1239, x1240, x1241, x1242, x1243, x1244, x1245, x1246, x1247, x1248, x1249, x1250, x1251, x1252, x1253, x1254, x1255, x1256, x1257, x1258, x1259, x1260, x1261, x1262, x1263, x1264, x1265, x1266, x1267, x1268, x1269, x1270, x1271, x1272, x1273, x1274, x1275, x1276, x1277, x1278, x1279, x1280, x1281, x1282, x1283, x1284, x1285, x1286, x1287, x1288, x1289, x1290, x1291, x1292, x1293, x1294, x1295, x1296, x1297, x1298, x1299, x1300, x1301, x1302, x1303, x1304, x1305, x1306, x1307, x1308, x1309, x1310, x1311, x1312, x1313, x1314, x1315, x1316, x1317, x1318, x1319, x1320, x1321, x1322, x1323, x1324, x1325, x1326, x1327, x1328, x1329, x1330, x1331, x1332, x1333, x1334, x1335, x1336, x1337, x1338, x1339, x1340, x1341, x1342, x1343, x1344, x1345, x1346, x1347, x1348, x1349, x1350, x1351, x1352, x1353, x1354, x1355, x1356, x1357, x1358, x1359, x1360, x1361, x1362, x1363, x1364, x1365, x1366, x1367, x1368, x1369, x1370, x1371, x1372, x1373, x1374, x1375, x1376, x1377, x1378, x1379, x1380, x1381, x1382, x1383, x1384, x1385, x1386, x1387, x1388, x1389, x1390, x1391, x1392, x1393, x1394, x1395, x1396, x1397, x1398, x1399, x1400, x1401, x1402, x1403, x1404, x1405, x1406, x1407, x1408, x1409, x1410, x1411, x1412, x1413, x1414, x1415, x1416, x1417, x1418, x1419, x1420, x1421, x1422, x1423, x1424, x1425, x1426, x1427, x1428, x1429, x1430, x1431, x1432, x1433, x1434, x1435, x1436, x1437, x1438, x1439, x1440, x1441, x1442, x1443, x1444, x1445, x1446, x1447, x1448, x1449, x1450, x1451, x1452, x1453, x1454, x1455, x1456, x1457, x1458, x1459, x1460, x1461, x1462, x1463, x1464, x1465, x1466, x1467, x1468, x1469, x1470, x1471, x1472, x1473, x1474, x1475, x1476, x1477, x1478, x1479, x1480, x1481, x1482, x1483, x1484, x1485, x1486, x1487, x1488, x1489, x1490, x1491, x1492, x1493, x1494, x1495, x1496, x1497, x1498, x1499, x1500, x1501, x1502, x1503, x1504, x1505, x1506, x1507, x1508, x1509, x1510, x1511, x1512, x1513, x1514, x1515, x1516, x1517, x1518, x1519, x1520, x1521, x1522, x1523, x1524, x1525, x1526, x1527, x1528, x1529, x1530, x1531, x1532, x1533, x1534, x1535, x1536, x1537, x1538, x1539, x1540, x1541, x1542, x1543, x1544, x1545, x1546, x1547, x1548, x1549, x1550, x1551, x1552, x1553, x1554, x1555, x1556, x1557, x1558, x1559, x1560, x1561, x1562, x1563, x1564, x1565, x1566, x1567, x1568, x1569, x1570, x1571, x1572, x1573, x1574, x1575, x1576, x1577, x1578, x1579, x1580, x1581, x1582, x1583, x1584, x1585, x1586, x1587, x1588, x1589, x1590, x1591, x1592, x1593, x1594, x1595, x1596, x1597, x1598, x1599, x1600, x1601, x1602, x1603, x1604, x1605, x1606, x1607, x1608, x1609, x1610, x1611, x1612, x1613, x1614, x1615, x1616, x1617, x1618, x1619, x1620, x1621, x1622, x1623, x1624, x1625, x1626, x1627, x1628, x1629, x1630, x1631, x1632, x1633, x1634, x1635, x1636, x1637, x1638, x1639, x1640, x1641, x1642, x1643, x1644, x1645, x1646, x1647, x1648, x1649, x1650, x1651, x1652, x1653, x1654, x1655, x1656, x1657, x1658, x1659, x1660, x1661, x1662, x1663, x1664, x1665, x1666, x1667, x1668, x1669, x1670, x1671, x1672, x1673, x1674, x1675, x1676, x1677, x1678, x1679, x1680, x1681, x1682, x1683, x1684, x1685, x1686, x1687, x1688, x1689, x1690, x1691, x1692, x1693, x1694, x1695, x1696, x1697, x1698, x1699, x1700, x1701, x1702, x1703, x1704, x1705, x1706, x1707, x1708, x1709, x1710, x1711, x1712, x1713, x1714, x1715, x1716, x1717, x1718, x1719, x1720, x1721, x1722, x1723, x1724, x1725, x1726, x1727, x1728, x1729, x1730, x1731, x1732, x1733, x1734, x1735, x1736, x1737, x1738, x1739, x1740, x1741, x1742, x1743, x1744, x1745, x1746, x1747, x1748, x1749, x1750, x1751, x1752, x1753, x1754, x1755, x1756, x1757, x1758, x1759, x1760, x1761, x1762, x1763, x1764, x1765, x1766, x1767, x1768, x1769, x1770, x1771, x1772, x1773, x1774, x1775, x1776, x1777, x1778, x1779, x1780, x1781, x1782, x1783, x1784, x1785, x1786, x1787, x1788, x1789, x1790, x1791, x1792, x1793, x1794, x1795, x1796, x1797, x1798, x1799, x1800, x1801, x1802, x1803, x1804, x1805, x1806, x1807, x1808, x1809, x1810, x1811, x1812, x1813, x1814, x1815, x1816, x1817, x1818, x1819, x1820, x1821, x1822, x1823, x1824, x1825, x1826, x1827, x1828, x1829, x1830, x1831, x1832, x1833, x1834, x1835, x1836, x1837, x1838, x1839, x1840, x1841, x1842, x1843, x1844, x1845, x1846, x1847, x1848, x1849, x1850, x1851, x1852, x1853, x1854, x1855, x1856, x1857, x1858, x1859, x1860, x1861, x1862, x1863, x1864, x1865, x1866, x1867, x1868, x1869, x1870, x1871, x1872, x1873, x1874, x1875, x1876, x1877, x1878, x1879, x1880, x1881, x1882, x1883, x1884, x1885, x1886, x1887, x1888, x1889, x1890, x1891, x1892, x1893, x1894, x1895, x1896, x1897, x1898, x1899, x1900, x1901, x1902, x1903, x1904, x1905, x1906, x1907, x1908, x1909, x1910, x1911, x1912, x1913, x1914, x1915, x1916, x1917, x1918, x1919, x1920, x1921, x1922, x1923, x1924, x1925, x1926, x1927, x1928, x1929, x1930, x1931, x1932, x1933, x1934, x1935, x1936, x1937, x1938, x1939, x1940, x1941, x1942, x1943, x1944, x1945, x1946, x1947, x1948, x1949, x1950, x1951, x1952, x1953, x1954, x1955, x1956, x1957, x1958, x1959, x1960, x1961, x1962, x1963, x1964, x1965, x1966, x1967, x1968, x1969, x1970, x1971, x1972, x1973, x1974, x1975, x1976, x1977, x1978, x1979, x1980, x1981, x1982, x1983, x1984, x1985, x1986, x1987, x1988, x1989, x1990, x1991, x1992, x1993, x1994, x1995, x1996, x1997, x1998, x1999, x2000, x2001, x2002, x2003, x2004, x2005, x2006, x2007, x2008, x2009, x2010, x2011, x2012, x2013, x2014, x2015, x2016, x2017, x2018, x2019, x2020, x2021, x2022, x2023, x2024, x2025, x2026, x2027, x2028, x2029, x2030, x2031, x2032, x2033, x2034, x2035, x2036, x2037, x2038, x2039, x2040, x2041, x2042, x2043, x2044, x2045, x2046, x2047, x2048, x2049, x2050, x2051, x2052, x2053, x2054, x2055, x2056, x2057, x2058, x2059, x2060, x2061, x2062, x2063, x2064, x2065, x2066, x2067, x2068, x2069, x2070, x2071, x2072, x2073, x2074, x2075, x2076, x2077, x2078, x2079, x2080, x2081, x2082, x2083, x2084, x2085, x2086, x2087, x2088, x2089, x2090, x2091, x2092, x2093, x2094, x2095, x2096, x2097, x2098, x2099, x2100, x2101, x2102, x2103, x2104, x2105, x2106, x2107, x2108, x2109, x2110, x2111, x2112, x2113, x2114, x2115, x2116, x2117, x2118, x2119, x2120, x2121, x2122, x2123, x2124, x2125, x2126, x2127, x2128, x2129, x2130, x2131, x2132, x2133, x2134, x2135, x2136, x2137, x2138, x2139, x2140, x2141, x2142, x2143, x2144, x2145, x2146, x2147, x2148, x2149, x2150, x2151, x2152, x2153, x2154, x2155, x2156, x2157, x2158, x2159, x2160, x2161, x2162, x2163, x2164, x2165, x2166, x2167, x2168, x2169, x2170, x2171, x2172, x2173, x2174, x2175, x2176, x2177, x2178, x2179, x2180, x2181, x2182, x2183, x2184, x2185, x2186, x2187, x2188, x2189, x2190, x2191, x2192, x2193, x2194, x2195, x2196, x2197, x2198, x2199, x2200, x2201, x2202, x2203, x2204, x2205, x2206, x2207, x2208, x2209, x2210, x2211, x2212, x2213, x2214, x2215, x2216, x2217, x2218, x2219, x2220, x2221, x2222, x2223, x2224, x2225, x2226, x2227, x2228, x2229, x2230, x2231, x2232, x2233, x2234, x2235, x2236, x2237, x2238, x2239, x2240, x2241, x2242, x2243, x2244, x2245, x2246, x2247, x2248, x2249, x2250, x2251, x2252, x2253, x2254, x2255, x2256, x2257, x2258, x2259, x2260, x2261, x2262, x2263, x2264, x2265, x2266, x2267, x2268, x2269, x2270, x2271, x2272, x2273, x2274, x2275, x2276, x2277, x2278, x2279, x2280, x2281, x2282, x2283, x2284, x2285, x2286, x2287, x2288, x2289, x2290, x2291, x2292, x2293, x2294, x2295, x2296, x2297, x2298, x2299, x2300, x2301, x2302, x2303, x2304, x2305, x2306, x2307, x2308, x2309, x2310, x2311, x2312, x2313, x2314, x2315, x2316, x2317, x2318, x2319, x2320, x2321, x2322, x2323, x2324, x2325, x2326, x2327, x2328, x2329, x2330, x2331, x2332, x2333, x2334, x2335, x2336, x2337, x2338, x2339, x2340, x2341, x2342, x2343, x2344, x2345, x2346, x2347, x2348, x2349, x2350, x2351, x2352, x2353, x2354, x2355, x2356, x2357, x2358, x2359, x2360, x2361, x2362, x2363, x2364, x2365, x2366, x2367, x2368, x2369, x2370, x2371, x2372, x2373, x2374, x2375, x2376, x2377, x2378, x2379, x2380, x2381, x2382, x2383, x2384, x2385, x2386, x2387, x2388, x2389, x2390, x2391, x2392, x2393, x2394, x2395, x2396, x2397, x2398, x2399, x2400, x2401, x2402, x2403, x2404, x2405, x2406, x2407, x2408, x2409, x2410, x2411, x2412, x2413, x2414, x2415, x2416, x2417, x2418, x2419, x2420, x2421, x2422, x2423, x2424, x2425, x2426, x2427, x2428, x2429, x2430, x2431, x2432, x2433, x2434, x2435, x2436, x2437, x2438, x2439, x2440, x2441, x2442, x2443, x2444, x2445, x2446, x2447, x2448, x2449, x2450, x2451, x2452, x2453, x2454, x2455, x2456, x2457, x2458, x2459, x2460, x2461, x2462, x2463, x2464, x2465, x2466, x2467, x2468, x2469, x2470, x2471, x2472, x2473, x2474, x2475, x2476, x2477, x2478, x2479, x2480, x2481, x2482, x2483, x2484, x2485, x2486, x2487, x2488, x2489, x2490, x2491, x2492, x2493, x2494, x2495, x2496, x2497, x2498, x2499, x2500, x2501, x2502, x2503, x2504, x2505, x2506, x2507, x2508, x2509, x2510, x2511, x2512, x2513, x2514, x2515, x2516, x2517, x2518, x2519, x2520, x2521, x2522, x2523, x2524, x2525, x2526, x2527, x2528, x2529, x2530, x2531, x2532, x2533, x2534, x2535, x2536, x2537, x2538, x2539, x2540, x2541, x2542, x2543, x2544, x2545, x2546, x2547, x2548, x2549, x2550, x2551, x2552, x2553, x2554, x2555, x2556, x2557, x2558, x2559, x2560, x2561, x2562, x2563, x2564, x2565, x2566, x2567, x2568, x2569, x2570, x2571, x2572, x2573, x2574, x2575, x2576, x2577, x2578, x2579, x2580, x2581, x2582, x2583, x2584, x2585, x2586, x2587, x2588, x2589, x2590, x2591, x2592, x2593, x2594, x2595, x2596, x2597, x2598, x2599, x2600, x2601, x2602, x2603, x2604, x2605, x2606, x2607, x2608, x2609, x2610, x2611, x2612, x2613, x2614, x2615, x2616, x2617, x2618, x2619, x2620, x2621, x2622, x2623, x2624, x2625, x2626, x2627, x2628, x2629, x2630, x2631, x2632, x2633, x2634, x2635, x2636, x2637, x2638, x2639, x2640, x2641, x2642, x2643, x2644, x2645, x2646, x2647, x2648, x2649, x2650, x2651, x2652, x2653, x2654, x2655, x2656, x2657, x2658, x2659, x2660, x2661, x2662, x2663, x2664, x2665, x2666, x2667, x2668, x2669, x2670, x2671, x2672, x2673, x2674, x2675, x2676, x2677, x2678, x2679, x2680, x2681, x2682, x2683, x2684, x2685, x2686, x2687, x2688, x2689, x2690, x2691, x2692, x2693, x2694, x2695, x2696, x2697, x2698, x2699, x2700, x2701, x2702, x2703, x2704, x2705, x2706, x2707, x2708, x2709, x2710, x2711, x2712, x2713, x2714, x2715, x2716, x2717, x2718, x2719, x2720, x2721, x2722, x2723, x2724, x2725, x2726, x2727, x2728, x2729, x2730, x2731, x2732, x2733, x2734, x2735, x2736, x2737, x2738, x2739, x2740, x2741, x2742, x2743, x2744, x2745, x2746, x2747, x2748, x2749, x2750, x2751, x2752, x2753, x2754, x2755, x2756, x2757, x2758, x2759, x2760, x2761, x2762, x2763, x2764, x2765, x2766, x2767, x2768, x2769, x2770, x2771, x2772, x2773, x2774, x2775, x2776, x2777, x2778, x2779, x2780, x2781, x2782, x2783, x2784, x2785, x2786, x2787, x2788, x2789, x2790, x2791, x2792, x2793, x2794, x2795, x2796, x2797, x2798, x2799, x2800, x2801, x2802, x2803, x2804, x2805, x2806, x2807, x2808, x2809, x2810, x2811, x2812, x2813, x2814, x2815, x2816, x2817, x2818, x2819, x2820, x2821, x2822, x2823, x2824, x2825, x2826, x2827, x2828, x2829, x2830, x2831, x2832, x2833, x2834, x2835, x2836, x2837, x2838, x2839, x2840, x2841, x2842, x2843, x2844, x2845, x2846, x2847, x2848, x2849, x2850, x2851, x2852, x2853, x2854, x2855, x2856, x2857, x2858, x2859, x2860, x2861, x2862, x2863, x2864, x2865, x2866, x2867, x2868, x2869, x2870, x2871, x2872, x2873, x2874, x2875, x2876, x2877, x2878, x2879, x2880, x2881, x2882, x2883, x2884, x2885, x2886, x2887, x2888, x2889, x2890, x2891, x2892, x2893, x2894, x2895, x2896, x2897, x2898, x2899, x2900, x2901, x2902, x2903, x2904, x2905, x2906, x2907, x2908, x2909, x2910, x2911, x2912, x2913, x2914, x2915, x2916, x2917, x2918, x2919, x2920, x2921, x2922, x2923, x2924, x2925, x2926, x2927, x2928, x2929, x2930, x2931, x2932, x2933, x2934, x2935, x2936, x2937, x2938, x2939, x2940, x2941, x2942, x2943, x2944, x2945, x2946, x2947, x2948, x2949, x2950, x2951, x2952, x2953, x2954, x2955, x2956, x2957, x2958, x2959, x2960, x2961, x2962, x2963, x2964, x2965, x2966, x2967, x2968, x2969, x2970, x2971, x2972, x2973, x2974, x2975, x2976, x2977, x2978, x2979, x2980, x2981, x2982, x2983, x2984, x2985, x2986, x2987, x2988, x2989, x2990, x2991, x2992, x2993, x2994, x2995, x2996, x2997, x2998, x2999, x3000;
  output y0;
  wire n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969;
  LUT3 #(.INIT(8'hE8)) lut_n3003 (.I0(x0), .I1(x1), .I2(x2), .O(n3003));
  LUT3 #(.INIT(8'hE8)) lut_n3004 (.I0(x6), .I1(x7), .I2(x8), .O(n3004));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3005 (.I0(x3), .I1(x4), .I2(x5), .I3(n3003), .I4(n3004), .O(n3005));
  LUT3 #(.INIT(8'hE8)) lut_n3006 (.I0(x12), .I1(x13), .I2(x14), .O(n3006));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3007 (.I0(x3), .I1(x4), .I2(x5), .I3(n3003), .I4(n3004), .O(n3007));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3008 (.I0(x9), .I1(x10), .I2(x11), .I3(n3006), .I4(n3007), .O(n3008));
  LUT3 #(.INIT(8'hE8)) lut_n3009 (.I0(x18), .I1(x19), .I2(x20), .O(n3009));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3010 (.I0(x9), .I1(x10), .I2(x11), .I3(n3006), .I4(n3007), .O(n3010));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3011 (.I0(x15), .I1(x16), .I2(x17), .I3(n3009), .I4(n3010), .O(n3011));
  LUT3 #(.INIT(8'hE8)) lut_n3012 (.I0(n3005), .I1(n3008), .I2(n3011), .O(n3012));
  LUT3 #(.INIT(8'hE8)) lut_n3013 (.I0(x24), .I1(x25), .I2(x26), .O(n3013));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3014 (.I0(x15), .I1(x16), .I2(x17), .I3(n3009), .I4(n3010), .O(n3014));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3015 (.I0(x21), .I1(x22), .I2(x23), .I3(n3013), .I4(n3014), .O(n3015));
  LUT3 #(.INIT(8'hE8)) lut_n3016 (.I0(x27), .I1(x28), .I2(x29), .O(n3016));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3017 (.I0(x21), .I1(x22), .I2(x23), .I3(n3013), .I4(n3014), .O(n3017));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3018 (.I0(x30), .I1(x31), .I2(x32), .I3(n3016), .I4(n3017), .O(n3018));
  LUT3 #(.INIT(8'h96)) lut_n3019 (.I0(n3005), .I1(n3008), .I2(n3011), .O(n3019));
  LUT3 #(.INIT(8'hE8)) lut_n3020 (.I0(n3015), .I1(n3018), .I2(n3019), .O(n3020));
  LUT3 #(.INIT(8'hE8)) lut_n3021 (.I0(x36), .I1(x37), .I2(x38), .O(n3021));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3022 (.I0(x30), .I1(x31), .I2(x32), .I3(n3016), .I4(n3017), .O(n3022));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3023 (.I0(x33), .I1(x34), .I2(x35), .I3(n3021), .I4(n3022), .O(n3023));
  LUT3 #(.INIT(8'hE8)) lut_n3024 (.I0(x42), .I1(x43), .I2(x44), .O(n3024));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3025 (.I0(x33), .I1(x34), .I2(x35), .I3(n3021), .I4(n3022), .O(n3025));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3026 (.I0(x39), .I1(x40), .I2(x41), .I3(n3024), .I4(n3025), .O(n3026));
  LUT3 #(.INIT(8'h96)) lut_n3027 (.I0(n3015), .I1(n3018), .I2(n3019), .O(n3027));
  LUT3 #(.INIT(8'hE8)) lut_n3028 (.I0(n3023), .I1(n3026), .I2(n3027), .O(n3028));
  LUT3 #(.INIT(8'hE8)) lut_n3029 (.I0(n3012), .I1(n3020), .I2(n3028), .O(n3029));
  LUT3 #(.INIT(8'hE8)) lut_n3030 (.I0(x48), .I1(x49), .I2(x50), .O(n3030));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3031 (.I0(x39), .I1(x40), .I2(x41), .I3(n3024), .I4(n3025), .O(n3031));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3032 (.I0(x45), .I1(x46), .I2(x47), .I3(n3030), .I4(n3031), .O(n3032));
  LUT3 #(.INIT(8'hE8)) lut_n3033 (.I0(x54), .I1(x55), .I2(x56), .O(n3033));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3034 (.I0(x45), .I1(x46), .I2(x47), .I3(n3030), .I4(n3031), .O(n3034));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3035 (.I0(x51), .I1(x52), .I2(x53), .I3(n3033), .I4(n3034), .O(n3035));
  LUT3 #(.INIT(8'h96)) lut_n3036 (.I0(n3023), .I1(n3026), .I2(n3027), .O(n3036));
  LUT3 #(.INIT(8'hE8)) lut_n3037 (.I0(n3032), .I1(n3035), .I2(n3036), .O(n3037));
  LUT3 #(.INIT(8'hE8)) lut_n3038 (.I0(x60), .I1(x61), .I2(x62), .O(n3038));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3039 (.I0(x51), .I1(x52), .I2(x53), .I3(n3033), .I4(n3034), .O(n3039));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3040 (.I0(x57), .I1(x58), .I2(x59), .I3(n3038), .I4(n3039), .O(n3040));
  LUT3 #(.INIT(8'hE8)) lut_n3041 (.I0(x66), .I1(x67), .I2(x68), .O(n3041));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3042 (.I0(x57), .I1(x58), .I2(x59), .I3(n3038), .I4(n3039), .O(n3042));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3043 (.I0(x63), .I1(x64), .I2(x65), .I3(n3041), .I4(n3042), .O(n3043));
  LUT3 #(.INIT(8'h96)) lut_n3044 (.I0(n3032), .I1(n3035), .I2(n3036), .O(n3044));
  LUT3 #(.INIT(8'hE8)) lut_n3045 (.I0(n3040), .I1(n3043), .I2(n3044), .O(n3045));
  LUT3 #(.INIT(8'h96)) lut_n3046 (.I0(n3012), .I1(n3020), .I2(n3028), .O(n3046));
  LUT3 #(.INIT(8'hE8)) lut_n3047 (.I0(n3037), .I1(n3045), .I2(n3046), .O(n3047));
  LUT3 #(.INIT(8'hE8)) lut_n3048 (.I0(x72), .I1(x73), .I2(x74), .O(n3048));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3049 (.I0(x63), .I1(x64), .I2(x65), .I3(n3041), .I4(n3042), .O(n3049));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3050 (.I0(x69), .I1(x70), .I2(x71), .I3(n3048), .I4(n3049), .O(n3050));
  LUT3 #(.INIT(8'hE8)) lut_n3051 (.I0(x78), .I1(x79), .I2(x80), .O(n3051));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3052 (.I0(x69), .I1(x70), .I2(x71), .I3(n3048), .I4(n3049), .O(n3052));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3053 (.I0(x75), .I1(x76), .I2(x77), .I3(n3051), .I4(n3052), .O(n3053));
  LUT3 #(.INIT(8'h96)) lut_n3054 (.I0(n3040), .I1(n3043), .I2(n3044), .O(n3054));
  LUT3 #(.INIT(8'hE8)) lut_n3055 (.I0(n3050), .I1(n3053), .I2(n3054), .O(n3055));
  LUT3 #(.INIT(8'hE8)) lut_n3056 (.I0(x84), .I1(x85), .I2(x86), .O(n3056));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3057 (.I0(x75), .I1(x76), .I2(x77), .I3(n3051), .I4(n3052), .O(n3057));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3058 (.I0(x81), .I1(x82), .I2(x83), .I3(n3056), .I4(n3057), .O(n3058));
  LUT3 #(.INIT(8'hE8)) lut_n3059 (.I0(x90), .I1(x91), .I2(x92), .O(n3059));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3060 (.I0(x81), .I1(x82), .I2(x83), .I3(n3056), .I4(n3057), .O(n3060));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3061 (.I0(x87), .I1(x88), .I2(x89), .I3(n3059), .I4(n3060), .O(n3061));
  LUT3 #(.INIT(8'h96)) lut_n3062 (.I0(n3050), .I1(n3053), .I2(n3054), .O(n3062));
  LUT3 #(.INIT(8'hE8)) lut_n3063 (.I0(n3058), .I1(n3061), .I2(n3062), .O(n3063));
  LUT3 #(.INIT(8'h96)) lut_n3064 (.I0(n3037), .I1(n3045), .I2(n3046), .O(n3064));
  LUT3 #(.INIT(8'hE8)) lut_n3065 (.I0(n3055), .I1(n3063), .I2(n3064), .O(n3065));
  LUT3 #(.INIT(8'hE8)) lut_n3066 (.I0(n3029), .I1(n3047), .I2(n3065), .O(n3066));
  LUT3 #(.INIT(8'hE8)) lut_n3067 (.I0(x96), .I1(x97), .I2(x98), .O(n3067));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3068 (.I0(x87), .I1(x88), .I2(x89), .I3(n3059), .I4(n3060), .O(n3068));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3069 (.I0(x93), .I1(x94), .I2(x95), .I3(n3067), .I4(n3068), .O(n3069));
  LUT3 #(.INIT(8'hE8)) lut_n3070 (.I0(x102), .I1(x103), .I2(x104), .O(n3070));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3071 (.I0(x93), .I1(x94), .I2(x95), .I3(n3067), .I4(n3068), .O(n3071));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3072 (.I0(x99), .I1(x100), .I2(x101), .I3(n3070), .I4(n3071), .O(n3072));
  LUT3 #(.INIT(8'h96)) lut_n3073 (.I0(n3058), .I1(n3061), .I2(n3062), .O(n3073));
  LUT3 #(.INIT(8'hE8)) lut_n3074 (.I0(n3069), .I1(n3072), .I2(n3073), .O(n3074));
  LUT3 #(.INIT(8'hE8)) lut_n3075 (.I0(x108), .I1(x109), .I2(x110), .O(n3075));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3076 (.I0(x99), .I1(x100), .I2(x101), .I3(n3070), .I4(n3071), .O(n3076));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3077 (.I0(x105), .I1(x106), .I2(x107), .I3(n3075), .I4(n3076), .O(n3077));
  LUT3 #(.INIT(8'hE8)) lut_n3078 (.I0(x114), .I1(x115), .I2(x116), .O(n3078));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3079 (.I0(x105), .I1(x106), .I2(x107), .I3(n3075), .I4(n3076), .O(n3079));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3080 (.I0(x111), .I1(x112), .I2(x113), .I3(n3078), .I4(n3079), .O(n3080));
  LUT3 #(.INIT(8'h96)) lut_n3081 (.I0(n3069), .I1(n3072), .I2(n3073), .O(n3081));
  LUT3 #(.INIT(8'hE8)) lut_n3082 (.I0(n3077), .I1(n3080), .I2(n3081), .O(n3082));
  LUT3 #(.INIT(8'h96)) lut_n3083 (.I0(n3055), .I1(n3063), .I2(n3064), .O(n3083));
  LUT3 #(.INIT(8'hE8)) lut_n3084 (.I0(n3074), .I1(n3082), .I2(n3083), .O(n3084));
  LUT3 #(.INIT(8'hE8)) lut_n3085 (.I0(x120), .I1(x121), .I2(x122), .O(n3085));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3086 (.I0(x111), .I1(x112), .I2(x113), .I3(n3078), .I4(n3079), .O(n3086));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3087 (.I0(x117), .I1(x118), .I2(x119), .I3(n3085), .I4(n3086), .O(n3087));
  LUT3 #(.INIT(8'hE8)) lut_n3088 (.I0(x126), .I1(x127), .I2(x128), .O(n3088));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3089 (.I0(x117), .I1(x118), .I2(x119), .I3(n3085), .I4(n3086), .O(n3089));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3090 (.I0(x123), .I1(x124), .I2(x125), .I3(n3088), .I4(n3089), .O(n3090));
  LUT3 #(.INIT(8'h96)) lut_n3091 (.I0(n3077), .I1(n3080), .I2(n3081), .O(n3091));
  LUT3 #(.INIT(8'hE8)) lut_n3092 (.I0(n3087), .I1(n3090), .I2(n3091), .O(n3092));
  LUT3 #(.INIT(8'hE8)) lut_n3093 (.I0(x132), .I1(x133), .I2(x134), .O(n3093));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3094 (.I0(x123), .I1(x124), .I2(x125), .I3(n3088), .I4(n3089), .O(n3094));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3095 (.I0(x129), .I1(x130), .I2(x131), .I3(n3093), .I4(n3094), .O(n3095));
  LUT3 #(.INIT(8'hE8)) lut_n3096 (.I0(x138), .I1(x139), .I2(x140), .O(n3096));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3097 (.I0(x129), .I1(x130), .I2(x131), .I3(n3093), .I4(n3094), .O(n3097));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3098 (.I0(x135), .I1(x136), .I2(x137), .I3(n3096), .I4(n3097), .O(n3098));
  LUT3 #(.INIT(8'h96)) lut_n3099 (.I0(n3087), .I1(n3090), .I2(n3091), .O(n3099));
  LUT3 #(.INIT(8'hE8)) lut_n3100 (.I0(n3095), .I1(n3098), .I2(n3099), .O(n3100));
  LUT3 #(.INIT(8'h96)) lut_n3101 (.I0(n3074), .I1(n3082), .I2(n3083), .O(n3101));
  LUT3 #(.INIT(8'hE8)) lut_n3102 (.I0(n3092), .I1(n3100), .I2(n3101), .O(n3102));
  LUT3 #(.INIT(8'h96)) lut_n3103 (.I0(n3029), .I1(n3047), .I2(n3065), .O(n3103));
  LUT3 #(.INIT(8'hE8)) lut_n3104 (.I0(n3084), .I1(n3102), .I2(n3103), .O(n3104));
  LUT3 #(.INIT(8'hE8)) lut_n3105 (.I0(x144), .I1(x145), .I2(x146), .O(n3105));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3106 (.I0(x135), .I1(x136), .I2(x137), .I3(n3096), .I4(n3097), .O(n3106));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3107 (.I0(x141), .I1(x142), .I2(x143), .I3(n3105), .I4(n3106), .O(n3107));
  LUT3 #(.INIT(8'hE8)) lut_n3108 (.I0(x150), .I1(x151), .I2(x152), .O(n3108));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3109 (.I0(x141), .I1(x142), .I2(x143), .I3(n3105), .I4(n3106), .O(n3109));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3110 (.I0(x147), .I1(x148), .I2(x149), .I3(n3108), .I4(n3109), .O(n3110));
  LUT3 #(.INIT(8'h96)) lut_n3111 (.I0(n3095), .I1(n3098), .I2(n3099), .O(n3111));
  LUT3 #(.INIT(8'hE8)) lut_n3112 (.I0(n3107), .I1(n3110), .I2(n3111), .O(n3112));
  LUT3 #(.INIT(8'hE8)) lut_n3113 (.I0(x156), .I1(x157), .I2(x158), .O(n3113));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3114 (.I0(x147), .I1(x148), .I2(x149), .I3(n3108), .I4(n3109), .O(n3114));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3115 (.I0(x153), .I1(x154), .I2(x155), .I3(n3113), .I4(n3114), .O(n3115));
  LUT3 #(.INIT(8'hE8)) lut_n3116 (.I0(x162), .I1(x163), .I2(x164), .O(n3116));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3117 (.I0(x153), .I1(x154), .I2(x155), .I3(n3113), .I4(n3114), .O(n3117));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3118 (.I0(x159), .I1(x160), .I2(x161), .I3(n3116), .I4(n3117), .O(n3118));
  LUT3 #(.INIT(8'h96)) lut_n3119 (.I0(n3107), .I1(n3110), .I2(n3111), .O(n3119));
  LUT3 #(.INIT(8'hE8)) lut_n3120 (.I0(n3115), .I1(n3118), .I2(n3119), .O(n3120));
  LUT3 #(.INIT(8'h96)) lut_n3121 (.I0(n3092), .I1(n3100), .I2(n3101), .O(n3121));
  LUT3 #(.INIT(8'hE8)) lut_n3122 (.I0(n3112), .I1(n3120), .I2(n3121), .O(n3122));
  LUT3 #(.INIT(8'hE8)) lut_n3123 (.I0(x168), .I1(x169), .I2(x170), .O(n3123));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3124 (.I0(x159), .I1(x160), .I2(x161), .I3(n3116), .I4(n3117), .O(n3124));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3125 (.I0(x165), .I1(x166), .I2(x167), .I3(n3123), .I4(n3124), .O(n3125));
  LUT3 #(.INIT(8'hE8)) lut_n3126 (.I0(x174), .I1(x175), .I2(x176), .O(n3126));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3127 (.I0(x165), .I1(x166), .I2(x167), .I3(n3123), .I4(n3124), .O(n3127));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3128 (.I0(x171), .I1(x172), .I2(x173), .I3(n3126), .I4(n3127), .O(n3128));
  LUT3 #(.INIT(8'h96)) lut_n3129 (.I0(n3115), .I1(n3118), .I2(n3119), .O(n3129));
  LUT3 #(.INIT(8'hE8)) lut_n3130 (.I0(n3125), .I1(n3128), .I2(n3129), .O(n3130));
  LUT3 #(.INIT(8'hE8)) lut_n3131 (.I0(x180), .I1(x181), .I2(x182), .O(n3131));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3132 (.I0(x171), .I1(x172), .I2(x173), .I3(n3126), .I4(n3127), .O(n3132));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3133 (.I0(x177), .I1(x178), .I2(x179), .I3(n3131), .I4(n3132), .O(n3133));
  LUT3 #(.INIT(8'hE8)) lut_n3134 (.I0(x186), .I1(x187), .I2(x188), .O(n3134));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3135 (.I0(x177), .I1(x178), .I2(x179), .I3(n3131), .I4(n3132), .O(n3135));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3136 (.I0(x183), .I1(x184), .I2(x185), .I3(n3134), .I4(n3135), .O(n3136));
  LUT3 #(.INIT(8'h96)) lut_n3137 (.I0(n3125), .I1(n3128), .I2(n3129), .O(n3137));
  LUT3 #(.INIT(8'hE8)) lut_n3138 (.I0(n3133), .I1(n3136), .I2(n3137), .O(n3138));
  LUT3 #(.INIT(8'h96)) lut_n3139 (.I0(n3112), .I1(n3120), .I2(n3121), .O(n3139));
  LUT3 #(.INIT(8'hE8)) lut_n3140 (.I0(n3130), .I1(n3138), .I2(n3139), .O(n3140));
  LUT3 #(.INIT(8'h96)) lut_n3141 (.I0(n3084), .I1(n3102), .I2(n3103), .O(n3141));
  LUT3 #(.INIT(8'hE8)) lut_n3142 (.I0(n3122), .I1(n3140), .I2(n3141), .O(n3142));
  LUT3 #(.INIT(8'hE8)) lut_n3143 (.I0(n3066), .I1(n3104), .I2(n3142), .O(n3143));
  LUT3 #(.INIT(8'hE8)) lut_n3144 (.I0(x192), .I1(x193), .I2(x194), .O(n3144));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3145 (.I0(x183), .I1(x184), .I2(x185), .I3(n3134), .I4(n3135), .O(n3145));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3146 (.I0(x189), .I1(x190), .I2(x191), .I3(n3144), .I4(n3145), .O(n3146));
  LUT3 #(.INIT(8'hE8)) lut_n3147 (.I0(x198), .I1(x199), .I2(x200), .O(n3147));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3148 (.I0(x189), .I1(x190), .I2(x191), .I3(n3144), .I4(n3145), .O(n3148));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3149 (.I0(x195), .I1(x196), .I2(x197), .I3(n3147), .I4(n3148), .O(n3149));
  LUT3 #(.INIT(8'h96)) lut_n3150 (.I0(n3133), .I1(n3136), .I2(n3137), .O(n3150));
  LUT3 #(.INIT(8'hE8)) lut_n3151 (.I0(n3146), .I1(n3149), .I2(n3150), .O(n3151));
  LUT3 #(.INIT(8'hE8)) lut_n3152 (.I0(x204), .I1(x205), .I2(x206), .O(n3152));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3153 (.I0(x195), .I1(x196), .I2(x197), .I3(n3147), .I4(n3148), .O(n3153));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3154 (.I0(x201), .I1(x202), .I2(x203), .I3(n3152), .I4(n3153), .O(n3154));
  LUT3 #(.INIT(8'hE8)) lut_n3155 (.I0(x210), .I1(x211), .I2(x212), .O(n3155));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3156 (.I0(x201), .I1(x202), .I2(x203), .I3(n3152), .I4(n3153), .O(n3156));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3157 (.I0(x207), .I1(x208), .I2(x209), .I3(n3155), .I4(n3156), .O(n3157));
  LUT3 #(.INIT(8'h96)) lut_n3158 (.I0(n3146), .I1(n3149), .I2(n3150), .O(n3158));
  LUT3 #(.INIT(8'hE8)) lut_n3159 (.I0(n3154), .I1(n3157), .I2(n3158), .O(n3159));
  LUT3 #(.INIT(8'h96)) lut_n3160 (.I0(n3130), .I1(n3138), .I2(n3139), .O(n3160));
  LUT3 #(.INIT(8'hE8)) lut_n3161 (.I0(n3151), .I1(n3159), .I2(n3160), .O(n3161));
  LUT3 #(.INIT(8'hE8)) lut_n3162 (.I0(x216), .I1(x217), .I2(x218), .O(n3162));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3163 (.I0(x207), .I1(x208), .I2(x209), .I3(n3155), .I4(n3156), .O(n3163));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3164 (.I0(x213), .I1(x214), .I2(x215), .I3(n3162), .I4(n3163), .O(n3164));
  LUT3 #(.INIT(8'hE8)) lut_n3165 (.I0(x222), .I1(x223), .I2(x224), .O(n3165));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3166 (.I0(x213), .I1(x214), .I2(x215), .I3(n3162), .I4(n3163), .O(n3166));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3167 (.I0(x219), .I1(x220), .I2(x221), .I3(n3165), .I4(n3166), .O(n3167));
  LUT3 #(.INIT(8'h96)) lut_n3168 (.I0(n3154), .I1(n3157), .I2(n3158), .O(n3168));
  LUT3 #(.INIT(8'hE8)) lut_n3169 (.I0(n3164), .I1(n3167), .I2(n3168), .O(n3169));
  LUT3 #(.INIT(8'hE8)) lut_n3170 (.I0(x228), .I1(x229), .I2(x230), .O(n3170));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3171 (.I0(x219), .I1(x220), .I2(x221), .I3(n3165), .I4(n3166), .O(n3171));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3172 (.I0(x225), .I1(x226), .I2(x227), .I3(n3170), .I4(n3171), .O(n3172));
  LUT3 #(.INIT(8'hE8)) lut_n3173 (.I0(x234), .I1(x235), .I2(x236), .O(n3173));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3174 (.I0(x225), .I1(x226), .I2(x227), .I3(n3170), .I4(n3171), .O(n3174));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3175 (.I0(x231), .I1(x232), .I2(x233), .I3(n3173), .I4(n3174), .O(n3175));
  LUT3 #(.INIT(8'h96)) lut_n3176 (.I0(n3164), .I1(n3167), .I2(n3168), .O(n3176));
  LUT3 #(.INIT(8'hE8)) lut_n3177 (.I0(n3172), .I1(n3175), .I2(n3176), .O(n3177));
  LUT3 #(.INIT(8'h96)) lut_n3178 (.I0(n3151), .I1(n3159), .I2(n3160), .O(n3178));
  LUT3 #(.INIT(8'hE8)) lut_n3179 (.I0(n3169), .I1(n3177), .I2(n3178), .O(n3179));
  LUT3 #(.INIT(8'h96)) lut_n3180 (.I0(n3122), .I1(n3140), .I2(n3141), .O(n3180));
  LUT3 #(.INIT(8'hE8)) lut_n3181 (.I0(n3161), .I1(n3179), .I2(n3180), .O(n3181));
  LUT3 #(.INIT(8'hE8)) lut_n3182 (.I0(x240), .I1(x241), .I2(x242), .O(n3182));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3183 (.I0(x231), .I1(x232), .I2(x233), .I3(n3173), .I4(n3174), .O(n3183));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3184 (.I0(x237), .I1(x238), .I2(x239), .I3(n3182), .I4(n3183), .O(n3184));
  LUT3 #(.INIT(8'hE8)) lut_n3185 (.I0(x246), .I1(x247), .I2(x248), .O(n3185));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3186 (.I0(x237), .I1(x238), .I2(x239), .I3(n3182), .I4(n3183), .O(n3186));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3187 (.I0(x243), .I1(x244), .I2(x245), .I3(n3185), .I4(n3186), .O(n3187));
  LUT3 #(.INIT(8'h96)) lut_n3188 (.I0(n3172), .I1(n3175), .I2(n3176), .O(n3188));
  LUT3 #(.INIT(8'hE8)) lut_n3189 (.I0(n3184), .I1(n3187), .I2(n3188), .O(n3189));
  LUT3 #(.INIT(8'hE8)) lut_n3190 (.I0(x252), .I1(x253), .I2(x254), .O(n3190));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3191 (.I0(x243), .I1(x244), .I2(x245), .I3(n3185), .I4(n3186), .O(n3191));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3192 (.I0(x249), .I1(x250), .I2(x251), .I3(n3190), .I4(n3191), .O(n3192));
  LUT3 #(.INIT(8'hE8)) lut_n3193 (.I0(x258), .I1(x259), .I2(x260), .O(n3193));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3194 (.I0(x249), .I1(x250), .I2(x251), .I3(n3190), .I4(n3191), .O(n3194));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3195 (.I0(x255), .I1(x256), .I2(x257), .I3(n3193), .I4(n3194), .O(n3195));
  LUT3 #(.INIT(8'h96)) lut_n3196 (.I0(n3184), .I1(n3187), .I2(n3188), .O(n3196));
  LUT3 #(.INIT(8'hE8)) lut_n3197 (.I0(n3192), .I1(n3195), .I2(n3196), .O(n3197));
  LUT3 #(.INIT(8'h96)) lut_n3198 (.I0(n3169), .I1(n3177), .I2(n3178), .O(n3198));
  LUT3 #(.INIT(8'hE8)) lut_n3199 (.I0(n3189), .I1(n3197), .I2(n3198), .O(n3199));
  LUT3 #(.INIT(8'hE8)) lut_n3200 (.I0(x264), .I1(x265), .I2(x266), .O(n3200));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3201 (.I0(x255), .I1(x256), .I2(x257), .I3(n3193), .I4(n3194), .O(n3201));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3202 (.I0(x261), .I1(x262), .I2(x263), .I3(n3200), .I4(n3201), .O(n3202));
  LUT3 #(.INIT(8'hE8)) lut_n3203 (.I0(x270), .I1(x271), .I2(x272), .O(n3203));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3204 (.I0(x261), .I1(x262), .I2(x263), .I3(n3200), .I4(n3201), .O(n3204));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3205 (.I0(x267), .I1(x268), .I2(x269), .I3(n3203), .I4(n3204), .O(n3205));
  LUT3 #(.INIT(8'h96)) lut_n3206 (.I0(n3192), .I1(n3195), .I2(n3196), .O(n3206));
  LUT3 #(.INIT(8'hE8)) lut_n3207 (.I0(n3202), .I1(n3205), .I2(n3206), .O(n3207));
  LUT3 #(.INIT(8'hE8)) lut_n3208 (.I0(x276), .I1(x277), .I2(x278), .O(n3208));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3209 (.I0(x267), .I1(x268), .I2(x269), .I3(n3203), .I4(n3204), .O(n3209));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3210 (.I0(x273), .I1(x274), .I2(x275), .I3(n3208), .I4(n3209), .O(n3210));
  LUT3 #(.INIT(8'hE8)) lut_n3211 (.I0(x282), .I1(x283), .I2(x284), .O(n3211));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3212 (.I0(x273), .I1(x274), .I2(x275), .I3(n3208), .I4(n3209), .O(n3212));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3213 (.I0(x279), .I1(x280), .I2(x281), .I3(n3211), .I4(n3212), .O(n3213));
  LUT3 #(.INIT(8'h96)) lut_n3214 (.I0(n3202), .I1(n3205), .I2(n3206), .O(n3214));
  LUT3 #(.INIT(8'hE8)) lut_n3215 (.I0(n3210), .I1(n3213), .I2(n3214), .O(n3215));
  LUT3 #(.INIT(8'h96)) lut_n3216 (.I0(n3189), .I1(n3197), .I2(n3198), .O(n3216));
  LUT3 #(.INIT(8'hE8)) lut_n3217 (.I0(n3207), .I1(n3215), .I2(n3216), .O(n3217));
  LUT3 #(.INIT(8'h96)) lut_n3218 (.I0(n3161), .I1(n3179), .I2(n3180), .O(n3218));
  LUT3 #(.INIT(8'hE8)) lut_n3219 (.I0(n3199), .I1(n3217), .I2(n3218), .O(n3219));
  LUT3 #(.INIT(8'h96)) lut_n3220 (.I0(n3066), .I1(n3104), .I2(n3142), .O(n3220));
  LUT3 #(.INIT(8'hE8)) lut_n3221 (.I0(n3181), .I1(n3219), .I2(n3220), .O(n3221));
  LUT3 #(.INIT(8'hE8)) lut_n3222 (.I0(x288), .I1(x289), .I2(x290), .O(n3222));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3223 (.I0(x279), .I1(x280), .I2(x281), .I3(n3211), .I4(n3212), .O(n3223));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3224 (.I0(x285), .I1(x286), .I2(x287), .I3(n3222), .I4(n3223), .O(n3224));
  LUT3 #(.INIT(8'hE8)) lut_n3225 (.I0(x294), .I1(x295), .I2(x296), .O(n3225));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3226 (.I0(x285), .I1(x286), .I2(x287), .I3(n3222), .I4(n3223), .O(n3226));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3227 (.I0(x291), .I1(x292), .I2(x293), .I3(n3225), .I4(n3226), .O(n3227));
  LUT3 #(.INIT(8'h96)) lut_n3228 (.I0(n3210), .I1(n3213), .I2(n3214), .O(n3228));
  LUT3 #(.INIT(8'hE8)) lut_n3229 (.I0(n3224), .I1(n3227), .I2(n3228), .O(n3229));
  LUT3 #(.INIT(8'hE8)) lut_n3230 (.I0(x297), .I1(x298), .I2(x299), .O(n3230));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3231 (.I0(x291), .I1(x292), .I2(x293), .I3(n3225), .I4(n3226), .O(n3231));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3232 (.I0(x300), .I1(x301), .I2(x302), .I3(n3230), .I4(n3231), .O(n3232));
  LUT3 #(.INIT(8'hE8)) lut_n3233 (.I0(x306), .I1(x307), .I2(x308), .O(n3233));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3234 (.I0(x300), .I1(x301), .I2(x302), .I3(n3230), .I4(n3231), .O(n3234));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3235 (.I0(x303), .I1(x304), .I2(x305), .I3(n3233), .I4(n3234), .O(n3235));
  LUT3 #(.INIT(8'h96)) lut_n3236 (.I0(n3224), .I1(n3227), .I2(n3228), .O(n3236));
  LUT3 #(.INIT(8'hE8)) lut_n3237 (.I0(n3232), .I1(n3235), .I2(n3236), .O(n3237));
  LUT3 #(.INIT(8'h96)) lut_n3238 (.I0(n3207), .I1(n3215), .I2(n3216), .O(n3238));
  LUT3 #(.INIT(8'hE8)) lut_n3239 (.I0(n3229), .I1(n3237), .I2(n3238), .O(n3239));
  LUT3 #(.INIT(8'hE8)) lut_n3240 (.I0(x312), .I1(x313), .I2(x314), .O(n3240));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3241 (.I0(x303), .I1(x304), .I2(x305), .I3(n3233), .I4(n3234), .O(n3241));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3242 (.I0(x309), .I1(x310), .I2(x311), .I3(n3240), .I4(n3241), .O(n3242));
  LUT3 #(.INIT(8'hE8)) lut_n3243 (.I0(x318), .I1(x319), .I2(x320), .O(n3243));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3244 (.I0(x309), .I1(x310), .I2(x311), .I3(n3240), .I4(n3241), .O(n3244));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3245 (.I0(x315), .I1(x316), .I2(x317), .I3(n3243), .I4(n3244), .O(n3245));
  LUT3 #(.INIT(8'h96)) lut_n3246 (.I0(n3232), .I1(n3235), .I2(n3236), .O(n3246));
  LUT3 #(.INIT(8'hE8)) lut_n3247 (.I0(n3242), .I1(n3245), .I2(n3246), .O(n3247));
  LUT3 #(.INIT(8'hE8)) lut_n3248 (.I0(x324), .I1(x325), .I2(x326), .O(n3248));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3249 (.I0(x315), .I1(x316), .I2(x317), .I3(n3243), .I4(n3244), .O(n3249));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3250 (.I0(x321), .I1(x322), .I2(x323), .I3(n3248), .I4(n3249), .O(n3250));
  LUT3 #(.INIT(8'hE8)) lut_n3251 (.I0(x330), .I1(x331), .I2(x332), .O(n3251));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3252 (.I0(x321), .I1(x322), .I2(x323), .I3(n3248), .I4(n3249), .O(n3252));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3253 (.I0(x327), .I1(x328), .I2(x329), .I3(n3251), .I4(n3252), .O(n3253));
  LUT3 #(.INIT(8'h96)) lut_n3254 (.I0(n3242), .I1(n3245), .I2(n3246), .O(n3254));
  LUT3 #(.INIT(8'hE8)) lut_n3255 (.I0(n3250), .I1(n3253), .I2(n3254), .O(n3255));
  LUT3 #(.INIT(8'h96)) lut_n3256 (.I0(n3229), .I1(n3237), .I2(n3238), .O(n3256));
  LUT3 #(.INIT(8'hE8)) lut_n3257 (.I0(n3247), .I1(n3255), .I2(n3256), .O(n3257));
  LUT3 #(.INIT(8'h96)) lut_n3258 (.I0(n3199), .I1(n3217), .I2(n3218), .O(n3258));
  LUT3 #(.INIT(8'hE8)) lut_n3259 (.I0(n3239), .I1(n3257), .I2(n3258), .O(n3259));
  LUT3 #(.INIT(8'hE8)) lut_n3260 (.I0(x336), .I1(x337), .I2(x338), .O(n3260));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3261 (.I0(x327), .I1(x328), .I2(x329), .I3(n3251), .I4(n3252), .O(n3261));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3262 (.I0(x333), .I1(x334), .I2(x335), .I3(n3260), .I4(n3261), .O(n3262));
  LUT3 #(.INIT(8'hE8)) lut_n3263 (.I0(x342), .I1(x343), .I2(x344), .O(n3263));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3264 (.I0(x333), .I1(x334), .I2(x335), .I3(n3260), .I4(n3261), .O(n3264));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3265 (.I0(x339), .I1(x340), .I2(x341), .I3(n3263), .I4(n3264), .O(n3265));
  LUT3 #(.INIT(8'h96)) lut_n3266 (.I0(n3250), .I1(n3253), .I2(n3254), .O(n3266));
  LUT3 #(.INIT(8'hE8)) lut_n3267 (.I0(n3262), .I1(n3265), .I2(n3266), .O(n3267));
  LUT3 #(.INIT(8'hE8)) lut_n3268 (.I0(x348), .I1(x349), .I2(x350), .O(n3268));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3269 (.I0(x339), .I1(x340), .I2(x341), .I3(n3263), .I4(n3264), .O(n3269));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3270 (.I0(x345), .I1(x346), .I2(x347), .I3(n3268), .I4(n3269), .O(n3270));
  LUT3 #(.INIT(8'hE8)) lut_n3271 (.I0(x354), .I1(x355), .I2(x356), .O(n3271));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3272 (.I0(x345), .I1(x346), .I2(x347), .I3(n3268), .I4(n3269), .O(n3272));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3273 (.I0(x351), .I1(x352), .I2(x353), .I3(n3271), .I4(n3272), .O(n3273));
  LUT3 #(.INIT(8'h96)) lut_n3274 (.I0(n3262), .I1(n3265), .I2(n3266), .O(n3274));
  LUT3 #(.INIT(8'hE8)) lut_n3275 (.I0(n3270), .I1(n3273), .I2(n3274), .O(n3275));
  LUT3 #(.INIT(8'h96)) lut_n3276 (.I0(n3247), .I1(n3255), .I2(n3256), .O(n3276));
  LUT3 #(.INIT(8'hE8)) lut_n3277 (.I0(n3267), .I1(n3275), .I2(n3276), .O(n3277));
  LUT3 #(.INIT(8'hE8)) lut_n3278 (.I0(x360), .I1(x361), .I2(x362), .O(n3278));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3279 (.I0(x351), .I1(x352), .I2(x353), .I3(n3271), .I4(n3272), .O(n3279));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3280 (.I0(x357), .I1(x358), .I2(x359), .I3(n3278), .I4(n3279), .O(n3280));
  LUT3 #(.INIT(8'hE8)) lut_n3281 (.I0(x366), .I1(x367), .I2(x368), .O(n3281));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3282 (.I0(x357), .I1(x358), .I2(x359), .I3(n3278), .I4(n3279), .O(n3282));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3283 (.I0(x363), .I1(x364), .I2(x365), .I3(n3281), .I4(n3282), .O(n3283));
  LUT3 #(.INIT(8'h96)) lut_n3284 (.I0(n3270), .I1(n3273), .I2(n3274), .O(n3284));
  LUT3 #(.INIT(8'hE8)) lut_n3285 (.I0(n3280), .I1(n3283), .I2(n3284), .O(n3285));
  LUT3 #(.INIT(8'hE8)) lut_n3286 (.I0(x372), .I1(x373), .I2(x374), .O(n3286));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3287 (.I0(x363), .I1(x364), .I2(x365), .I3(n3281), .I4(n3282), .O(n3287));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3288 (.I0(x369), .I1(x370), .I2(x371), .I3(n3286), .I4(n3287), .O(n3288));
  LUT3 #(.INIT(8'hE8)) lut_n3289 (.I0(x378), .I1(x379), .I2(x380), .O(n3289));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3290 (.I0(x369), .I1(x370), .I2(x371), .I3(n3286), .I4(n3287), .O(n3290));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3291 (.I0(x375), .I1(x376), .I2(x377), .I3(n3289), .I4(n3290), .O(n3291));
  LUT3 #(.INIT(8'h96)) lut_n3292 (.I0(n3280), .I1(n3283), .I2(n3284), .O(n3292));
  LUT3 #(.INIT(8'hE8)) lut_n3293 (.I0(n3288), .I1(n3291), .I2(n3292), .O(n3293));
  LUT3 #(.INIT(8'h96)) lut_n3294 (.I0(n3267), .I1(n3275), .I2(n3276), .O(n3294));
  LUT3 #(.INIT(8'hE8)) lut_n3295 (.I0(n3285), .I1(n3293), .I2(n3294), .O(n3295));
  LUT3 #(.INIT(8'h96)) lut_n3296 (.I0(n3239), .I1(n3257), .I2(n3258), .O(n3296));
  LUT3 #(.INIT(8'hE8)) lut_n3297 (.I0(n3277), .I1(n3295), .I2(n3296), .O(n3297));
  LUT3 #(.INIT(8'h96)) lut_n3298 (.I0(n3181), .I1(n3219), .I2(n3220), .O(n3298));
  LUT3 #(.INIT(8'hE8)) lut_n3299 (.I0(n3259), .I1(n3297), .I2(n3298), .O(n3299));
  LUT3 #(.INIT(8'hE8)) lut_n3300 (.I0(n3143), .I1(n3221), .I2(n3299), .O(n3300));
  LUT3 #(.INIT(8'hE8)) lut_n3301 (.I0(x384), .I1(x385), .I2(x386), .O(n3301));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3302 (.I0(x375), .I1(x376), .I2(x377), .I3(n3289), .I4(n3290), .O(n3302));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3303 (.I0(x381), .I1(x382), .I2(x383), .I3(n3301), .I4(n3302), .O(n3303));
  LUT3 #(.INIT(8'hE8)) lut_n3304 (.I0(x390), .I1(x391), .I2(x392), .O(n3304));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3305 (.I0(x381), .I1(x382), .I2(x383), .I3(n3301), .I4(n3302), .O(n3305));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3306 (.I0(x387), .I1(x388), .I2(x389), .I3(n3304), .I4(n3305), .O(n3306));
  LUT3 #(.INIT(8'h96)) lut_n3307 (.I0(n3288), .I1(n3291), .I2(n3292), .O(n3307));
  LUT3 #(.INIT(8'hE8)) lut_n3308 (.I0(n3303), .I1(n3306), .I2(n3307), .O(n3308));
  LUT3 #(.INIT(8'hE8)) lut_n3309 (.I0(x396), .I1(x397), .I2(x398), .O(n3309));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3310 (.I0(x387), .I1(x388), .I2(x389), .I3(n3304), .I4(n3305), .O(n3310));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3311 (.I0(x393), .I1(x394), .I2(x395), .I3(n3309), .I4(n3310), .O(n3311));
  LUT3 #(.INIT(8'hE8)) lut_n3312 (.I0(x402), .I1(x403), .I2(x404), .O(n3312));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3313 (.I0(x393), .I1(x394), .I2(x395), .I3(n3309), .I4(n3310), .O(n3313));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3314 (.I0(x399), .I1(x400), .I2(x401), .I3(n3312), .I4(n3313), .O(n3314));
  LUT3 #(.INIT(8'h96)) lut_n3315 (.I0(n3303), .I1(n3306), .I2(n3307), .O(n3315));
  LUT3 #(.INIT(8'hE8)) lut_n3316 (.I0(n3311), .I1(n3314), .I2(n3315), .O(n3316));
  LUT3 #(.INIT(8'h96)) lut_n3317 (.I0(n3285), .I1(n3293), .I2(n3294), .O(n3317));
  LUT3 #(.INIT(8'hE8)) lut_n3318 (.I0(n3308), .I1(n3316), .I2(n3317), .O(n3318));
  LUT3 #(.INIT(8'hE8)) lut_n3319 (.I0(x408), .I1(x409), .I2(x410), .O(n3319));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3320 (.I0(x399), .I1(x400), .I2(x401), .I3(n3312), .I4(n3313), .O(n3320));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3321 (.I0(x405), .I1(x406), .I2(x407), .I3(n3319), .I4(n3320), .O(n3321));
  LUT3 #(.INIT(8'hE8)) lut_n3322 (.I0(x414), .I1(x415), .I2(x416), .O(n3322));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3323 (.I0(x405), .I1(x406), .I2(x407), .I3(n3319), .I4(n3320), .O(n3323));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3324 (.I0(x411), .I1(x412), .I2(x413), .I3(n3322), .I4(n3323), .O(n3324));
  LUT3 #(.INIT(8'h96)) lut_n3325 (.I0(n3311), .I1(n3314), .I2(n3315), .O(n3325));
  LUT3 #(.INIT(8'hE8)) lut_n3326 (.I0(n3321), .I1(n3324), .I2(n3325), .O(n3326));
  LUT3 #(.INIT(8'hE8)) lut_n3327 (.I0(x420), .I1(x421), .I2(x422), .O(n3327));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3328 (.I0(x411), .I1(x412), .I2(x413), .I3(n3322), .I4(n3323), .O(n3328));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3329 (.I0(x417), .I1(x418), .I2(x419), .I3(n3327), .I4(n3328), .O(n3329));
  LUT3 #(.INIT(8'hE8)) lut_n3330 (.I0(x426), .I1(x427), .I2(x428), .O(n3330));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3331 (.I0(x417), .I1(x418), .I2(x419), .I3(n3327), .I4(n3328), .O(n3331));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3332 (.I0(x423), .I1(x424), .I2(x425), .I3(n3330), .I4(n3331), .O(n3332));
  LUT3 #(.INIT(8'h96)) lut_n3333 (.I0(n3321), .I1(n3324), .I2(n3325), .O(n3333));
  LUT3 #(.INIT(8'hE8)) lut_n3334 (.I0(n3329), .I1(n3332), .I2(n3333), .O(n3334));
  LUT3 #(.INIT(8'h96)) lut_n3335 (.I0(n3308), .I1(n3316), .I2(n3317), .O(n3335));
  LUT3 #(.INIT(8'hE8)) lut_n3336 (.I0(n3326), .I1(n3334), .I2(n3335), .O(n3336));
  LUT3 #(.INIT(8'h96)) lut_n3337 (.I0(n3277), .I1(n3295), .I2(n3296), .O(n3337));
  LUT3 #(.INIT(8'hE8)) lut_n3338 (.I0(n3318), .I1(n3336), .I2(n3337), .O(n3338));
  LUT3 #(.INIT(8'hE8)) lut_n3339 (.I0(x432), .I1(x433), .I2(x434), .O(n3339));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3340 (.I0(x423), .I1(x424), .I2(x425), .I3(n3330), .I4(n3331), .O(n3340));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3341 (.I0(x429), .I1(x430), .I2(x431), .I3(n3339), .I4(n3340), .O(n3341));
  LUT3 #(.INIT(8'hE8)) lut_n3342 (.I0(x438), .I1(x439), .I2(x440), .O(n3342));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3343 (.I0(x429), .I1(x430), .I2(x431), .I3(n3339), .I4(n3340), .O(n3343));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3344 (.I0(x435), .I1(x436), .I2(x437), .I3(n3342), .I4(n3343), .O(n3344));
  LUT3 #(.INIT(8'h96)) lut_n3345 (.I0(n3329), .I1(n3332), .I2(n3333), .O(n3345));
  LUT3 #(.INIT(8'hE8)) lut_n3346 (.I0(n3341), .I1(n3344), .I2(n3345), .O(n3346));
  LUT3 #(.INIT(8'hE8)) lut_n3347 (.I0(x444), .I1(x445), .I2(x446), .O(n3347));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3348 (.I0(x435), .I1(x436), .I2(x437), .I3(n3342), .I4(n3343), .O(n3348));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3349 (.I0(x441), .I1(x442), .I2(x443), .I3(n3347), .I4(n3348), .O(n3349));
  LUT3 #(.INIT(8'hE8)) lut_n3350 (.I0(x450), .I1(x451), .I2(x452), .O(n3350));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3351 (.I0(x441), .I1(x442), .I2(x443), .I3(n3347), .I4(n3348), .O(n3351));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3352 (.I0(x447), .I1(x448), .I2(x449), .I3(n3350), .I4(n3351), .O(n3352));
  LUT3 #(.INIT(8'h96)) lut_n3353 (.I0(n3341), .I1(n3344), .I2(n3345), .O(n3353));
  LUT3 #(.INIT(8'hE8)) lut_n3354 (.I0(n3349), .I1(n3352), .I2(n3353), .O(n3354));
  LUT3 #(.INIT(8'h96)) lut_n3355 (.I0(n3326), .I1(n3334), .I2(n3335), .O(n3355));
  LUT3 #(.INIT(8'hE8)) lut_n3356 (.I0(n3346), .I1(n3354), .I2(n3355), .O(n3356));
  LUT3 #(.INIT(8'hE8)) lut_n3357 (.I0(x456), .I1(x457), .I2(x458), .O(n3357));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3358 (.I0(x447), .I1(x448), .I2(x449), .I3(n3350), .I4(n3351), .O(n3358));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3359 (.I0(x453), .I1(x454), .I2(x455), .I3(n3357), .I4(n3358), .O(n3359));
  LUT3 #(.INIT(8'hE8)) lut_n3360 (.I0(x462), .I1(x463), .I2(x464), .O(n3360));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3361 (.I0(x453), .I1(x454), .I2(x455), .I3(n3357), .I4(n3358), .O(n3361));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3362 (.I0(x459), .I1(x460), .I2(x461), .I3(n3360), .I4(n3361), .O(n3362));
  LUT3 #(.INIT(8'h96)) lut_n3363 (.I0(n3349), .I1(n3352), .I2(n3353), .O(n3363));
  LUT3 #(.INIT(8'hE8)) lut_n3364 (.I0(n3359), .I1(n3362), .I2(n3363), .O(n3364));
  LUT3 #(.INIT(8'hE8)) lut_n3365 (.I0(x468), .I1(x469), .I2(x470), .O(n3365));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3366 (.I0(x459), .I1(x460), .I2(x461), .I3(n3360), .I4(n3361), .O(n3366));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3367 (.I0(x465), .I1(x466), .I2(x467), .I3(n3365), .I4(n3366), .O(n3367));
  LUT3 #(.INIT(8'hE8)) lut_n3368 (.I0(x474), .I1(x475), .I2(x476), .O(n3368));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3369 (.I0(x465), .I1(x466), .I2(x467), .I3(n3365), .I4(n3366), .O(n3369));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3370 (.I0(x471), .I1(x472), .I2(x473), .I3(n3368), .I4(n3369), .O(n3370));
  LUT3 #(.INIT(8'h96)) lut_n3371 (.I0(n3359), .I1(n3362), .I2(n3363), .O(n3371));
  LUT3 #(.INIT(8'hE8)) lut_n3372 (.I0(n3367), .I1(n3370), .I2(n3371), .O(n3372));
  LUT3 #(.INIT(8'h96)) lut_n3373 (.I0(n3346), .I1(n3354), .I2(n3355), .O(n3373));
  LUT3 #(.INIT(8'hE8)) lut_n3374 (.I0(n3364), .I1(n3372), .I2(n3373), .O(n3374));
  LUT3 #(.INIT(8'h96)) lut_n3375 (.I0(n3318), .I1(n3336), .I2(n3337), .O(n3375));
  LUT3 #(.INIT(8'hE8)) lut_n3376 (.I0(n3356), .I1(n3374), .I2(n3375), .O(n3376));
  LUT3 #(.INIT(8'h96)) lut_n3377 (.I0(n3259), .I1(n3297), .I2(n3298), .O(n3377));
  LUT3 #(.INIT(8'hE8)) lut_n3378 (.I0(n3338), .I1(n3376), .I2(n3377), .O(n3378));
  LUT3 #(.INIT(8'hE8)) lut_n3379 (.I0(x480), .I1(x481), .I2(x482), .O(n3379));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3380 (.I0(x471), .I1(x472), .I2(x473), .I3(n3368), .I4(n3369), .O(n3380));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3381 (.I0(x477), .I1(x478), .I2(x479), .I3(n3379), .I4(n3380), .O(n3381));
  LUT3 #(.INIT(8'hE8)) lut_n3382 (.I0(x486), .I1(x487), .I2(x488), .O(n3382));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3383 (.I0(x477), .I1(x478), .I2(x479), .I3(n3379), .I4(n3380), .O(n3383));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3384 (.I0(x483), .I1(x484), .I2(x485), .I3(n3382), .I4(n3383), .O(n3384));
  LUT3 #(.INIT(8'h96)) lut_n3385 (.I0(n3367), .I1(n3370), .I2(n3371), .O(n3385));
  LUT3 #(.INIT(8'hE8)) lut_n3386 (.I0(n3381), .I1(n3384), .I2(n3385), .O(n3386));
  LUT3 #(.INIT(8'hE8)) lut_n3387 (.I0(x492), .I1(x493), .I2(x494), .O(n3387));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3388 (.I0(x483), .I1(x484), .I2(x485), .I3(n3382), .I4(n3383), .O(n3388));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3389 (.I0(x489), .I1(x490), .I2(x491), .I3(n3387), .I4(n3388), .O(n3389));
  LUT3 #(.INIT(8'hE8)) lut_n3390 (.I0(x498), .I1(x499), .I2(x500), .O(n3390));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3391 (.I0(x489), .I1(x490), .I2(x491), .I3(n3387), .I4(n3388), .O(n3391));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3392 (.I0(x495), .I1(x496), .I2(x497), .I3(n3390), .I4(n3391), .O(n3392));
  LUT3 #(.INIT(8'h96)) lut_n3393 (.I0(n3381), .I1(n3384), .I2(n3385), .O(n3393));
  LUT3 #(.INIT(8'hE8)) lut_n3394 (.I0(n3389), .I1(n3392), .I2(n3393), .O(n3394));
  LUT3 #(.INIT(8'h96)) lut_n3395 (.I0(n3364), .I1(n3372), .I2(n3373), .O(n3395));
  LUT3 #(.INIT(8'hE8)) lut_n3396 (.I0(n3386), .I1(n3394), .I2(n3395), .O(n3396));
  LUT3 #(.INIT(8'hE8)) lut_n3397 (.I0(x504), .I1(x505), .I2(x506), .O(n3397));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3398 (.I0(x495), .I1(x496), .I2(x497), .I3(n3390), .I4(n3391), .O(n3398));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3399 (.I0(x501), .I1(x502), .I2(x503), .I3(n3397), .I4(n3398), .O(n3399));
  LUT3 #(.INIT(8'hE8)) lut_n3400 (.I0(x510), .I1(x511), .I2(x512), .O(n3400));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3401 (.I0(x501), .I1(x502), .I2(x503), .I3(n3397), .I4(n3398), .O(n3401));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3402 (.I0(x507), .I1(x508), .I2(x509), .I3(n3400), .I4(n3401), .O(n3402));
  LUT3 #(.INIT(8'h96)) lut_n3403 (.I0(n3389), .I1(n3392), .I2(n3393), .O(n3403));
  LUT3 #(.INIT(8'hE8)) lut_n3404 (.I0(n3399), .I1(n3402), .I2(n3403), .O(n3404));
  LUT3 #(.INIT(8'hE8)) lut_n3405 (.I0(x516), .I1(x517), .I2(x518), .O(n3405));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3406 (.I0(x507), .I1(x508), .I2(x509), .I3(n3400), .I4(n3401), .O(n3406));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3407 (.I0(x513), .I1(x514), .I2(x515), .I3(n3405), .I4(n3406), .O(n3407));
  LUT3 #(.INIT(8'hE8)) lut_n3408 (.I0(x522), .I1(x523), .I2(x524), .O(n3408));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3409 (.I0(x513), .I1(x514), .I2(x515), .I3(n3405), .I4(n3406), .O(n3409));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3410 (.I0(x519), .I1(x520), .I2(x521), .I3(n3408), .I4(n3409), .O(n3410));
  LUT3 #(.INIT(8'h96)) lut_n3411 (.I0(n3399), .I1(n3402), .I2(n3403), .O(n3411));
  LUT3 #(.INIT(8'hE8)) lut_n3412 (.I0(n3407), .I1(n3410), .I2(n3411), .O(n3412));
  LUT3 #(.INIT(8'h96)) lut_n3413 (.I0(n3386), .I1(n3394), .I2(n3395), .O(n3413));
  LUT3 #(.INIT(8'hE8)) lut_n3414 (.I0(n3404), .I1(n3412), .I2(n3413), .O(n3414));
  LUT3 #(.INIT(8'h96)) lut_n3415 (.I0(n3356), .I1(n3374), .I2(n3375), .O(n3415));
  LUT3 #(.INIT(8'hE8)) lut_n3416 (.I0(n3396), .I1(n3414), .I2(n3415), .O(n3416));
  LUT3 #(.INIT(8'hE8)) lut_n3417 (.I0(x528), .I1(x529), .I2(x530), .O(n3417));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3418 (.I0(x519), .I1(x520), .I2(x521), .I3(n3408), .I4(n3409), .O(n3418));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3419 (.I0(x525), .I1(x526), .I2(x527), .I3(n3417), .I4(n3418), .O(n3419));
  LUT3 #(.INIT(8'hE8)) lut_n3420 (.I0(x534), .I1(x535), .I2(x536), .O(n3420));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3421 (.I0(x525), .I1(x526), .I2(x527), .I3(n3417), .I4(n3418), .O(n3421));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3422 (.I0(x531), .I1(x532), .I2(x533), .I3(n3420), .I4(n3421), .O(n3422));
  LUT3 #(.INIT(8'h96)) lut_n3423 (.I0(n3407), .I1(n3410), .I2(n3411), .O(n3423));
  LUT3 #(.INIT(8'hE8)) lut_n3424 (.I0(n3419), .I1(n3422), .I2(n3423), .O(n3424));
  LUT3 #(.INIT(8'hE8)) lut_n3425 (.I0(x540), .I1(x541), .I2(x542), .O(n3425));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3426 (.I0(x531), .I1(x532), .I2(x533), .I3(n3420), .I4(n3421), .O(n3426));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3427 (.I0(x537), .I1(x538), .I2(x539), .I3(n3425), .I4(n3426), .O(n3427));
  LUT3 #(.INIT(8'hE8)) lut_n3428 (.I0(x546), .I1(x547), .I2(x548), .O(n3428));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3429 (.I0(x537), .I1(x538), .I2(x539), .I3(n3425), .I4(n3426), .O(n3429));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3430 (.I0(x543), .I1(x544), .I2(x545), .I3(n3428), .I4(n3429), .O(n3430));
  LUT3 #(.INIT(8'h96)) lut_n3431 (.I0(n3419), .I1(n3422), .I2(n3423), .O(n3431));
  LUT3 #(.INIT(8'hE8)) lut_n3432 (.I0(n3427), .I1(n3430), .I2(n3431), .O(n3432));
  LUT3 #(.INIT(8'h96)) lut_n3433 (.I0(n3404), .I1(n3412), .I2(n3413), .O(n3433));
  LUT3 #(.INIT(8'hE8)) lut_n3434 (.I0(n3424), .I1(n3432), .I2(n3433), .O(n3434));
  LUT3 #(.INIT(8'hE8)) lut_n3435 (.I0(x552), .I1(x553), .I2(x554), .O(n3435));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3436 (.I0(x543), .I1(x544), .I2(x545), .I3(n3428), .I4(n3429), .O(n3436));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3437 (.I0(x549), .I1(x550), .I2(x551), .I3(n3435), .I4(n3436), .O(n3437));
  LUT3 #(.INIT(8'hE8)) lut_n3438 (.I0(x558), .I1(x559), .I2(x560), .O(n3438));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3439 (.I0(x549), .I1(x550), .I2(x551), .I3(n3435), .I4(n3436), .O(n3439));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3440 (.I0(x555), .I1(x556), .I2(x557), .I3(n3438), .I4(n3439), .O(n3440));
  LUT3 #(.INIT(8'h96)) lut_n3441 (.I0(n3427), .I1(n3430), .I2(n3431), .O(n3441));
  LUT3 #(.INIT(8'hE8)) lut_n3442 (.I0(n3437), .I1(n3440), .I2(n3441), .O(n3442));
  LUT3 #(.INIT(8'hE8)) lut_n3443 (.I0(x564), .I1(x565), .I2(x566), .O(n3443));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3444 (.I0(x555), .I1(x556), .I2(x557), .I3(n3438), .I4(n3439), .O(n3444));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3445 (.I0(x561), .I1(x562), .I2(x563), .I3(n3443), .I4(n3444), .O(n3445));
  LUT3 #(.INIT(8'hE8)) lut_n3446 (.I0(x570), .I1(x571), .I2(x572), .O(n3446));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3447 (.I0(x561), .I1(x562), .I2(x563), .I3(n3443), .I4(n3444), .O(n3447));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3448 (.I0(x567), .I1(x568), .I2(x569), .I3(n3446), .I4(n3447), .O(n3448));
  LUT3 #(.INIT(8'h96)) lut_n3449 (.I0(n3437), .I1(n3440), .I2(n3441), .O(n3449));
  LUT3 #(.INIT(8'hE8)) lut_n3450 (.I0(n3445), .I1(n3448), .I2(n3449), .O(n3450));
  LUT3 #(.INIT(8'h96)) lut_n3451 (.I0(n3424), .I1(n3432), .I2(n3433), .O(n3451));
  LUT3 #(.INIT(8'hE8)) lut_n3452 (.I0(n3442), .I1(n3450), .I2(n3451), .O(n3452));
  LUT3 #(.INIT(8'h96)) lut_n3453 (.I0(n3396), .I1(n3414), .I2(n3415), .O(n3453));
  LUT3 #(.INIT(8'hE8)) lut_n3454 (.I0(n3434), .I1(n3452), .I2(n3453), .O(n3454));
  LUT3 #(.INIT(8'h96)) lut_n3455 (.I0(n3338), .I1(n3376), .I2(n3377), .O(n3455));
  LUT3 #(.INIT(8'hE8)) lut_n3456 (.I0(n3416), .I1(n3454), .I2(n3455), .O(n3456));
  LUT3 #(.INIT(8'h96)) lut_n3457 (.I0(n3143), .I1(n3221), .I2(n3299), .O(n3457));
  LUT3 #(.INIT(8'hE8)) lut_n3458 (.I0(n3378), .I1(n3456), .I2(n3457), .O(n3458));
  LUT3 #(.INIT(8'hE8)) lut_n3459 (.I0(x576), .I1(x577), .I2(x578), .O(n3459));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3460 (.I0(x567), .I1(x568), .I2(x569), .I3(n3446), .I4(n3447), .O(n3460));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3461 (.I0(x573), .I1(x574), .I2(x575), .I3(n3459), .I4(n3460), .O(n3461));
  LUT3 #(.INIT(8'hE8)) lut_n3462 (.I0(x582), .I1(x583), .I2(x584), .O(n3462));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3463 (.I0(x573), .I1(x574), .I2(x575), .I3(n3459), .I4(n3460), .O(n3463));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3464 (.I0(x579), .I1(x580), .I2(x581), .I3(n3462), .I4(n3463), .O(n3464));
  LUT3 #(.INIT(8'h96)) lut_n3465 (.I0(n3445), .I1(n3448), .I2(n3449), .O(n3465));
  LUT3 #(.INIT(8'hE8)) lut_n3466 (.I0(n3461), .I1(n3464), .I2(n3465), .O(n3466));
  LUT3 #(.INIT(8'hE8)) lut_n3467 (.I0(x588), .I1(x589), .I2(x590), .O(n3467));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3468 (.I0(x579), .I1(x580), .I2(x581), .I3(n3462), .I4(n3463), .O(n3468));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3469 (.I0(x585), .I1(x586), .I2(x587), .I3(n3467), .I4(n3468), .O(n3469));
  LUT3 #(.INIT(8'hE8)) lut_n3470 (.I0(x594), .I1(x595), .I2(x596), .O(n3470));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3471 (.I0(x585), .I1(x586), .I2(x587), .I3(n3467), .I4(n3468), .O(n3471));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3472 (.I0(x591), .I1(x592), .I2(x593), .I3(n3470), .I4(n3471), .O(n3472));
  LUT3 #(.INIT(8'h96)) lut_n3473 (.I0(n3461), .I1(n3464), .I2(n3465), .O(n3473));
  LUT3 #(.INIT(8'hE8)) lut_n3474 (.I0(n3469), .I1(n3472), .I2(n3473), .O(n3474));
  LUT3 #(.INIT(8'h96)) lut_n3475 (.I0(n3442), .I1(n3450), .I2(n3451), .O(n3475));
  LUT3 #(.INIT(8'hE8)) lut_n3476 (.I0(n3466), .I1(n3474), .I2(n3475), .O(n3476));
  LUT3 #(.INIT(8'hE8)) lut_n3477 (.I0(x600), .I1(x601), .I2(x602), .O(n3477));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3478 (.I0(x591), .I1(x592), .I2(x593), .I3(n3470), .I4(n3471), .O(n3478));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3479 (.I0(x597), .I1(x598), .I2(x599), .I3(n3477), .I4(n3478), .O(n3479));
  LUT3 #(.INIT(8'hE8)) lut_n3480 (.I0(x606), .I1(x607), .I2(x608), .O(n3480));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3481 (.I0(x597), .I1(x598), .I2(x599), .I3(n3477), .I4(n3478), .O(n3481));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3482 (.I0(x603), .I1(x604), .I2(x605), .I3(n3480), .I4(n3481), .O(n3482));
  LUT3 #(.INIT(8'h96)) lut_n3483 (.I0(n3469), .I1(n3472), .I2(n3473), .O(n3483));
  LUT3 #(.INIT(8'hE8)) lut_n3484 (.I0(n3479), .I1(n3482), .I2(n3483), .O(n3484));
  LUT3 #(.INIT(8'hE8)) lut_n3485 (.I0(x612), .I1(x613), .I2(x614), .O(n3485));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3486 (.I0(x603), .I1(x604), .I2(x605), .I3(n3480), .I4(n3481), .O(n3486));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3487 (.I0(x609), .I1(x610), .I2(x611), .I3(n3485), .I4(n3486), .O(n3487));
  LUT3 #(.INIT(8'hE8)) lut_n3488 (.I0(x618), .I1(x619), .I2(x620), .O(n3488));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3489 (.I0(x609), .I1(x610), .I2(x611), .I3(n3485), .I4(n3486), .O(n3489));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3490 (.I0(x615), .I1(x616), .I2(x617), .I3(n3488), .I4(n3489), .O(n3490));
  LUT3 #(.INIT(8'h96)) lut_n3491 (.I0(n3479), .I1(n3482), .I2(n3483), .O(n3491));
  LUT3 #(.INIT(8'hE8)) lut_n3492 (.I0(n3487), .I1(n3490), .I2(n3491), .O(n3492));
  LUT3 #(.INIT(8'h96)) lut_n3493 (.I0(n3466), .I1(n3474), .I2(n3475), .O(n3493));
  LUT3 #(.INIT(8'hE8)) lut_n3494 (.I0(n3484), .I1(n3492), .I2(n3493), .O(n3494));
  LUT3 #(.INIT(8'h96)) lut_n3495 (.I0(n3434), .I1(n3452), .I2(n3453), .O(n3495));
  LUT3 #(.INIT(8'hE8)) lut_n3496 (.I0(n3476), .I1(n3494), .I2(n3495), .O(n3496));
  LUT3 #(.INIT(8'hE8)) lut_n3497 (.I0(x624), .I1(x625), .I2(x626), .O(n3497));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3498 (.I0(x615), .I1(x616), .I2(x617), .I3(n3488), .I4(n3489), .O(n3498));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3499 (.I0(x621), .I1(x622), .I2(x623), .I3(n3497), .I4(n3498), .O(n3499));
  LUT3 #(.INIT(8'hE8)) lut_n3500 (.I0(x630), .I1(x631), .I2(x632), .O(n3500));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3501 (.I0(x621), .I1(x622), .I2(x623), .I3(n3497), .I4(n3498), .O(n3501));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3502 (.I0(x627), .I1(x628), .I2(x629), .I3(n3500), .I4(n3501), .O(n3502));
  LUT3 #(.INIT(8'h96)) lut_n3503 (.I0(n3487), .I1(n3490), .I2(n3491), .O(n3503));
  LUT3 #(.INIT(8'hE8)) lut_n3504 (.I0(n3499), .I1(n3502), .I2(n3503), .O(n3504));
  LUT3 #(.INIT(8'hE8)) lut_n3505 (.I0(x636), .I1(x637), .I2(x638), .O(n3505));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3506 (.I0(x627), .I1(x628), .I2(x629), .I3(n3500), .I4(n3501), .O(n3506));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3507 (.I0(x633), .I1(x634), .I2(x635), .I3(n3505), .I4(n3506), .O(n3507));
  LUT3 #(.INIT(8'hE8)) lut_n3508 (.I0(x642), .I1(x643), .I2(x644), .O(n3508));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3509 (.I0(x633), .I1(x634), .I2(x635), .I3(n3505), .I4(n3506), .O(n3509));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3510 (.I0(x639), .I1(x640), .I2(x641), .I3(n3508), .I4(n3509), .O(n3510));
  LUT3 #(.INIT(8'h96)) lut_n3511 (.I0(n3499), .I1(n3502), .I2(n3503), .O(n3511));
  LUT3 #(.INIT(8'hE8)) lut_n3512 (.I0(n3507), .I1(n3510), .I2(n3511), .O(n3512));
  LUT3 #(.INIT(8'h96)) lut_n3513 (.I0(n3484), .I1(n3492), .I2(n3493), .O(n3513));
  LUT3 #(.INIT(8'hE8)) lut_n3514 (.I0(n3504), .I1(n3512), .I2(n3513), .O(n3514));
  LUT3 #(.INIT(8'hE8)) lut_n3515 (.I0(x648), .I1(x649), .I2(x650), .O(n3515));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3516 (.I0(x639), .I1(x640), .I2(x641), .I3(n3508), .I4(n3509), .O(n3516));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3517 (.I0(x645), .I1(x646), .I2(x647), .I3(n3515), .I4(n3516), .O(n3517));
  LUT3 #(.INIT(8'hE8)) lut_n3518 (.I0(x654), .I1(x655), .I2(x656), .O(n3518));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3519 (.I0(x645), .I1(x646), .I2(x647), .I3(n3515), .I4(n3516), .O(n3519));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3520 (.I0(x651), .I1(x652), .I2(x653), .I3(n3518), .I4(n3519), .O(n3520));
  LUT3 #(.INIT(8'h96)) lut_n3521 (.I0(n3507), .I1(n3510), .I2(n3511), .O(n3521));
  LUT3 #(.INIT(8'hE8)) lut_n3522 (.I0(n3517), .I1(n3520), .I2(n3521), .O(n3522));
  LUT3 #(.INIT(8'hE8)) lut_n3523 (.I0(x660), .I1(x661), .I2(x662), .O(n3523));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3524 (.I0(x651), .I1(x652), .I2(x653), .I3(n3518), .I4(n3519), .O(n3524));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3525 (.I0(x657), .I1(x658), .I2(x659), .I3(n3523), .I4(n3524), .O(n3525));
  LUT3 #(.INIT(8'hE8)) lut_n3526 (.I0(x666), .I1(x667), .I2(x668), .O(n3526));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3527 (.I0(x657), .I1(x658), .I2(x659), .I3(n3523), .I4(n3524), .O(n3527));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3528 (.I0(x663), .I1(x664), .I2(x665), .I3(n3526), .I4(n3527), .O(n3528));
  LUT3 #(.INIT(8'h96)) lut_n3529 (.I0(n3517), .I1(n3520), .I2(n3521), .O(n3529));
  LUT3 #(.INIT(8'hE8)) lut_n3530 (.I0(n3525), .I1(n3528), .I2(n3529), .O(n3530));
  LUT3 #(.INIT(8'h96)) lut_n3531 (.I0(n3504), .I1(n3512), .I2(n3513), .O(n3531));
  LUT3 #(.INIT(8'hE8)) lut_n3532 (.I0(n3522), .I1(n3530), .I2(n3531), .O(n3532));
  LUT3 #(.INIT(8'h96)) lut_n3533 (.I0(n3476), .I1(n3494), .I2(n3495), .O(n3533));
  LUT3 #(.INIT(8'hE8)) lut_n3534 (.I0(n3514), .I1(n3532), .I2(n3533), .O(n3534));
  LUT3 #(.INIT(8'h96)) lut_n3535 (.I0(n3416), .I1(n3454), .I2(n3455), .O(n3535));
  LUT3 #(.INIT(8'hE8)) lut_n3536 (.I0(n3496), .I1(n3534), .I2(n3535), .O(n3536));
  LUT3 #(.INIT(8'hE8)) lut_n3537 (.I0(x672), .I1(x673), .I2(x674), .O(n3537));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3538 (.I0(x663), .I1(x664), .I2(x665), .I3(n3526), .I4(n3527), .O(n3538));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3539 (.I0(x669), .I1(x670), .I2(x671), .I3(n3537), .I4(n3538), .O(n3539));
  LUT3 #(.INIT(8'hE8)) lut_n3540 (.I0(x678), .I1(x679), .I2(x680), .O(n3540));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3541 (.I0(x669), .I1(x670), .I2(x671), .I3(n3537), .I4(n3538), .O(n3541));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3542 (.I0(x675), .I1(x676), .I2(x677), .I3(n3540), .I4(n3541), .O(n3542));
  LUT3 #(.INIT(8'h96)) lut_n3543 (.I0(n3525), .I1(n3528), .I2(n3529), .O(n3543));
  LUT3 #(.INIT(8'hE8)) lut_n3544 (.I0(n3539), .I1(n3542), .I2(n3543), .O(n3544));
  LUT3 #(.INIT(8'hE8)) lut_n3545 (.I0(x684), .I1(x685), .I2(x686), .O(n3545));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3546 (.I0(x675), .I1(x676), .I2(x677), .I3(n3540), .I4(n3541), .O(n3546));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3547 (.I0(x681), .I1(x682), .I2(x683), .I3(n3545), .I4(n3546), .O(n3547));
  LUT3 #(.INIT(8'hE8)) lut_n3548 (.I0(x690), .I1(x691), .I2(x692), .O(n3548));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3549 (.I0(x681), .I1(x682), .I2(x683), .I3(n3545), .I4(n3546), .O(n3549));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3550 (.I0(x687), .I1(x688), .I2(x689), .I3(n3548), .I4(n3549), .O(n3550));
  LUT3 #(.INIT(8'h96)) lut_n3551 (.I0(n3539), .I1(n3542), .I2(n3543), .O(n3551));
  LUT3 #(.INIT(8'hE8)) lut_n3552 (.I0(n3547), .I1(n3550), .I2(n3551), .O(n3552));
  LUT3 #(.INIT(8'h96)) lut_n3553 (.I0(n3522), .I1(n3530), .I2(n3531), .O(n3553));
  LUT3 #(.INIT(8'hE8)) lut_n3554 (.I0(n3544), .I1(n3552), .I2(n3553), .O(n3554));
  LUT3 #(.INIT(8'hE8)) lut_n3555 (.I0(x696), .I1(x697), .I2(x698), .O(n3555));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3556 (.I0(x687), .I1(x688), .I2(x689), .I3(n3548), .I4(n3549), .O(n3556));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3557 (.I0(x693), .I1(x694), .I2(x695), .I3(n3555), .I4(n3556), .O(n3557));
  LUT3 #(.INIT(8'hE8)) lut_n3558 (.I0(x702), .I1(x703), .I2(x704), .O(n3558));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3559 (.I0(x693), .I1(x694), .I2(x695), .I3(n3555), .I4(n3556), .O(n3559));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3560 (.I0(x699), .I1(x700), .I2(x701), .I3(n3558), .I4(n3559), .O(n3560));
  LUT3 #(.INIT(8'h96)) lut_n3561 (.I0(n3547), .I1(n3550), .I2(n3551), .O(n3561));
  LUT3 #(.INIT(8'hE8)) lut_n3562 (.I0(n3557), .I1(n3560), .I2(n3561), .O(n3562));
  LUT3 #(.INIT(8'hE8)) lut_n3563 (.I0(x708), .I1(x709), .I2(x710), .O(n3563));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3564 (.I0(x699), .I1(x700), .I2(x701), .I3(n3558), .I4(n3559), .O(n3564));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3565 (.I0(x705), .I1(x706), .I2(x707), .I3(n3563), .I4(n3564), .O(n3565));
  LUT3 #(.INIT(8'hE8)) lut_n3566 (.I0(x714), .I1(x715), .I2(x716), .O(n3566));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3567 (.I0(x705), .I1(x706), .I2(x707), .I3(n3563), .I4(n3564), .O(n3567));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3568 (.I0(x711), .I1(x712), .I2(x713), .I3(n3566), .I4(n3567), .O(n3568));
  LUT3 #(.INIT(8'h96)) lut_n3569 (.I0(n3557), .I1(n3560), .I2(n3561), .O(n3569));
  LUT3 #(.INIT(8'hE8)) lut_n3570 (.I0(n3565), .I1(n3568), .I2(n3569), .O(n3570));
  LUT3 #(.INIT(8'h96)) lut_n3571 (.I0(n3544), .I1(n3552), .I2(n3553), .O(n3571));
  LUT3 #(.INIT(8'hE8)) lut_n3572 (.I0(n3562), .I1(n3570), .I2(n3571), .O(n3572));
  LUT3 #(.INIT(8'h96)) lut_n3573 (.I0(n3514), .I1(n3532), .I2(n3533), .O(n3573));
  LUT3 #(.INIT(8'hE8)) lut_n3574 (.I0(n3554), .I1(n3572), .I2(n3573), .O(n3574));
  LUT3 #(.INIT(8'hE8)) lut_n3575 (.I0(x720), .I1(x721), .I2(x722), .O(n3575));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3576 (.I0(x711), .I1(x712), .I2(x713), .I3(n3566), .I4(n3567), .O(n3576));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3577 (.I0(x717), .I1(x718), .I2(x719), .I3(n3575), .I4(n3576), .O(n3577));
  LUT3 #(.INIT(8'hE8)) lut_n3578 (.I0(x726), .I1(x727), .I2(x728), .O(n3578));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3579 (.I0(x717), .I1(x718), .I2(x719), .I3(n3575), .I4(n3576), .O(n3579));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3580 (.I0(x723), .I1(x724), .I2(x725), .I3(n3578), .I4(n3579), .O(n3580));
  LUT3 #(.INIT(8'h96)) lut_n3581 (.I0(n3565), .I1(n3568), .I2(n3569), .O(n3581));
  LUT3 #(.INIT(8'hE8)) lut_n3582 (.I0(n3577), .I1(n3580), .I2(n3581), .O(n3582));
  LUT3 #(.INIT(8'hE8)) lut_n3583 (.I0(x732), .I1(x733), .I2(x734), .O(n3583));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3584 (.I0(x723), .I1(x724), .I2(x725), .I3(n3578), .I4(n3579), .O(n3584));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3585 (.I0(x729), .I1(x730), .I2(x731), .I3(n3583), .I4(n3584), .O(n3585));
  LUT3 #(.INIT(8'hE8)) lut_n3586 (.I0(x738), .I1(x739), .I2(x740), .O(n3586));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3587 (.I0(x729), .I1(x730), .I2(x731), .I3(n3583), .I4(n3584), .O(n3587));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3588 (.I0(x735), .I1(x736), .I2(x737), .I3(n3586), .I4(n3587), .O(n3588));
  LUT3 #(.INIT(8'h96)) lut_n3589 (.I0(n3577), .I1(n3580), .I2(n3581), .O(n3589));
  LUT3 #(.INIT(8'hE8)) lut_n3590 (.I0(n3585), .I1(n3588), .I2(n3589), .O(n3590));
  LUT3 #(.INIT(8'h96)) lut_n3591 (.I0(n3562), .I1(n3570), .I2(n3571), .O(n3591));
  LUT3 #(.INIT(8'hE8)) lut_n3592 (.I0(n3582), .I1(n3590), .I2(n3591), .O(n3592));
  LUT3 #(.INIT(8'hE8)) lut_n3593 (.I0(x744), .I1(x745), .I2(x746), .O(n3593));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3594 (.I0(x735), .I1(x736), .I2(x737), .I3(n3586), .I4(n3587), .O(n3594));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3595 (.I0(x741), .I1(x742), .I2(x743), .I3(n3593), .I4(n3594), .O(n3595));
  LUT3 #(.INIT(8'hE8)) lut_n3596 (.I0(x750), .I1(x751), .I2(x752), .O(n3596));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3597 (.I0(x741), .I1(x742), .I2(x743), .I3(n3593), .I4(n3594), .O(n3597));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3598 (.I0(x747), .I1(x748), .I2(x749), .I3(n3596), .I4(n3597), .O(n3598));
  LUT3 #(.INIT(8'h96)) lut_n3599 (.I0(n3585), .I1(n3588), .I2(n3589), .O(n3599));
  LUT3 #(.INIT(8'hE8)) lut_n3600 (.I0(n3595), .I1(n3598), .I2(n3599), .O(n3600));
  LUT3 #(.INIT(8'hE8)) lut_n3601 (.I0(x756), .I1(x757), .I2(x758), .O(n3601));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3602 (.I0(x747), .I1(x748), .I2(x749), .I3(n3596), .I4(n3597), .O(n3602));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3603 (.I0(x753), .I1(x754), .I2(x755), .I3(n3601), .I4(n3602), .O(n3603));
  LUT3 #(.INIT(8'hE8)) lut_n3604 (.I0(x762), .I1(x763), .I2(x764), .O(n3604));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3605 (.I0(x753), .I1(x754), .I2(x755), .I3(n3601), .I4(n3602), .O(n3605));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3606 (.I0(x759), .I1(x760), .I2(x761), .I3(n3604), .I4(n3605), .O(n3606));
  LUT3 #(.INIT(8'h96)) lut_n3607 (.I0(n3595), .I1(n3598), .I2(n3599), .O(n3607));
  LUT3 #(.INIT(8'hE8)) lut_n3608 (.I0(n3603), .I1(n3606), .I2(n3607), .O(n3608));
  LUT3 #(.INIT(8'h96)) lut_n3609 (.I0(n3582), .I1(n3590), .I2(n3591), .O(n3609));
  LUT3 #(.INIT(8'hE8)) lut_n3610 (.I0(n3600), .I1(n3608), .I2(n3609), .O(n3610));
  LUT3 #(.INIT(8'h96)) lut_n3611 (.I0(n3554), .I1(n3572), .I2(n3573), .O(n3611));
  LUT3 #(.INIT(8'hE8)) lut_n3612 (.I0(n3592), .I1(n3610), .I2(n3611), .O(n3612));
  LUT3 #(.INIT(8'h96)) lut_n3613 (.I0(n3496), .I1(n3534), .I2(n3535), .O(n3613));
  LUT3 #(.INIT(8'hE8)) lut_n3614 (.I0(n3574), .I1(n3612), .I2(n3613), .O(n3614));
  LUT3 #(.INIT(8'h96)) lut_n3615 (.I0(n3378), .I1(n3456), .I2(n3457), .O(n3615));
  LUT3 #(.INIT(8'hE8)) lut_n3616 (.I0(n3536), .I1(n3614), .I2(n3615), .O(n3616));
  LUT3 #(.INIT(8'hE8)) lut_n3617 (.I0(n3300), .I1(n3458), .I2(n3616), .O(n3617));
  LUT3 #(.INIT(8'hE8)) lut_n3618 (.I0(x768), .I1(x769), .I2(x770), .O(n3618));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3619 (.I0(x759), .I1(x760), .I2(x761), .I3(n3604), .I4(n3605), .O(n3619));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3620 (.I0(x765), .I1(x766), .I2(x767), .I3(n3618), .I4(n3619), .O(n3620));
  LUT3 #(.INIT(8'hE8)) lut_n3621 (.I0(x774), .I1(x775), .I2(x776), .O(n3621));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3622 (.I0(x765), .I1(x766), .I2(x767), .I3(n3618), .I4(n3619), .O(n3622));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3623 (.I0(x771), .I1(x772), .I2(x773), .I3(n3621), .I4(n3622), .O(n3623));
  LUT3 #(.INIT(8'h96)) lut_n3624 (.I0(n3603), .I1(n3606), .I2(n3607), .O(n3624));
  LUT3 #(.INIT(8'hE8)) lut_n3625 (.I0(n3620), .I1(n3623), .I2(n3624), .O(n3625));
  LUT3 #(.INIT(8'hE8)) lut_n3626 (.I0(x780), .I1(x781), .I2(x782), .O(n3626));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3627 (.I0(x771), .I1(x772), .I2(x773), .I3(n3621), .I4(n3622), .O(n3627));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3628 (.I0(x777), .I1(x778), .I2(x779), .I3(n3626), .I4(n3627), .O(n3628));
  LUT3 #(.INIT(8'hE8)) lut_n3629 (.I0(x786), .I1(x787), .I2(x788), .O(n3629));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3630 (.I0(x777), .I1(x778), .I2(x779), .I3(n3626), .I4(n3627), .O(n3630));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3631 (.I0(x783), .I1(x784), .I2(x785), .I3(n3629), .I4(n3630), .O(n3631));
  LUT3 #(.INIT(8'h96)) lut_n3632 (.I0(n3620), .I1(n3623), .I2(n3624), .O(n3632));
  LUT3 #(.INIT(8'hE8)) lut_n3633 (.I0(n3628), .I1(n3631), .I2(n3632), .O(n3633));
  LUT3 #(.INIT(8'h96)) lut_n3634 (.I0(n3600), .I1(n3608), .I2(n3609), .O(n3634));
  LUT3 #(.INIT(8'hE8)) lut_n3635 (.I0(n3625), .I1(n3633), .I2(n3634), .O(n3635));
  LUT3 #(.INIT(8'hE8)) lut_n3636 (.I0(x792), .I1(x793), .I2(x794), .O(n3636));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3637 (.I0(x783), .I1(x784), .I2(x785), .I3(n3629), .I4(n3630), .O(n3637));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3638 (.I0(x789), .I1(x790), .I2(x791), .I3(n3636), .I4(n3637), .O(n3638));
  LUT3 #(.INIT(8'hE8)) lut_n3639 (.I0(x798), .I1(x799), .I2(x800), .O(n3639));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3640 (.I0(x789), .I1(x790), .I2(x791), .I3(n3636), .I4(n3637), .O(n3640));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3641 (.I0(x795), .I1(x796), .I2(x797), .I3(n3639), .I4(n3640), .O(n3641));
  LUT3 #(.INIT(8'h96)) lut_n3642 (.I0(n3628), .I1(n3631), .I2(n3632), .O(n3642));
  LUT3 #(.INIT(8'hE8)) lut_n3643 (.I0(n3638), .I1(n3641), .I2(n3642), .O(n3643));
  LUT3 #(.INIT(8'hE8)) lut_n3644 (.I0(x804), .I1(x805), .I2(x806), .O(n3644));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3645 (.I0(x795), .I1(x796), .I2(x797), .I3(n3639), .I4(n3640), .O(n3645));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3646 (.I0(x801), .I1(x802), .I2(x803), .I3(n3644), .I4(n3645), .O(n3646));
  LUT3 #(.INIT(8'hE8)) lut_n3647 (.I0(x810), .I1(x811), .I2(x812), .O(n3647));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3648 (.I0(x801), .I1(x802), .I2(x803), .I3(n3644), .I4(n3645), .O(n3648));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3649 (.I0(x807), .I1(x808), .I2(x809), .I3(n3647), .I4(n3648), .O(n3649));
  LUT3 #(.INIT(8'h96)) lut_n3650 (.I0(n3638), .I1(n3641), .I2(n3642), .O(n3650));
  LUT3 #(.INIT(8'hE8)) lut_n3651 (.I0(n3646), .I1(n3649), .I2(n3650), .O(n3651));
  LUT3 #(.INIT(8'h96)) lut_n3652 (.I0(n3625), .I1(n3633), .I2(n3634), .O(n3652));
  LUT3 #(.INIT(8'hE8)) lut_n3653 (.I0(n3643), .I1(n3651), .I2(n3652), .O(n3653));
  LUT3 #(.INIT(8'h96)) lut_n3654 (.I0(n3592), .I1(n3610), .I2(n3611), .O(n3654));
  LUT3 #(.INIT(8'hE8)) lut_n3655 (.I0(n3635), .I1(n3653), .I2(n3654), .O(n3655));
  LUT3 #(.INIT(8'hE8)) lut_n3656 (.I0(x816), .I1(x817), .I2(x818), .O(n3656));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3657 (.I0(x807), .I1(x808), .I2(x809), .I3(n3647), .I4(n3648), .O(n3657));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3658 (.I0(x813), .I1(x814), .I2(x815), .I3(n3656), .I4(n3657), .O(n3658));
  LUT3 #(.INIT(8'hE8)) lut_n3659 (.I0(x822), .I1(x823), .I2(x824), .O(n3659));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3660 (.I0(x813), .I1(x814), .I2(x815), .I3(n3656), .I4(n3657), .O(n3660));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3661 (.I0(x819), .I1(x820), .I2(x821), .I3(n3659), .I4(n3660), .O(n3661));
  LUT3 #(.INIT(8'h96)) lut_n3662 (.I0(n3646), .I1(n3649), .I2(n3650), .O(n3662));
  LUT3 #(.INIT(8'hE8)) lut_n3663 (.I0(n3658), .I1(n3661), .I2(n3662), .O(n3663));
  LUT3 #(.INIT(8'hE8)) lut_n3664 (.I0(x828), .I1(x829), .I2(x830), .O(n3664));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3665 (.I0(x819), .I1(x820), .I2(x821), .I3(n3659), .I4(n3660), .O(n3665));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3666 (.I0(x825), .I1(x826), .I2(x827), .I3(n3664), .I4(n3665), .O(n3666));
  LUT3 #(.INIT(8'hE8)) lut_n3667 (.I0(x834), .I1(x835), .I2(x836), .O(n3667));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3668 (.I0(x825), .I1(x826), .I2(x827), .I3(n3664), .I4(n3665), .O(n3668));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3669 (.I0(x831), .I1(x832), .I2(x833), .I3(n3667), .I4(n3668), .O(n3669));
  LUT3 #(.INIT(8'h96)) lut_n3670 (.I0(n3658), .I1(n3661), .I2(n3662), .O(n3670));
  LUT3 #(.INIT(8'hE8)) lut_n3671 (.I0(n3666), .I1(n3669), .I2(n3670), .O(n3671));
  LUT3 #(.INIT(8'h96)) lut_n3672 (.I0(n3643), .I1(n3651), .I2(n3652), .O(n3672));
  LUT3 #(.INIT(8'hE8)) lut_n3673 (.I0(n3663), .I1(n3671), .I2(n3672), .O(n3673));
  LUT3 #(.INIT(8'hE8)) lut_n3674 (.I0(x840), .I1(x841), .I2(x842), .O(n3674));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3675 (.I0(x831), .I1(x832), .I2(x833), .I3(n3667), .I4(n3668), .O(n3675));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3676 (.I0(x837), .I1(x838), .I2(x839), .I3(n3674), .I4(n3675), .O(n3676));
  LUT3 #(.INIT(8'hE8)) lut_n3677 (.I0(x846), .I1(x847), .I2(x848), .O(n3677));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3678 (.I0(x837), .I1(x838), .I2(x839), .I3(n3674), .I4(n3675), .O(n3678));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3679 (.I0(x843), .I1(x844), .I2(x845), .I3(n3677), .I4(n3678), .O(n3679));
  LUT3 #(.INIT(8'h96)) lut_n3680 (.I0(n3666), .I1(n3669), .I2(n3670), .O(n3680));
  LUT3 #(.INIT(8'hE8)) lut_n3681 (.I0(n3676), .I1(n3679), .I2(n3680), .O(n3681));
  LUT3 #(.INIT(8'hE8)) lut_n3682 (.I0(x852), .I1(x853), .I2(x854), .O(n3682));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3683 (.I0(x843), .I1(x844), .I2(x845), .I3(n3677), .I4(n3678), .O(n3683));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3684 (.I0(x849), .I1(x850), .I2(x851), .I3(n3682), .I4(n3683), .O(n3684));
  LUT3 #(.INIT(8'hE8)) lut_n3685 (.I0(x858), .I1(x859), .I2(x860), .O(n3685));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3686 (.I0(x849), .I1(x850), .I2(x851), .I3(n3682), .I4(n3683), .O(n3686));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3687 (.I0(x855), .I1(x856), .I2(x857), .I3(n3685), .I4(n3686), .O(n3687));
  LUT3 #(.INIT(8'h96)) lut_n3688 (.I0(n3676), .I1(n3679), .I2(n3680), .O(n3688));
  LUT3 #(.INIT(8'hE8)) lut_n3689 (.I0(n3684), .I1(n3687), .I2(n3688), .O(n3689));
  LUT3 #(.INIT(8'h96)) lut_n3690 (.I0(n3663), .I1(n3671), .I2(n3672), .O(n3690));
  LUT3 #(.INIT(8'hE8)) lut_n3691 (.I0(n3681), .I1(n3689), .I2(n3690), .O(n3691));
  LUT3 #(.INIT(8'h96)) lut_n3692 (.I0(n3635), .I1(n3653), .I2(n3654), .O(n3692));
  LUT3 #(.INIT(8'hE8)) lut_n3693 (.I0(n3673), .I1(n3691), .I2(n3692), .O(n3693));
  LUT3 #(.INIT(8'h96)) lut_n3694 (.I0(n3574), .I1(n3612), .I2(n3613), .O(n3694));
  LUT3 #(.INIT(8'hE8)) lut_n3695 (.I0(n3655), .I1(n3693), .I2(n3694), .O(n3695));
  LUT3 #(.INIT(8'hE8)) lut_n3696 (.I0(x864), .I1(x865), .I2(x866), .O(n3696));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3697 (.I0(x855), .I1(x856), .I2(x857), .I3(n3685), .I4(n3686), .O(n3697));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3698 (.I0(x861), .I1(x862), .I2(x863), .I3(n3696), .I4(n3697), .O(n3698));
  LUT3 #(.INIT(8'hE8)) lut_n3699 (.I0(x870), .I1(x871), .I2(x872), .O(n3699));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3700 (.I0(x861), .I1(x862), .I2(x863), .I3(n3696), .I4(n3697), .O(n3700));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3701 (.I0(x867), .I1(x868), .I2(x869), .I3(n3699), .I4(n3700), .O(n3701));
  LUT3 #(.INIT(8'h96)) lut_n3702 (.I0(n3684), .I1(n3687), .I2(n3688), .O(n3702));
  LUT3 #(.INIT(8'hE8)) lut_n3703 (.I0(n3698), .I1(n3701), .I2(n3702), .O(n3703));
  LUT3 #(.INIT(8'hE8)) lut_n3704 (.I0(x876), .I1(x877), .I2(x878), .O(n3704));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3705 (.I0(x867), .I1(x868), .I2(x869), .I3(n3699), .I4(n3700), .O(n3705));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3706 (.I0(x873), .I1(x874), .I2(x875), .I3(n3704), .I4(n3705), .O(n3706));
  LUT3 #(.INIT(8'hE8)) lut_n3707 (.I0(x882), .I1(x883), .I2(x884), .O(n3707));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3708 (.I0(x873), .I1(x874), .I2(x875), .I3(n3704), .I4(n3705), .O(n3708));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3709 (.I0(x879), .I1(x880), .I2(x881), .I3(n3707), .I4(n3708), .O(n3709));
  LUT3 #(.INIT(8'h96)) lut_n3710 (.I0(n3698), .I1(n3701), .I2(n3702), .O(n3710));
  LUT3 #(.INIT(8'hE8)) lut_n3711 (.I0(n3706), .I1(n3709), .I2(n3710), .O(n3711));
  LUT3 #(.INIT(8'h96)) lut_n3712 (.I0(n3681), .I1(n3689), .I2(n3690), .O(n3712));
  LUT3 #(.INIT(8'hE8)) lut_n3713 (.I0(n3703), .I1(n3711), .I2(n3712), .O(n3713));
  LUT3 #(.INIT(8'hE8)) lut_n3714 (.I0(x888), .I1(x889), .I2(x890), .O(n3714));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3715 (.I0(x879), .I1(x880), .I2(x881), .I3(n3707), .I4(n3708), .O(n3715));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3716 (.I0(x885), .I1(x886), .I2(x887), .I3(n3714), .I4(n3715), .O(n3716));
  LUT3 #(.INIT(8'hE8)) lut_n3717 (.I0(x894), .I1(x895), .I2(x896), .O(n3717));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3718 (.I0(x885), .I1(x886), .I2(x887), .I3(n3714), .I4(n3715), .O(n3718));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3719 (.I0(x891), .I1(x892), .I2(x893), .I3(n3717), .I4(n3718), .O(n3719));
  LUT3 #(.INIT(8'h96)) lut_n3720 (.I0(n3706), .I1(n3709), .I2(n3710), .O(n3720));
  LUT3 #(.INIT(8'hE8)) lut_n3721 (.I0(n3716), .I1(n3719), .I2(n3720), .O(n3721));
  LUT3 #(.INIT(8'hE8)) lut_n3722 (.I0(x900), .I1(x901), .I2(x902), .O(n3722));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3723 (.I0(x891), .I1(x892), .I2(x893), .I3(n3717), .I4(n3718), .O(n3723));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3724 (.I0(x897), .I1(x898), .I2(x899), .I3(n3722), .I4(n3723), .O(n3724));
  LUT3 #(.INIT(8'hE8)) lut_n3725 (.I0(x906), .I1(x907), .I2(x908), .O(n3725));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3726 (.I0(x897), .I1(x898), .I2(x899), .I3(n3722), .I4(n3723), .O(n3726));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3727 (.I0(x903), .I1(x904), .I2(x905), .I3(n3725), .I4(n3726), .O(n3727));
  LUT3 #(.INIT(8'h96)) lut_n3728 (.I0(n3716), .I1(n3719), .I2(n3720), .O(n3728));
  LUT3 #(.INIT(8'hE8)) lut_n3729 (.I0(n3724), .I1(n3727), .I2(n3728), .O(n3729));
  LUT3 #(.INIT(8'h96)) lut_n3730 (.I0(n3703), .I1(n3711), .I2(n3712), .O(n3730));
  LUT3 #(.INIT(8'hE8)) lut_n3731 (.I0(n3721), .I1(n3729), .I2(n3730), .O(n3731));
  LUT3 #(.INIT(8'h96)) lut_n3732 (.I0(n3673), .I1(n3691), .I2(n3692), .O(n3732));
  LUT3 #(.INIT(8'hE8)) lut_n3733 (.I0(n3713), .I1(n3731), .I2(n3732), .O(n3733));
  LUT3 #(.INIT(8'hE8)) lut_n3734 (.I0(x912), .I1(x913), .I2(x914), .O(n3734));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3735 (.I0(x903), .I1(x904), .I2(x905), .I3(n3725), .I4(n3726), .O(n3735));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3736 (.I0(x909), .I1(x910), .I2(x911), .I3(n3734), .I4(n3735), .O(n3736));
  LUT3 #(.INIT(8'hE8)) lut_n3737 (.I0(x918), .I1(x919), .I2(x920), .O(n3737));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3738 (.I0(x909), .I1(x910), .I2(x911), .I3(n3734), .I4(n3735), .O(n3738));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3739 (.I0(x915), .I1(x916), .I2(x917), .I3(n3737), .I4(n3738), .O(n3739));
  LUT3 #(.INIT(8'h96)) lut_n3740 (.I0(n3724), .I1(n3727), .I2(n3728), .O(n3740));
  LUT3 #(.INIT(8'hE8)) lut_n3741 (.I0(n3736), .I1(n3739), .I2(n3740), .O(n3741));
  LUT3 #(.INIT(8'hE8)) lut_n3742 (.I0(x924), .I1(x925), .I2(x926), .O(n3742));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3743 (.I0(x915), .I1(x916), .I2(x917), .I3(n3737), .I4(n3738), .O(n3743));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3744 (.I0(x921), .I1(x922), .I2(x923), .I3(n3742), .I4(n3743), .O(n3744));
  LUT3 #(.INIT(8'hE8)) lut_n3745 (.I0(x930), .I1(x931), .I2(x932), .O(n3745));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3746 (.I0(x921), .I1(x922), .I2(x923), .I3(n3742), .I4(n3743), .O(n3746));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3747 (.I0(x927), .I1(x928), .I2(x929), .I3(n3745), .I4(n3746), .O(n3747));
  LUT3 #(.INIT(8'h96)) lut_n3748 (.I0(n3736), .I1(n3739), .I2(n3740), .O(n3748));
  LUT3 #(.INIT(8'hE8)) lut_n3749 (.I0(n3744), .I1(n3747), .I2(n3748), .O(n3749));
  LUT3 #(.INIT(8'h96)) lut_n3750 (.I0(n3721), .I1(n3729), .I2(n3730), .O(n3750));
  LUT3 #(.INIT(8'hE8)) lut_n3751 (.I0(n3741), .I1(n3749), .I2(n3750), .O(n3751));
  LUT3 #(.INIT(8'hE8)) lut_n3752 (.I0(x936), .I1(x937), .I2(x938), .O(n3752));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3753 (.I0(x927), .I1(x928), .I2(x929), .I3(n3745), .I4(n3746), .O(n3753));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3754 (.I0(x933), .I1(x934), .I2(x935), .I3(n3752), .I4(n3753), .O(n3754));
  LUT3 #(.INIT(8'hE8)) lut_n3755 (.I0(x942), .I1(x943), .I2(x944), .O(n3755));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3756 (.I0(x933), .I1(x934), .I2(x935), .I3(n3752), .I4(n3753), .O(n3756));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3757 (.I0(x939), .I1(x940), .I2(x941), .I3(n3755), .I4(n3756), .O(n3757));
  LUT3 #(.INIT(8'h96)) lut_n3758 (.I0(n3744), .I1(n3747), .I2(n3748), .O(n3758));
  LUT3 #(.INIT(8'hE8)) lut_n3759 (.I0(n3754), .I1(n3757), .I2(n3758), .O(n3759));
  LUT3 #(.INIT(8'hE8)) lut_n3760 (.I0(x948), .I1(x949), .I2(x950), .O(n3760));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3761 (.I0(x939), .I1(x940), .I2(x941), .I3(n3755), .I4(n3756), .O(n3761));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3762 (.I0(x945), .I1(x946), .I2(x947), .I3(n3760), .I4(n3761), .O(n3762));
  LUT3 #(.INIT(8'hE8)) lut_n3763 (.I0(x954), .I1(x955), .I2(x956), .O(n3763));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3764 (.I0(x945), .I1(x946), .I2(x947), .I3(n3760), .I4(n3761), .O(n3764));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3765 (.I0(x951), .I1(x952), .I2(x953), .I3(n3763), .I4(n3764), .O(n3765));
  LUT3 #(.INIT(8'h96)) lut_n3766 (.I0(n3754), .I1(n3757), .I2(n3758), .O(n3766));
  LUT3 #(.INIT(8'hE8)) lut_n3767 (.I0(n3762), .I1(n3765), .I2(n3766), .O(n3767));
  LUT3 #(.INIT(8'h96)) lut_n3768 (.I0(n3741), .I1(n3749), .I2(n3750), .O(n3768));
  LUT3 #(.INIT(8'hE8)) lut_n3769 (.I0(n3759), .I1(n3767), .I2(n3768), .O(n3769));
  LUT3 #(.INIT(8'h96)) lut_n3770 (.I0(n3713), .I1(n3731), .I2(n3732), .O(n3770));
  LUT3 #(.INIT(8'hE8)) lut_n3771 (.I0(n3751), .I1(n3769), .I2(n3770), .O(n3771));
  LUT3 #(.INIT(8'h96)) lut_n3772 (.I0(n3655), .I1(n3693), .I2(n3694), .O(n3772));
  LUT3 #(.INIT(8'hE8)) lut_n3773 (.I0(n3733), .I1(n3771), .I2(n3772), .O(n3773));
  LUT3 #(.INIT(8'h96)) lut_n3774 (.I0(n3536), .I1(n3614), .I2(n3615), .O(n3774));
  LUT3 #(.INIT(8'hE8)) lut_n3775 (.I0(n3695), .I1(n3773), .I2(n3774), .O(n3775));
  LUT3 #(.INIT(8'hE8)) lut_n3776 (.I0(x960), .I1(x961), .I2(x962), .O(n3776));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3777 (.I0(x951), .I1(x952), .I2(x953), .I3(n3763), .I4(n3764), .O(n3777));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3778 (.I0(x957), .I1(x958), .I2(x959), .I3(n3776), .I4(n3777), .O(n3778));
  LUT3 #(.INIT(8'hE8)) lut_n3779 (.I0(x966), .I1(x967), .I2(x968), .O(n3779));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3780 (.I0(x957), .I1(x958), .I2(x959), .I3(n3776), .I4(n3777), .O(n3780));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3781 (.I0(x963), .I1(x964), .I2(x965), .I3(n3779), .I4(n3780), .O(n3781));
  LUT3 #(.INIT(8'h96)) lut_n3782 (.I0(n3762), .I1(n3765), .I2(n3766), .O(n3782));
  LUT3 #(.INIT(8'hE8)) lut_n3783 (.I0(n3778), .I1(n3781), .I2(n3782), .O(n3783));
  LUT3 #(.INIT(8'hE8)) lut_n3784 (.I0(x972), .I1(x973), .I2(x974), .O(n3784));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3785 (.I0(x963), .I1(x964), .I2(x965), .I3(n3779), .I4(n3780), .O(n3785));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3786 (.I0(x969), .I1(x970), .I2(x971), .I3(n3784), .I4(n3785), .O(n3786));
  LUT3 #(.INIT(8'hE8)) lut_n3787 (.I0(x978), .I1(x979), .I2(x980), .O(n3787));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3788 (.I0(x969), .I1(x970), .I2(x971), .I3(n3784), .I4(n3785), .O(n3788));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3789 (.I0(x975), .I1(x976), .I2(x977), .I3(n3787), .I4(n3788), .O(n3789));
  LUT3 #(.INIT(8'h96)) lut_n3790 (.I0(n3778), .I1(n3781), .I2(n3782), .O(n3790));
  LUT3 #(.INIT(8'hE8)) lut_n3791 (.I0(n3786), .I1(n3789), .I2(n3790), .O(n3791));
  LUT3 #(.INIT(8'h96)) lut_n3792 (.I0(n3759), .I1(n3767), .I2(n3768), .O(n3792));
  LUT3 #(.INIT(8'hE8)) lut_n3793 (.I0(n3783), .I1(n3791), .I2(n3792), .O(n3793));
  LUT3 #(.INIT(8'hE8)) lut_n3794 (.I0(x984), .I1(x985), .I2(x986), .O(n3794));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3795 (.I0(x975), .I1(x976), .I2(x977), .I3(n3787), .I4(n3788), .O(n3795));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3796 (.I0(x981), .I1(x982), .I2(x983), .I3(n3794), .I4(n3795), .O(n3796));
  LUT3 #(.INIT(8'hE8)) lut_n3797 (.I0(x990), .I1(x991), .I2(x992), .O(n3797));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3798 (.I0(x981), .I1(x982), .I2(x983), .I3(n3794), .I4(n3795), .O(n3798));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3799 (.I0(x987), .I1(x988), .I2(x989), .I3(n3797), .I4(n3798), .O(n3799));
  LUT3 #(.INIT(8'h96)) lut_n3800 (.I0(n3786), .I1(n3789), .I2(n3790), .O(n3800));
  LUT3 #(.INIT(8'hE8)) lut_n3801 (.I0(n3796), .I1(n3799), .I2(n3800), .O(n3801));
  LUT3 #(.INIT(8'hE8)) lut_n3802 (.I0(x996), .I1(x997), .I2(x998), .O(n3802));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3803 (.I0(x987), .I1(x988), .I2(x989), .I3(n3797), .I4(n3798), .O(n3803));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3804 (.I0(x993), .I1(x994), .I2(x995), .I3(n3802), .I4(n3803), .O(n3804));
  LUT3 #(.INIT(8'hE8)) lut_n3805 (.I0(x1002), .I1(x1003), .I2(x1004), .O(n3805));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3806 (.I0(x993), .I1(x994), .I2(x995), .I3(n3802), .I4(n3803), .O(n3806));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3807 (.I0(x999), .I1(x1000), .I2(x1001), .I3(n3805), .I4(n3806), .O(n3807));
  LUT3 #(.INIT(8'h96)) lut_n3808 (.I0(n3796), .I1(n3799), .I2(n3800), .O(n3808));
  LUT3 #(.INIT(8'hE8)) lut_n3809 (.I0(n3804), .I1(n3807), .I2(n3808), .O(n3809));
  LUT3 #(.INIT(8'h96)) lut_n3810 (.I0(n3783), .I1(n3791), .I2(n3792), .O(n3810));
  LUT3 #(.INIT(8'hE8)) lut_n3811 (.I0(n3801), .I1(n3809), .I2(n3810), .O(n3811));
  LUT3 #(.INIT(8'h96)) lut_n3812 (.I0(n3751), .I1(n3769), .I2(n3770), .O(n3812));
  LUT3 #(.INIT(8'hE8)) lut_n3813 (.I0(n3793), .I1(n3811), .I2(n3812), .O(n3813));
  LUT3 #(.INIT(8'hE8)) lut_n3814 (.I0(x1008), .I1(x1009), .I2(x1010), .O(n3814));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3815 (.I0(x999), .I1(x1000), .I2(x1001), .I3(n3805), .I4(n3806), .O(n3815));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3816 (.I0(x1005), .I1(x1006), .I2(x1007), .I3(n3814), .I4(n3815), .O(n3816));
  LUT3 #(.INIT(8'hE8)) lut_n3817 (.I0(x1014), .I1(x1015), .I2(x1016), .O(n3817));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3818 (.I0(x1005), .I1(x1006), .I2(x1007), .I3(n3814), .I4(n3815), .O(n3818));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3819 (.I0(x1011), .I1(x1012), .I2(x1013), .I3(n3817), .I4(n3818), .O(n3819));
  LUT3 #(.INIT(8'h96)) lut_n3820 (.I0(n3804), .I1(n3807), .I2(n3808), .O(n3820));
  LUT3 #(.INIT(8'hE8)) lut_n3821 (.I0(n3816), .I1(n3819), .I2(n3820), .O(n3821));
  LUT3 #(.INIT(8'hE8)) lut_n3822 (.I0(x1020), .I1(x1021), .I2(x1022), .O(n3822));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3823 (.I0(x1011), .I1(x1012), .I2(x1013), .I3(n3817), .I4(n3818), .O(n3823));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3824 (.I0(x1017), .I1(x1018), .I2(x1019), .I3(n3822), .I4(n3823), .O(n3824));
  LUT3 #(.INIT(8'hE8)) lut_n3825 (.I0(x1026), .I1(x1027), .I2(x1028), .O(n3825));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3826 (.I0(x1017), .I1(x1018), .I2(x1019), .I3(n3822), .I4(n3823), .O(n3826));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3827 (.I0(x1023), .I1(x1024), .I2(x1025), .I3(n3825), .I4(n3826), .O(n3827));
  LUT3 #(.INIT(8'h96)) lut_n3828 (.I0(n3816), .I1(n3819), .I2(n3820), .O(n3828));
  LUT3 #(.INIT(8'hE8)) lut_n3829 (.I0(n3824), .I1(n3827), .I2(n3828), .O(n3829));
  LUT3 #(.INIT(8'h96)) lut_n3830 (.I0(n3801), .I1(n3809), .I2(n3810), .O(n3830));
  LUT3 #(.INIT(8'hE8)) lut_n3831 (.I0(n3821), .I1(n3829), .I2(n3830), .O(n3831));
  LUT3 #(.INIT(8'hE8)) lut_n3832 (.I0(x1032), .I1(x1033), .I2(x1034), .O(n3832));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3833 (.I0(x1023), .I1(x1024), .I2(x1025), .I3(n3825), .I4(n3826), .O(n3833));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3834 (.I0(x1029), .I1(x1030), .I2(x1031), .I3(n3832), .I4(n3833), .O(n3834));
  LUT3 #(.INIT(8'hE8)) lut_n3835 (.I0(x1038), .I1(x1039), .I2(x1040), .O(n3835));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3836 (.I0(x1029), .I1(x1030), .I2(x1031), .I3(n3832), .I4(n3833), .O(n3836));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3837 (.I0(x1035), .I1(x1036), .I2(x1037), .I3(n3835), .I4(n3836), .O(n3837));
  LUT3 #(.INIT(8'h96)) lut_n3838 (.I0(n3824), .I1(n3827), .I2(n3828), .O(n3838));
  LUT3 #(.INIT(8'hE8)) lut_n3839 (.I0(n3834), .I1(n3837), .I2(n3838), .O(n3839));
  LUT3 #(.INIT(8'hE8)) lut_n3840 (.I0(x1044), .I1(x1045), .I2(x1046), .O(n3840));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3841 (.I0(x1035), .I1(x1036), .I2(x1037), .I3(n3835), .I4(n3836), .O(n3841));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3842 (.I0(x1041), .I1(x1042), .I2(x1043), .I3(n3840), .I4(n3841), .O(n3842));
  LUT3 #(.INIT(8'hE8)) lut_n3843 (.I0(x1050), .I1(x1051), .I2(x1052), .O(n3843));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3844 (.I0(x1041), .I1(x1042), .I2(x1043), .I3(n3840), .I4(n3841), .O(n3844));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3845 (.I0(x1047), .I1(x1048), .I2(x1049), .I3(n3843), .I4(n3844), .O(n3845));
  LUT3 #(.INIT(8'h96)) lut_n3846 (.I0(n3834), .I1(n3837), .I2(n3838), .O(n3846));
  LUT3 #(.INIT(8'hE8)) lut_n3847 (.I0(n3842), .I1(n3845), .I2(n3846), .O(n3847));
  LUT3 #(.INIT(8'h96)) lut_n3848 (.I0(n3821), .I1(n3829), .I2(n3830), .O(n3848));
  LUT3 #(.INIT(8'hE8)) lut_n3849 (.I0(n3839), .I1(n3847), .I2(n3848), .O(n3849));
  LUT3 #(.INIT(8'h96)) lut_n3850 (.I0(n3793), .I1(n3811), .I2(n3812), .O(n3850));
  LUT3 #(.INIT(8'hE8)) lut_n3851 (.I0(n3831), .I1(n3849), .I2(n3850), .O(n3851));
  LUT3 #(.INIT(8'h96)) lut_n3852 (.I0(n3733), .I1(n3771), .I2(n3772), .O(n3852));
  LUT3 #(.INIT(8'hE8)) lut_n3853 (.I0(n3813), .I1(n3851), .I2(n3852), .O(n3853));
  LUT3 #(.INIT(8'hE8)) lut_n3854 (.I0(x1056), .I1(x1057), .I2(x1058), .O(n3854));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3855 (.I0(x1047), .I1(x1048), .I2(x1049), .I3(n3843), .I4(n3844), .O(n3855));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3856 (.I0(x1053), .I1(x1054), .I2(x1055), .I3(n3854), .I4(n3855), .O(n3856));
  LUT3 #(.INIT(8'hE8)) lut_n3857 (.I0(x1062), .I1(x1063), .I2(x1064), .O(n3857));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3858 (.I0(x1053), .I1(x1054), .I2(x1055), .I3(n3854), .I4(n3855), .O(n3858));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3859 (.I0(x1059), .I1(x1060), .I2(x1061), .I3(n3857), .I4(n3858), .O(n3859));
  LUT3 #(.INIT(8'h96)) lut_n3860 (.I0(n3842), .I1(n3845), .I2(n3846), .O(n3860));
  LUT3 #(.INIT(8'hE8)) lut_n3861 (.I0(n3856), .I1(n3859), .I2(n3860), .O(n3861));
  LUT3 #(.INIT(8'hE8)) lut_n3862 (.I0(x1068), .I1(x1069), .I2(x1070), .O(n3862));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3863 (.I0(x1059), .I1(x1060), .I2(x1061), .I3(n3857), .I4(n3858), .O(n3863));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3864 (.I0(x1065), .I1(x1066), .I2(x1067), .I3(n3862), .I4(n3863), .O(n3864));
  LUT3 #(.INIT(8'hE8)) lut_n3865 (.I0(x1074), .I1(x1075), .I2(x1076), .O(n3865));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3866 (.I0(x1065), .I1(x1066), .I2(x1067), .I3(n3862), .I4(n3863), .O(n3866));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3867 (.I0(x1071), .I1(x1072), .I2(x1073), .I3(n3865), .I4(n3866), .O(n3867));
  LUT3 #(.INIT(8'h96)) lut_n3868 (.I0(n3856), .I1(n3859), .I2(n3860), .O(n3868));
  LUT3 #(.INIT(8'hE8)) lut_n3869 (.I0(n3864), .I1(n3867), .I2(n3868), .O(n3869));
  LUT3 #(.INIT(8'h96)) lut_n3870 (.I0(n3839), .I1(n3847), .I2(n3848), .O(n3870));
  LUT3 #(.INIT(8'hE8)) lut_n3871 (.I0(n3861), .I1(n3869), .I2(n3870), .O(n3871));
  LUT3 #(.INIT(8'hE8)) lut_n3872 (.I0(x1080), .I1(x1081), .I2(x1082), .O(n3872));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3873 (.I0(x1071), .I1(x1072), .I2(x1073), .I3(n3865), .I4(n3866), .O(n3873));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3874 (.I0(x1077), .I1(x1078), .I2(x1079), .I3(n3872), .I4(n3873), .O(n3874));
  LUT3 #(.INIT(8'hE8)) lut_n3875 (.I0(x1086), .I1(x1087), .I2(x1088), .O(n3875));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3876 (.I0(x1077), .I1(x1078), .I2(x1079), .I3(n3872), .I4(n3873), .O(n3876));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3877 (.I0(x1083), .I1(x1084), .I2(x1085), .I3(n3875), .I4(n3876), .O(n3877));
  LUT3 #(.INIT(8'h96)) lut_n3878 (.I0(n3864), .I1(n3867), .I2(n3868), .O(n3878));
  LUT3 #(.INIT(8'hE8)) lut_n3879 (.I0(n3874), .I1(n3877), .I2(n3878), .O(n3879));
  LUT3 #(.INIT(8'hE8)) lut_n3880 (.I0(x1092), .I1(x1093), .I2(x1094), .O(n3880));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3881 (.I0(x1083), .I1(x1084), .I2(x1085), .I3(n3875), .I4(n3876), .O(n3881));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3882 (.I0(x1089), .I1(x1090), .I2(x1091), .I3(n3880), .I4(n3881), .O(n3882));
  LUT3 #(.INIT(8'hE8)) lut_n3883 (.I0(x1098), .I1(x1099), .I2(x1100), .O(n3883));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3884 (.I0(x1089), .I1(x1090), .I2(x1091), .I3(n3880), .I4(n3881), .O(n3884));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3885 (.I0(x1095), .I1(x1096), .I2(x1097), .I3(n3883), .I4(n3884), .O(n3885));
  LUT3 #(.INIT(8'h96)) lut_n3886 (.I0(n3874), .I1(n3877), .I2(n3878), .O(n3886));
  LUT3 #(.INIT(8'hE8)) lut_n3887 (.I0(n3882), .I1(n3885), .I2(n3886), .O(n3887));
  LUT3 #(.INIT(8'h96)) lut_n3888 (.I0(n3861), .I1(n3869), .I2(n3870), .O(n3888));
  LUT3 #(.INIT(8'hE8)) lut_n3889 (.I0(n3879), .I1(n3887), .I2(n3888), .O(n3889));
  LUT3 #(.INIT(8'h96)) lut_n3890 (.I0(n3831), .I1(n3849), .I2(n3850), .O(n3890));
  LUT3 #(.INIT(8'hE8)) lut_n3891 (.I0(n3871), .I1(n3889), .I2(n3890), .O(n3891));
  LUT3 #(.INIT(8'hE8)) lut_n3892 (.I0(x1104), .I1(x1105), .I2(x1106), .O(n3892));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3893 (.I0(x1095), .I1(x1096), .I2(x1097), .I3(n3883), .I4(n3884), .O(n3893));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3894 (.I0(x1101), .I1(x1102), .I2(x1103), .I3(n3892), .I4(n3893), .O(n3894));
  LUT3 #(.INIT(8'hE8)) lut_n3895 (.I0(x1110), .I1(x1111), .I2(x1112), .O(n3895));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3896 (.I0(x1101), .I1(x1102), .I2(x1103), .I3(n3892), .I4(n3893), .O(n3896));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3897 (.I0(x1107), .I1(x1108), .I2(x1109), .I3(n3895), .I4(n3896), .O(n3897));
  LUT3 #(.INIT(8'h96)) lut_n3898 (.I0(n3882), .I1(n3885), .I2(n3886), .O(n3898));
  LUT3 #(.INIT(8'hE8)) lut_n3899 (.I0(n3894), .I1(n3897), .I2(n3898), .O(n3899));
  LUT3 #(.INIT(8'hE8)) lut_n3900 (.I0(x1116), .I1(x1117), .I2(x1118), .O(n3900));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3901 (.I0(x1107), .I1(x1108), .I2(x1109), .I3(n3895), .I4(n3896), .O(n3901));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3902 (.I0(x1113), .I1(x1114), .I2(x1115), .I3(n3900), .I4(n3901), .O(n3902));
  LUT3 #(.INIT(8'hE8)) lut_n3903 (.I0(x1122), .I1(x1123), .I2(x1124), .O(n3903));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3904 (.I0(x1113), .I1(x1114), .I2(x1115), .I3(n3900), .I4(n3901), .O(n3904));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3905 (.I0(x1119), .I1(x1120), .I2(x1121), .I3(n3903), .I4(n3904), .O(n3905));
  LUT3 #(.INIT(8'h96)) lut_n3906 (.I0(n3894), .I1(n3897), .I2(n3898), .O(n3906));
  LUT3 #(.INIT(8'hE8)) lut_n3907 (.I0(n3902), .I1(n3905), .I2(n3906), .O(n3907));
  LUT3 #(.INIT(8'h96)) lut_n3908 (.I0(n3879), .I1(n3887), .I2(n3888), .O(n3908));
  LUT3 #(.INIT(8'hE8)) lut_n3909 (.I0(n3899), .I1(n3907), .I2(n3908), .O(n3909));
  LUT3 #(.INIT(8'hE8)) lut_n3910 (.I0(x1128), .I1(x1129), .I2(x1130), .O(n3910));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3911 (.I0(x1119), .I1(x1120), .I2(x1121), .I3(n3903), .I4(n3904), .O(n3911));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3912 (.I0(x1125), .I1(x1126), .I2(x1127), .I3(n3910), .I4(n3911), .O(n3912));
  LUT3 #(.INIT(8'hE8)) lut_n3913 (.I0(x1134), .I1(x1135), .I2(x1136), .O(n3913));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3914 (.I0(x1125), .I1(x1126), .I2(x1127), .I3(n3910), .I4(n3911), .O(n3914));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3915 (.I0(x1131), .I1(x1132), .I2(x1133), .I3(n3913), .I4(n3914), .O(n3915));
  LUT3 #(.INIT(8'h96)) lut_n3916 (.I0(n3902), .I1(n3905), .I2(n3906), .O(n3916));
  LUT3 #(.INIT(8'hE8)) lut_n3917 (.I0(n3912), .I1(n3915), .I2(n3916), .O(n3917));
  LUT3 #(.INIT(8'hE8)) lut_n3918 (.I0(x1140), .I1(x1141), .I2(x1142), .O(n3918));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3919 (.I0(x1131), .I1(x1132), .I2(x1133), .I3(n3913), .I4(n3914), .O(n3919));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3920 (.I0(x1137), .I1(x1138), .I2(x1139), .I3(n3918), .I4(n3919), .O(n3920));
  LUT3 #(.INIT(8'hE8)) lut_n3921 (.I0(x1146), .I1(x1147), .I2(x1148), .O(n3921));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3922 (.I0(x1137), .I1(x1138), .I2(x1139), .I3(n3918), .I4(n3919), .O(n3922));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3923 (.I0(x1143), .I1(x1144), .I2(x1145), .I3(n3921), .I4(n3922), .O(n3923));
  LUT3 #(.INIT(8'h96)) lut_n3924 (.I0(n3912), .I1(n3915), .I2(n3916), .O(n3924));
  LUT3 #(.INIT(8'hE8)) lut_n3925 (.I0(n3920), .I1(n3923), .I2(n3924), .O(n3925));
  LUT3 #(.INIT(8'h96)) lut_n3926 (.I0(n3899), .I1(n3907), .I2(n3908), .O(n3926));
  LUT3 #(.INIT(8'hE8)) lut_n3927 (.I0(n3917), .I1(n3925), .I2(n3926), .O(n3927));
  LUT3 #(.INIT(8'h96)) lut_n3928 (.I0(n3871), .I1(n3889), .I2(n3890), .O(n3928));
  LUT3 #(.INIT(8'hE8)) lut_n3929 (.I0(n3909), .I1(n3927), .I2(n3928), .O(n3929));
  LUT3 #(.INIT(8'h96)) lut_n3930 (.I0(n3813), .I1(n3851), .I2(n3852), .O(n3930));
  LUT3 #(.INIT(8'hE8)) lut_n3931 (.I0(n3891), .I1(n3929), .I2(n3930), .O(n3931));
  LUT3 #(.INIT(8'h96)) lut_n3932 (.I0(n3695), .I1(n3773), .I2(n3774), .O(n3932));
  LUT3 #(.INIT(8'hE8)) lut_n3933 (.I0(n3853), .I1(n3931), .I2(n3932), .O(n3933));
  LUT3 #(.INIT(8'h96)) lut_n3934 (.I0(n3300), .I1(n3458), .I2(n3616), .O(n3934));
  LUT3 #(.INIT(8'hE8)) lut_n3935 (.I0(n3775), .I1(n3933), .I2(n3934), .O(n3935));
  LUT3 #(.INIT(8'hE8)) lut_n3936 (.I0(x1152), .I1(x1153), .I2(x1154), .O(n3936));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3937 (.I0(x1143), .I1(x1144), .I2(x1145), .I3(n3921), .I4(n3922), .O(n3937));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3938 (.I0(x1149), .I1(x1150), .I2(x1151), .I3(n3936), .I4(n3937), .O(n3938));
  LUT3 #(.INIT(8'hE8)) lut_n3939 (.I0(x1158), .I1(x1159), .I2(x1160), .O(n3939));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3940 (.I0(x1149), .I1(x1150), .I2(x1151), .I3(n3936), .I4(n3937), .O(n3940));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3941 (.I0(x1155), .I1(x1156), .I2(x1157), .I3(n3939), .I4(n3940), .O(n3941));
  LUT3 #(.INIT(8'h96)) lut_n3942 (.I0(n3920), .I1(n3923), .I2(n3924), .O(n3942));
  LUT3 #(.INIT(8'hE8)) lut_n3943 (.I0(n3938), .I1(n3941), .I2(n3942), .O(n3943));
  LUT3 #(.INIT(8'hE8)) lut_n3944 (.I0(x1164), .I1(x1165), .I2(x1166), .O(n3944));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3945 (.I0(x1155), .I1(x1156), .I2(x1157), .I3(n3939), .I4(n3940), .O(n3945));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3946 (.I0(x1161), .I1(x1162), .I2(x1163), .I3(n3944), .I4(n3945), .O(n3946));
  LUT3 #(.INIT(8'hE8)) lut_n3947 (.I0(x1170), .I1(x1171), .I2(x1172), .O(n3947));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3948 (.I0(x1161), .I1(x1162), .I2(x1163), .I3(n3944), .I4(n3945), .O(n3948));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3949 (.I0(x1167), .I1(x1168), .I2(x1169), .I3(n3947), .I4(n3948), .O(n3949));
  LUT3 #(.INIT(8'h96)) lut_n3950 (.I0(n3938), .I1(n3941), .I2(n3942), .O(n3950));
  LUT3 #(.INIT(8'hE8)) lut_n3951 (.I0(n3946), .I1(n3949), .I2(n3950), .O(n3951));
  LUT3 #(.INIT(8'h96)) lut_n3952 (.I0(n3917), .I1(n3925), .I2(n3926), .O(n3952));
  LUT3 #(.INIT(8'hE8)) lut_n3953 (.I0(n3943), .I1(n3951), .I2(n3952), .O(n3953));
  LUT3 #(.INIT(8'hE8)) lut_n3954 (.I0(x1176), .I1(x1177), .I2(x1178), .O(n3954));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3955 (.I0(x1167), .I1(x1168), .I2(x1169), .I3(n3947), .I4(n3948), .O(n3955));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3956 (.I0(x1173), .I1(x1174), .I2(x1175), .I3(n3954), .I4(n3955), .O(n3956));
  LUT3 #(.INIT(8'hE8)) lut_n3957 (.I0(x1182), .I1(x1183), .I2(x1184), .O(n3957));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3958 (.I0(x1173), .I1(x1174), .I2(x1175), .I3(n3954), .I4(n3955), .O(n3958));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3959 (.I0(x1179), .I1(x1180), .I2(x1181), .I3(n3957), .I4(n3958), .O(n3959));
  LUT3 #(.INIT(8'h96)) lut_n3960 (.I0(n3946), .I1(n3949), .I2(n3950), .O(n3960));
  LUT3 #(.INIT(8'hE8)) lut_n3961 (.I0(n3956), .I1(n3959), .I2(n3960), .O(n3961));
  LUT3 #(.INIT(8'hE8)) lut_n3962 (.I0(x1188), .I1(x1189), .I2(x1190), .O(n3962));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3963 (.I0(x1179), .I1(x1180), .I2(x1181), .I3(n3957), .I4(n3958), .O(n3963));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3964 (.I0(x1185), .I1(x1186), .I2(x1187), .I3(n3962), .I4(n3963), .O(n3964));
  LUT3 #(.INIT(8'hE8)) lut_n3965 (.I0(x1194), .I1(x1195), .I2(x1196), .O(n3965));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3966 (.I0(x1185), .I1(x1186), .I2(x1187), .I3(n3962), .I4(n3963), .O(n3966));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3967 (.I0(x1191), .I1(x1192), .I2(x1193), .I3(n3965), .I4(n3966), .O(n3967));
  LUT3 #(.INIT(8'h96)) lut_n3968 (.I0(n3956), .I1(n3959), .I2(n3960), .O(n3968));
  LUT3 #(.INIT(8'hE8)) lut_n3969 (.I0(n3964), .I1(n3967), .I2(n3968), .O(n3969));
  LUT3 #(.INIT(8'h96)) lut_n3970 (.I0(n3943), .I1(n3951), .I2(n3952), .O(n3970));
  LUT3 #(.INIT(8'hE8)) lut_n3971 (.I0(n3961), .I1(n3969), .I2(n3970), .O(n3971));
  LUT3 #(.INIT(8'h96)) lut_n3972 (.I0(n3909), .I1(n3927), .I2(n3928), .O(n3972));
  LUT3 #(.INIT(8'hE8)) lut_n3973 (.I0(n3953), .I1(n3971), .I2(n3972), .O(n3973));
  LUT3 #(.INIT(8'hE8)) lut_n3974 (.I0(x1200), .I1(x1201), .I2(x1202), .O(n3974));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3975 (.I0(x1191), .I1(x1192), .I2(x1193), .I3(n3965), .I4(n3966), .O(n3975));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3976 (.I0(x1197), .I1(x1198), .I2(x1199), .I3(n3974), .I4(n3975), .O(n3976));
  LUT3 #(.INIT(8'hE8)) lut_n3977 (.I0(x1206), .I1(x1207), .I2(x1208), .O(n3977));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3978 (.I0(x1197), .I1(x1198), .I2(x1199), .I3(n3974), .I4(n3975), .O(n3978));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3979 (.I0(x1203), .I1(x1204), .I2(x1205), .I3(n3977), .I4(n3978), .O(n3979));
  LUT3 #(.INIT(8'h96)) lut_n3980 (.I0(n3964), .I1(n3967), .I2(n3968), .O(n3980));
  LUT3 #(.INIT(8'hE8)) lut_n3981 (.I0(n3976), .I1(n3979), .I2(n3980), .O(n3981));
  LUT3 #(.INIT(8'hE8)) lut_n3982 (.I0(x1212), .I1(x1213), .I2(x1214), .O(n3982));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3983 (.I0(x1203), .I1(x1204), .I2(x1205), .I3(n3977), .I4(n3978), .O(n3983));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3984 (.I0(x1209), .I1(x1210), .I2(x1211), .I3(n3982), .I4(n3983), .O(n3984));
  LUT3 #(.INIT(8'hE8)) lut_n3985 (.I0(x1218), .I1(x1219), .I2(x1220), .O(n3985));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3986 (.I0(x1209), .I1(x1210), .I2(x1211), .I3(n3982), .I4(n3983), .O(n3986));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3987 (.I0(x1215), .I1(x1216), .I2(x1217), .I3(n3985), .I4(n3986), .O(n3987));
  LUT3 #(.INIT(8'h96)) lut_n3988 (.I0(n3976), .I1(n3979), .I2(n3980), .O(n3988));
  LUT3 #(.INIT(8'hE8)) lut_n3989 (.I0(n3984), .I1(n3987), .I2(n3988), .O(n3989));
  LUT3 #(.INIT(8'h96)) lut_n3990 (.I0(n3961), .I1(n3969), .I2(n3970), .O(n3990));
  LUT3 #(.INIT(8'hE8)) lut_n3991 (.I0(n3981), .I1(n3989), .I2(n3990), .O(n3991));
  LUT3 #(.INIT(8'hE8)) lut_n3992 (.I0(x1224), .I1(x1225), .I2(x1226), .O(n3992));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3993 (.I0(x1215), .I1(x1216), .I2(x1217), .I3(n3985), .I4(n3986), .O(n3993));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3994 (.I0(x1221), .I1(x1222), .I2(x1223), .I3(n3992), .I4(n3993), .O(n3994));
  LUT3 #(.INIT(8'hE8)) lut_n3995 (.I0(x1230), .I1(x1231), .I2(x1232), .O(n3995));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3996 (.I0(x1221), .I1(x1222), .I2(x1223), .I3(n3992), .I4(n3993), .O(n3996));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3997 (.I0(x1227), .I1(x1228), .I2(x1229), .I3(n3995), .I4(n3996), .O(n3997));
  LUT3 #(.INIT(8'h96)) lut_n3998 (.I0(n3984), .I1(n3987), .I2(n3988), .O(n3998));
  LUT3 #(.INIT(8'hE8)) lut_n3999 (.I0(n3994), .I1(n3997), .I2(n3998), .O(n3999));
  LUT3 #(.INIT(8'hE8)) lut_n4000 (.I0(x1236), .I1(x1237), .I2(x1238), .O(n4000));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4001 (.I0(x1227), .I1(x1228), .I2(x1229), .I3(n3995), .I4(n3996), .O(n4001));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4002 (.I0(x1233), .I1(x1234), .I2(x1235), .I3(n4000), .I4(n4001), .O(n4002));
  LUT3 #(.INIT(8'hE8)) lut_n4003 (.I0(x1242), .I1(x1243), .I2(x1244), .O(n4003));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4004 (.I0(x1233), .I1(x1234), .I2(x1235), .I3(n4000), .I4(n4001), .O(n4004));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4005 (.I0(x1239), .I1(x1240), .I2(x1241), .I3(n4003), .I4(n4004), .O(n4005));
  LUT3 #(.INIT(8'h96)) lut_n4006 (.I0(n3994), .I1(n3997), .I2(n3998), .O(n4006));
  LUT3 #(.INIT(8'hE8)) lut_n4007 (.I0(n4002), .I1(n4005), .I2(n4006), .O(n4007));
  LUT3 #(.INIT(8'h96)) lut_n4008 (.I0(n3981), .I1(n3989), .I2(n3990), .O(n4008));
  LUT3 #(.INIT(8'hE8)) lut_n4009 (.I0(n3999), .I1(n4007), .I2(n4008), .O(n4009));
  LUT3 #(.INIT(8'h96)) lut_n4010 (.I0(n3953), .I1(n3971), .I2(n3972), .O(n4010));
  LUT3 #(.INIT(8'hE8)) lut_n4011 (.I0(n3991), .I1(n4009), .I2(n4010), .O(n4011));
  LUT3 #(.INIT(8'h96)) lut_n4012 (.I0(n3891), .I1(n3929), .I2(n3930), .O(n4012));
  LUT3 #(.INIT(8'hE8)) lut_n4013 (.I0(n3973), .I1(n4011), .I2(n4012), .O(n4013));
  LUT3 #(.INIT(8'hE8)) lut_n4014 (.I0(x1248), .I1(x1249), .I2(x1250), .O(n4014));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4015 (.I0(x1239), .I1(x1240), .I2(x1241), .I3(n4003), .I4(n4004), .O(n4015));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4016 (.I0(x1245), .I1(x1246), .I2(x1247), .I3(n4014), .I4(n4015), .O(n4016));
  LUT3 #(.INIT(8'hE8)) lut_n4017 (.I0(x1254), .I1(x1255), .I2(x1256), .O(n4017));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4018 (.I0(x1245), .I1(x1246), .I2(x1247), .I3(n4014), .I4(n4015), .O(n4018));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4019 (.I0(x1251), .I1(x1252), .I2(x1253), .I3(n4017), .I4(n4018), .O(n4019));
  LUT3 #(.INIT(8'h96)) lut_n4020 (.I0(n4002), .I1(n4005), .I2(n4006), .O(n4020));
  LUT3 #(.INIT(8'hE8)) lut_n4021 (.I0(n4016), .I1(n4019), .I2(n4020), .O(n4021));
  LUT3 #(.INIT(8'hE8)) lut_n4022 (.I0(x1260), .I1(x1261), .I2(x1262), .O(n4022));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4023 (.I0(x1251), .I1(x1252), .I2(x1253), .I3(n4017), .I4(n4018), .O(n4023));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4024 (.I0(x1257), .I1(x1258), .I2(x1259), .I3(n4022), .I4(n4023), .O(n4024));
  LUT3 #(.INIT(8'hE8)) lut_n4025 (.I0(x1266), .I1(x1267), .I2(x1268), .O(n4025));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4026 (.I0(x1257), .I1(x1258), .I2(x1259), .I3(n4022), .I4(n4023), .O(n4026));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4027 (.I0(x1263), .I1(x1264), .I2(x1265), .I3(n4025), .I4(n4026), .O(n4027));
  LUT3 #(.INIT(8'h96)) lut_n4028 (.I0(n4016), .I1(n4019), .I2(n4020), .O(n4028));
  LUT3 #(.INIT(8'hE8)) lut_n4029 (.I0(n4024), .I1(n4027), .I2(n4028), .O(n4029));
  LUT3 #(.INIT(8'h96)) lut_n4030 (.I0(n3999), .I1(n4007), .I2(n4008), .O(n4030));
  LUT3 #(.INIT(8'hE8)) lut_n4031 (.I0(n4021), .I1(n4029), .I2(n4030), .O(n4031));
  LUT3 #(.INIT(8'hE8)) lut_n4032 (.I0(x1272), .I1(x1273), .I2(x1274), .O(n4032));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4033 (.I0(x1263), .I1(x1264), .I2(x1265), .I3(n4025), .I4(n4026), .O(n4033));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4034 (.I0(x1269), .I1(x1270), .I2(x1271), .I3(n4032), .I4(n4033), .O(n4034));
  LUT3 #(.INIT(8'hE8)) lut_n4035 (.I0(x1278), .I1(x1279), .I2(x1280), .O(n4035));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4036 (.I0(x1269), .I1(x1270), .I2(x1271), .I3(n4032), .I4(n4033), .O(n4036));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4037 (.I0(x1275), .I1(x1276), .I2(x1277), .I3(n4035), .I4(n4036), .O(n4037));
  LUT3 #(.INIT(8'h96)) lut_n4038 (.I0(n4024), .I1(n4027), .I2(n4028), .O(n4038));
  LUT3 #(.INIT(8'hE8)) lut_n4039 (.I0(n4034), .I1(n4037), .I2(n4038), .O(n4039));
  LUT3 #(.INIT(8'hE8)) lut_n4040 (.I0(x1284), .I1(x1285), .I2(x1286), .O(n4040));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4041 (.I0(x1275), .I1(x1276), .I2(x1277), .I3(n4035), .I4(n4036), .O(n4041));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4042 (.I0(x1281), .I1(x1282), .I2(x1283), .I3(n4040), .I4(n4041), .O(n4042));
  LUT3 #(.INIT(8'hE8)) lut_n4043 (.I0(x1290), .I1(x1291), .I2(x1292), .O(n4043));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4044 (.I0(x1281), .I1(x1282), .I2(x1283), .I3(n4040), .I4(n4041), .O(n4044));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4045 (.I0(x1287), .I1(x1288), .I2(x1289), .I3(n4043), .I4(n4044), .O(n4045));
  LUT3 #(.INIT(8'h96)) lut_n4046 (.I0(n4034), .I1(n4037), .I2(n4038), .O(n4046));
  LUT3 #(.INIT(8'hE8)) lut_n4047 (.I0(n4042), .I1(n4045), .I2(n4046), .O(n4047));
  LUT3 #(.INIT(8'h96)) lut_n4048 (.I0(n4021), .I1(n4029), .I2(n4030), .O(n4048));
  LUT3 #(.INIT(8'hE8)) lut_n4049 (.I0(n4039), .I1(n4047), .I2(n4048), .O(n4049));
  LUT3 #(.INIT(8'h96)) lut_n4050 (.I0(n3991), .I1(n4009), .I2(n4010), .O(n4050));
  LUT3 #(.INIT(8'hE8)) lut_n4051 (.I0(n4031), .I1(n4049), .I2(n4050), .O(n4051));
  LUT3 #(.INIT(8'hE8)) lut_n4052 (.I0(x1296), .I1(x1297), .I2(x1298), .O(n4052));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4053 (.I0(x1287), .I1(x1288), .I2(x1289), .I3(n4043), .I4(n4044), .O(n4053));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4054 (.I0(x1293), .I1(x1294), .I2(x1295), .I3(n4052), .I4(n4053), .O(n4054));
  LUT3 #(.INIT(8'hE8)) lut_n4055 (.I0(x1302), .I1(x1303), .I2(x1304), .O(n4055));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4056 (.I0(x1293), .I1(x1294), .I2(x1295), .I3(n4052), .I4(n4053), .O(n4056));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4057 (.I0(x1299), .I1(x1300), .I2(x1301), .I3(n4055), .I4(n4056), .O(n4057));
  LUT3 #(.INIT(8'h96)) lut_n4058 (.I0(n4042), .I1(n4045), .I2(n4046), .O(n4058));
  LUT3 #(.INIT(8'hE8)) lut_n4059 (.I0(n4054), .I1(n4057), .I2(n4058), .O(n4059));
  LUT3 #(.INIT(8'hE8)) lut_n4060 (.I0(x1308), .I1(x1309), .I2(x1310), .O(n4060));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4061 (.I0(x1299), .I1(x1300), .I2(x1301), .I3(n4055), .I4(n4056), .O(n4061));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4062 (.I0(x1305), .I1(x1306), .I2(x1307), .I3(n4060), .I4(n4061), .O(n4062));
  LUT3 #(.INIT(8'hE8)) lut_n4063 (.I0(x1314), .I1(x1315), .I2(x1316), .O(n4063));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4064 (.I0(x1305), .I1(x1306), .I2(x1307), .I3(n4060), .I4(n4061), .O(n4064));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4065 (.I0(x1311), .I1(x1312), .I2(x1313), .I3(n4063), .I4(n4064), .O(n4065));
  LUT3 #(.INIT(8'h96)) lut_n4066 (.I0(n4054), .I1(n4057), .I2(n4058), .O(n4066));
  LUT3 #(.INIT(8'hE8)) lut_n4067 (.I0(n4062), .I1(n4065), .I2(n4066), .O(n4067));
  LUT3 #(.INIT(8'h96)) lut_n4068 (.I0(n4039), .I1(n4047), .I2(n4048), .O(n4068));
  LUT3 #(.INIT(8'hE8)) lut_n4069 (.I0(n4059), .I1(n4067), .I2(n4068), .O(n4069));
  LUT3 #(.INIT(8'hE8)) lut_n4070 (.I0(x1320), .I1(x1321), .I2(x1322), .O(n4070));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4071 (.I0(x1311), .I1(x1312), .I2(x1313), .I3(n4063), .I4(n4064), .O(n4071));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4072 (.I0(x1317), .I1(x1318), .I2(x1319), .I3(n4070), .I4(n4071), .O(n4072));
  LUT3 #(.INIT(8'hE8)) lut_n4073 (.I0(x1326), .I1(x1327), .I2(x1328), .O(n4073));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4074 (.I0(x1317), .I1(x1318), .I2(x1319), .I3(n4070), .I4(n4071), .O(n4074));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4075 (.I0(x1323), .I1(x1324), .I2(x1325), .I3(n4073), .I4(n4074), .O(n4075));
  LUT3 #(.INIT(8'h96)) lut_n4076 (.I0(n4062), .I1(n4065), .I2(n4066), .O(n4076));
  LUT3 #(.INIT(8'hE8)) lut_n4077 (.I0(n4072), .I1(n4075), .I2(n4076), .O(n4077));
  LUT3 #(.INIT(8'hE8)) lut_n4078 (.I0(x1332), .I1(x1333), .I2(x1334), .O(n4078));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4079 (.I0(x1323), .I1(x1324), .I2(x1325), .I3(n4073), .I4(n4074), .O(n4079));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4080 (.I0(x1329), .I1(x1330), .I2(x1331), .I3(n4078), .I4(n4079), .O(n4080));
  LUT3 #(.INIT(8'hE8)) lut_n4081 (.I0(x1338), .I1(x1339), .I2(x1340), .O(n4081));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4082 (.I0(x1329), .I1(x1330), .I2(x1331), .I3(n4078), .I4(n4079), .O(n4082));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4083 (.I0(x1335), .I1(x1336), .I2(x1337), .I3(n4081), .I4(n4082), .O(n4083));
  LUT3 #(.INIT(8'h96)) lut_n4084 (.I0(n4072), .I1(n4075), .I2(n4076), .O(n4084));
  LUT3 #(.INIT(8'hE8)) lut_n4085 (.I0(n4080), .I1(n4083), .I2(n4084), .O(n4085));
  LUT3 #(.INIT(8'h96)) lut_n4086 (.I0(n4059), .I1(n4067), .I2(n4068), .O(n4086));
  LUT3 #(.INIT(8'hE8)) lut_n4087 (.I0(n4077), .I1(n4085), .I2(n4086), .O(n4087));
  LUT3 #(.INIT(8'h96)) lut_n4088 (.I0(n4031), .I1(n4049), .I2(n4050), .O(n4088));
  LUT3 #(.INIT(8'hE8)) lut_n4089 (.I0(n4069), .I1(n4087), .I2(n4088), .O(n4089));
  LUT3 #(.INIT(8'h96)) lut_n4090 (.I0(n3973), .I1(n4011), .I2(n4012), .O(n4090));
  LUT3 #(.INIT(8'hE8)) lut_n4091 (.I0(n4051), .I1(n4089), .I2(n4090), .O(n4091));
  LUT3 #(.INIT(8'h96)) lut_n4092 (.I0(n3853), .I1(n3931), .I2(n3932), .O(n4092));
  LUT3 #(.INIT(8'hE8)) lut_n4093 (.I0(n4013), .I1(n4091), .I2(n4092), .O(n4093));
  LUT3 #(.INIT(8'hE8)) lut_n4094 (.I0(x1344), .I1(x1345), .I2(x1346), .O(n4094));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4095 (.I0(x1335), .I1(x1336), .I2(x1337), .I3(n4081), .I4(n4082), .O(n4095));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4096 (.I0(x1341), .I1(x1342), .I2(x1343), .I3(n4094), .I4(n4095), .O(n4096));
  LUT3 #(.INIT(8'hE8)) lut_n4097 (.I0(x1350), .I1(x1351), .I2(x1352), .O(n4097));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4098 (.I0(x1341), .I1(x1342), .I2(x1343), .I3(n4094), .I4(n4095), .O(n4098));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4099 (.I0(x1347), .I1(x1348), .I2(x1349), .I3(n4097), .I4(n4098), .O(n4099));
  LUT3 #(.INIT(8'h96)) lut_n4100 (.I0(n4080), .I1(n4083), .I2(n4084), .O(n4100));
  LUT3 #(.INIT(8'hE8)) lut_n4101 (.I0(n4096), .I1(n4099), .I2(n4100), .O(n4101));
  LUT3 #(.INIT(8'hE8)) lut_n4102 (.I0(x1356), .I1(x1357), .I2(x1358), .O(n4102));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4103 (.I0(x1347), .I1(x1348), .I2(x1349), .I3(n4097), .I4(n4098), .O(n4103));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4104 (.I0(x1353), .I1(x1354), .I2(x1355), .I3(n4102), .I4(n4103), .O(n4104));
  LUT3 #(.INIT(8'hE8)) lut_n4105 (.I0(x1362), .I1(x1363), .I2(x1364), .O(n4105));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4106 (.I0(x1353), .I1(x1354), .I2(x1355), .I3(n4102), .I4(n4103), .O(n4106));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4107 (.I0(x1359), .I1(x1360), .I2(x1361), .I3(n4105), .I4(n4106), .O(n4107));
  LUT3 #(.INIT(8'h96)) lut_n4108 (.I0(n4096), .I1(n4099), .I2(n4100), .O(n4108));
  LUT3 #(.INIT(8'hE8)) lut_n4109 (.I0(n4104), .I1(n4107), .I2(n4108), .O(n4109));
  LUT3 #(.INIT(8'h96)) lut_n4110 (.I0(n4077), .I1(n4085), .I2(n4086), .O(n4110));
  LUT3 #(.INIT(8'hE8)) lut_n4111 (.I0(n4101), .I1(n4109), .I2(n4110), .O(n4111));
  LUT3 #(.INIT(8'hE8)) lut_n4112 (.I0(x1368), .I1(x1369), .I2(x1370), .O(n4112));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4113 (.I0(x1359), .I1(x1360), .I2(x1361), .I3(n4105), .I4(n4106), .O(n4113));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4114 (.I0(x1365), .I1(x1366), .I2(x1367), .I3(n4112), .I4(n4113), .O(n4114));
  LUT3 #(.INIT(8'hE8)) lut_n4115 (.I0(x1374), .I1(x1375), .I2(x1376), .O(n4115));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4116 (.I0(x1365), .I1(x1366), .I2(x1367), .I3(n4112), .I4(n4113), .O(n4116));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4117 (.I0(x1371), .I1(x1372), .I2(x1373), .I3(n4115), .I4(n4116), .O(n4117));
  LUT3 #(.INIT(8'h96)) lut_n4118 (.I0(n4104), .I1(n4107), .I2(n4108), .O(n4118));
  LUT3 #(.INIT(8'hE8)) lut_n4119 (.I0(n4114), .I1(n4117), .I2(n4118), .O(n4119));
  LUT3 #(.INIT(8'hE8)) lut_n4120 (.I0(x1380), .I1(x1381), .I2(x1382), .O(n4120));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4121 (.I0(x1371), .I1(x1372), .I2(x1373), .I3(n4115), .I4(n4116), .O(n4121));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4122 (.I0(x1377), .I1(x1378), .I2(x1379), .I3(n4120), .I4(n4121), .O(n4122));
  LUT3 #(.INIT(8'hE8)) lut_n4123 (.I0(x1386), .I1(x1387), .I2(x1388), .O(n4123));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4124 (.I0(x1377), .I1(x1378), .I2(x1379), .I3(n4120), .I4(n4121), .O(n4124));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4125 (.I0(x1383), .I1(x1384), .I2(x1385), .I3(n4123), .I4(n4124), .O(n4125));
  LUT3 #(.INIT(8'h96)) lut_n4126 (.I0(n4114), .I1(n4117), .I2(n4118), .O(n4126));
  LUT3 #(.INIT(8'hE8)) lut_n4127 (.I0(n4122), .I1(n4125), .I2(n4126), .O(n4127));
  LUT3 #(.INIT(8'h96)) lut_n4128 (.I0(n4101), .I1(n4109), .I2(n4110), .O(n4128));
  LUT3 #(.INIT(8'hE8)) lut_n4129 (.I0(n4119), .I1(n4127), .I2(n4128), .O(n4129));
  LUT3 #(.INIT(8'h96)) lut_n4130 (.I0(n4069), .I1(n4087), .I2(n4088), .O(n4130));
  LUT3 #(.INIT(8'hE8)) lut_n4131 (.I0(n4111), .I1(n4129), .I2(n4130), .O(n4131));
  LUT3 #(.INIT(8'hE8)) lut_n4132 (.I0(x1392), .I1(x1393), .I2(x1394), .O(n4132));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4133 (.I0(x1383), .I1(x1384), .I2(x1385), .I3(n4123), .I4(n4124), .O(n4133));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4134 (.I0(x1389), .I1(x1390), .I2(x1391), .I3(n4132), .I4(n4133), .O(n4134));
  LUT3 #(.INIT(8'hE8)) lut_n4135 (.I0(x1398), .I1(x1399), .I2(x1400), .O(n4135));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4136 (.I0(x1389), .I1(x1390), .I2(x1391), .I3(n4132), .I4(n4133), .O(n4136));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4137 (.I0(x1395), .I1(x1396), .I2(x1397), .I3(n4135), .I4(n4136), .O(n4137));
  LUT3 #(.INIT(8'h96)) lut_n4138 (.I0(n4122), .I1(n4125), .I2(n4126), .O(n4138));
  LUT3 #(.INIT(8'hE8)) lut_n4139 (.I0(n4134), .I1(n4137), .I2(n4138), .O(n4139));
  LUT3 #(.INIT(8'hE8)) lut_n4140 (.I0(x1404), .I1(x1405), .I2(x1406), .O(n4140));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4141 (.I0(x1395), .I1(x1396), .I2(x1397), .I3(n4135), .I4(n4136), .O(n4141));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4142 (.I0(x1401), .I1(x1402), .I2(x1403), .I3(n4140), .I4(n4141), .O(n4142));
  LUT3 #(.INIT(8'hE8)) lut_n4143 (.I0(x1410), .I1(x1411), .I2(x1412), .O(n4143));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4144 (.I0(x1401), .I1(x1402), .I2(x1403), .I3(n4140), .I4(n4141), .O(n4144));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4145 (.I0(x1407), .I1(x1408), .I2(x1409), .I3(n4143), .I4(n4144), .O(n4145));
  LUT3 #(.INIT(8'h96)) lut_n4146 (.I0(n4134), .I1(n4137), .I2(n4138), .O(n4146));
  LUT3 #(.INIT(8'hE8)) lut_n4147 (.I0(n4142), .I1(n4145), .I2(n4146), .O(n4147));
  LUT3 #(.INIT(8'h96)) lut_n4148 (.I0(n4119), .I1(n4127), .I2(n4128), .O(n4148));
  LUT3 #(.INIT(8'hE8)) lut_n4149 (.I0(n4139), .I1(n4147), .I2(n4148), .O(n4149));
  LUT3 #(.INIT(8'hE8)) lut_n4150 (.I0(x1416), .I1(x1417), .I2(x1418), .O(n4150));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4151 (.I0(x1407), .I1(x1408), .I2(x1409), .I3(n4143), .I4(n4144), .O(n4151));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4152 (.I0(x1413), .I1(x1414), .I2(x1415), .I3(n4150), .I4(n4151), .O(n4152));
  LUT3 #(.INIT(8'hE8)) lut_n4153 (.I0(x1422), .I1(x1423), .I2(x1424), .O(n4153));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4154 (.I0(x1413), .I1(x1414), .I2(x1415), .I3(n4150), .I4(n4151), .O(n4154));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4155 (.I0(x1419), .I1(x1420), .I2(x1421), .I3(n4153), .I4(n4154), .O(n4155));
  LUT3 #(.INIT(8'h96)) lut_n4156 (.I0(n4142), .I1(n4145), .I2(n4146), .O(n4156));
  LUT3 #(.INIT(8'hE8)) lut_n4157 (.I0(n4152), .I1(n4155), .I2(n4156), .O(n4157));
  LUT3 #(.INIT(8'hE8)) lut_n4158 (.I0(x1428), .I1(x1429), .I2(x1430), .O(n4158));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4159 (.I0(x1419), .I1(x1420), .I2(x1421), .I3(n4153), .I4(n4154), .O(n4159));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4160 (.I0(x1425), .I1(x1426), .I2(x1427), .I3(n4158), .I4(n4159), .O(n4160));
  LUT3 #(.INIT(8'hE8)) lut_n4161 (.I0(x1434), .I1(x1435), .I2(x1436), .O(n4161));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4162 (.I0(x1425), .I1(x1426), .I2(x1427), .I3(n4158), .I4(n4159), .O(n4162));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4163 (.I0(x1431), .I1(x1432), .I2(x1433), .I3(n4161), .I4(n4162), .O(n4163));
  LUT3 #(.INIT(8'h96)) lut_n4164 (.I0(n4152), .I1(n4155), .I2(n4156), .O(n4164));
  LUT3 #(.INIT(8'hE8)) lut_n4165 (.I0(n4160), .I1(n4163), .I2(n4164), .O(n4165));
  LUT3 #(.INIT(8'h96)) lut_n4166 (.I0(n4139), .I1(n4147), .I2(n4148), .O(n4166));
  LUT3 #(.INIT(8'hE8)) lut_n4167 (.I0(n4157), .I1(n4165), .I2(n4166), .O(n4167));
  LUT3 #(.INIT(8'h96)) lut_n4168 (.I0(n4111), .I1(n4129), .I2(n4130), .O(n4168));
  LUT3 #(.INIT(8'hE8)) lut_n4169 (.I0(n4149), .I1(n4167), .I2(n4168), .O(n4169));
  LUT3 #(.INIT(8'h96)) lut_n4170 (.I0(n4051), .I1(n4089), .I2(n4090), .O(n4170));
  LUT3 #(.INIT(8'hE8)) lut_n4171 (.I0(n4131), .I1(n4169), .I2(n4170), .O(n4171));
  LUT3 #(.INIT(8'hE8)) lut_n4172 (.I0(x1440), .I1(x1441), .I2(x1442), .O(n4172));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4173 (.I0(x1431), .I1(x1432), .I2(x1433), .I3(n4161), .I4(n4162), .O(n4173));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4174 (.I0(x1437), .I1(x1438), .I2(x1439), .I3(n4172), .I4(n4173), .O(n4174));
  LUT3 #(.INIT(8'hE8)) lut_n4175 (.I0(x1446), .I1(x1447), .I2(x1448), .O(n4175));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4176 (.I0(x1437), .I1(x1438), .I2(x1439), .I3(n4172), .I4(n4173), .O(n4176));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4177 (.I0(x1443), .I1(x1444), .I2(x1445), .I3(n4175), .I4(n4176), .O(n4177));
  LUT3 #(.INIT(8'h96)) lut_n4178 (.I0(n4160), .I1(n4163), .I2(n4164), .O(n4178));
  LUT3 #(.INIT(8'hE8)) lut_n4179 (.I0(n4174), .I1(n4177), .I2(n4178), .O(n4179));
  LUT3 #(.INIT(8'hE8)) lut_n4180 (.I0(x1452), .I1(x1453), .I2(x1454), .O(n4180));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4181 (.I0(x1443), .I1(x1444), .I2(x1445), .I3(n4175), .I4(n4176), .O(n4181));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4182 (.I0(x1449), .I1(x1450), .I2(x1451), .I3(n4180), .I4(n4181), .O(n4182));
  LUT3 #(.INIT(8'hE8)) lut_n4183 (.I0(x1458), .I1(x1459), .I2(x1460), .O(n4183));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4184 (.I0(x1449), .I1(x1450), .I2(x1451), .I3(n4180), .I4(n4181), .O(n4184));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4185 (.I0(x1455), .I1(x1456), .I2(x1457), .I3(n4183), .I4(n4184), .O(n4185));
  LUT3 #(.INIT(8'h96)) lut_n4186 (.I0(n4174), .I1(n4177), .I2(n4178), .O(n4186));
  LUT3 #(.INIT(8'hE8)) lut_n4187 (.I0(n4182), .I1(n4185), .I2(n4186), .O(n4187));
  LUT3 #(.INIT(8'h96)) lut_n4188 (.I0(n4157), .I1(n4165), .I2(n4166), .O(n4188));
  LUT3 #(.INIT(8'hE8)) lut_n4189 (.I0(n4179), .I1(n4187), .I2(n4188), .O(n4189));
  LUT3 #(.INIT(8'hE8)) lut_n4190 (.I0(x1464), .I1(x1465), .I2(x1466), .O(n4190));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4191 (.I0(x1455), .I1(x1456), .I2(x1457), .I3(n4183), .I4(n4184), .O(n4191));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4192 (.I0(x1461), .I1(x1462), .I2(x1463), .I3(n4190), .I4(n4191), .O(n4192));
  LUT3 #(.INIT(8'hE8)) lut_n4193 (.I0(x1470), .I1(x1471), .I2(x1472), .O(n4193));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4194 (.I0(x1461), .I1(x1462), .I2(x1463), .I3(n4190), .I4(n4191), .O(n4194));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4195 (.I0(x1467), .I1(x1468), .I2(x1469), .I3(n4193), .I4(n4194), .O(n4195));
  LUT3 #(.INIT(8'h96)) lut_n4196 (.I0(n4182), .I1(n4185), .I2(n4186), .O(n4196));
  LUT3 #(.INIT(8'hE8)) lut_n4197 (.I0(n4192), .I1(n4195), .I2(n4196), .O(n4197));
  LUT3 #(.INIT(8'hE8)) lut_n4198 (.I0(x1476), .I1(x1477), .I2(x1478), .O(n4198));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4199 (.I0(x1467), .I1(x1468), .I2(x1469), .I3(n4193), .I4(n4194), .O(n4199));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4200 (.I0(x1473), .I1(x1474), .I2(x1475), .I3(n4198), .I4(n4199), .O(n4200));
  LUT3 #(.INIT(8'hE8)) lut_n4201 (.I0(x1482), .I1(x1483), .I2(x1484), .O(n4201));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4202 (.I0(x1473), .I1(x1474), .I2(x1475), .I3(n4198), .I4(n4199), .O(n4202));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4203 (.I0(x1479), .I1(x1480), .I2(x1481), .I3(n4201), .I4(n4202), .O(n4203));
  LUT3 #(.INIT(8'h96)) lut_n4204 (.I0(n4192), .I1(n4195), .I2(n4196), .O(n4204));
  LUT3 #(.INIT(8'hE8)) lut_n4205 (.I0(n4200), .I1(n4203), .I2(n4204), .O(n4205));
  LUT3 #(.INIT(8'h96)) lut_n4206 (.I0(n4179), .I1(n4187), .I2(n4188), .O(n4206));
  LUT3 #(.INIT(8'hE8)) lut_n4207 (.I0(n4197), .I1(n4205), .I2(n4206), .O(n4207));
  LUT3 #(.INIT(8'h96)) lut_n4208 (.I0(n4149), .I1(n4167), .I2(n4168), .O(n4208));
  LUT3 #(.INIT(8'hE8)) lut_n4209 (.I0(n4189), .I1(n4207), .I2(n4208), .O(n4209));
  LUT3 #(.INIT(8'hE8)) lut_n4210 (.I0(x1488), .I1(x1489), .I2(x1490), .O(n4210));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4211 (.I0(x1479), .I1(x1480), .I2(x1481), .I3(n4201), .I4(n4202), .O(n4211));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4212 (.I0(x1485), .I1(x1486), .I2(x1487), .I3(n4210), .I4(n4211), .O(n4212));
  LUT3 #(.INIT(8'hE8)) lut_n4213 (.I0(x1494), .I1(x1495), .I2(x1496), .O(n4213));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4214 (.I0(x1485), .I1(x1486), .I2(x1487), .I3(n4210), .I4(n4211), .O(n4214));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4215 (.I0(x1491), .I1(x1492), .I2(x1493), .I3(n4213), .I4(n4214), .O(n4215));
  LUT3 #(.INIT(8'h96)) lut_n4216 (.I0(n4200), .I1(n4203), .I2(n4204), .O(n4216));
  LUT3 #(.INIT(8'hE8)) lut_n4217 (.I0(n4212), .I1(n4215), .I2(n4216), .O(n4217));
  LUT3 #(.INIT(8'hE8)) lut_n4218 (.I0(x1500), .I1(x1501), .I2(x1502), .O(n4218));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4219 (.I0(x1491), .I1(x1492), .I2(x1493), .I3(n4213), .I4(n4214), .O(n4219));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4220 (.I0(x1497), .I1(x1498), .I2(x1499), .I3(n4218), .I4(n4219), .O(n4220));
  LUT3 #(.INIT(8'hE8)) lut_n4221 (.I0(x1506), .I1(x1507), .I2(x1508), .O(n4221));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4222 (.I0(x1497), .I1(x1498), .I2(x1499), .I3(n4218), .I4(n4219), .O(n4222));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4223 (.I0(x1503), .I1(x1504), .I2(x1505), .I3(n4221), .I4(n4222), .O(n4223));
  LUT3 #(.INIT(8'h96)) lut_n4224 (.I0(n4212), .I1(n4215), .I2(n4216), .O(n4224));
  LUT3 #(.INIT(8'hE8)) lut_n4225 (.I0(n4220), .I1(n4223), .I2(n4224), .O(n4225));
  LUT3 #(.INIT(8'h96)) lut_n4226 (.I0(n4197), .I1(n4205), .I2(n4206), .O(n4226));
  LUT3 #(.INIT(8'hE8)) lut_n4227 (.I0(n4217), .I1(n4225), .I2(n4226), .O(n4227));
  LUT3 #(.INIT(8'hE8)) lut_n4228 (.I0(x1512), .I1(x1513), .I2(x1514), .O(n4228));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4229 (.I0(x1503), .I1(x1504), .I2(x1505), .I3(n4221), .I4(n4222), .O(n4229));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4230 (.I0(x1509), .I1(x1510), .I2(x1511), .I3(n4228), .I4(n4229), .O(n4230));
  LUT3 #(.INIT(8'hE8)) lut_n4231 (.I0(x1518), .I1(x1519), .I2(x1520), .O(n4231));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4232 (.I0(x1509), .I1(x1510), .I2(x1511), .I3(n4228), .I4(n4229), .O(n4232));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4233 (.I0(x1515), .I1(x1516), .I2(x1517), .I3(n4231), .I4(n4232), .O(n4233));
  LUT3 #(.INIT(8'h96)) lut_n4234 (.I0(n4220), .I1(n4223), .I2(n4224), .O(n4234));
  LUT3 #(.INIT(8'hE8)) lut_n4235 (.I0(n4230), .I1(n4233), .I2(n4234), .O(n4235));
  LUT3 #(.INIT(8'hE8)) lut_n4236 (.I0(x1524), .I1(x1525), .I2(x1526), .O(n4236));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4237 (.I0(x1515), .I1(x1516), .I2(x1517), .I3(n4231), .I4(n4232), .O(n4237));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4238 (.I0(x1521), .I1(x1522), .I2(x1523), .I3(n4236), .I4(n4237), .O(n4238));
  LUT3 #(.INIT(8'hE8)) lut_n4239 (.I0(x1530), .I1(x1531), .I2(x1532), .O(n4239));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4240 (.I0(x1521), .I1(x1522), .I2(x1523), .I3(n4236), .I4(n4237), .O(n4240));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4241 (.I0(x1527), .I1(x1528), .I2(x1529), .I3(n4239), .I4(n4240), .O(n4241));
  LUT3 #(.INIT(8'h96)) lut_n4242 (.I0(n4230), .I1(n4233), .I2(n4234), .O(n4242));
  LUT3 #(.INIT(8'hE8)) lut_n4243 (.I0(n4238), .I1(n4241), .I2(n4242), .O(n4243));
  LUT3 #(.INIT(8'h96)) lut_n4244 (.I0(n4217), .I1(n4225), .I2(n4226), .O(n4244));
  LUT3 #(.INIT(8'hE8)) lut_n4245 (.I0(n4235), .I1(n4243), .I2(n4244), .O(n4245));
  LUT3 #(.INIT(8'h96)) lut_n4246 (.I0(n4189), .I1(n4207), .I2(n4208), .O(n4246));
  LUT3 #(.INIT(8'hE8)) lut_n4247 (.I0(n4227), .I1(n4245), .I2(n4246), .O(n4247));
  LUT3 #(.INIT(8'h96)) lut_n4248 (.I0(n4131), .I1(n4169), .I2(n4170), .O(n4248));
  LUT3 #(.INIT(8'hE8)) lut_n4249 (.I0(n4209), .I1(n4247), .I2(n4248), .O(n4249));
  LUT3 #(.INIT(8'h96)) lut_n4250 (.I0(n4013), .I1(n4091), .I2(n4092), .O(n4250));
  LUT3 #(.INIT(8'hE8)) lut_n4251 (.I0(n4171), .I1(n4249), .I2(n4250), .O(n4251));
  LUT3 #(.INIT(8'h96)) lut_n4252 (.I0(n3775), .I1(n3933), .I2(n3934), .O(n4252));
  LUT3 #(.INIT(8'hE8)) lut_n4253 (.I0(n4093), .I1(n4251), .I2(n4252), .O(n4253));
  LUT3 #(.INIT(8'hE8)) lut_n4254 (.I0(n3617), .I1(n3935), .I2(n4253), .O(n4254));
  LUT3 #(.INIT(8'hE8)) lut_n4255 (.I0(x1536), .I1(x1537), .I2(x1538), .O(n4255));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4256 (.I0(x1527), .I1(x1528), .I2(x1529), .I3(n4239), .I4(n4240), .O(n4256));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4257 (.I0(x1533), .I1(x1534), .I2(x1535), .I3(n4255), .I4(n4256), .O(n4257));
  LUT3 #(.INIT(8'hE8)) lut_n4258 (.I0(x1542), .I1(x1543), .I2(x1544), .O(n4258));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4259 (.I0(x1533), .I1(x1534), .I2(x1535), .I3(n4255), .I4(n4256), .O(n4259));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4260 (.I0(x1539), .I1(x1540), .I2(x1541), .I3(n4258), .I4(n4259), .O(n4260));
  LUT3 #(.INIT(8'h96)) lut_n4261 (.I0(n4238), .I1(n4241), .I2(n4242), .O(n4261));
  LUT3 #(.INIT(8'hE8)) lut_n4262 (.I0(n4257), .I1(n4260), .I2(n4261), .O(n4262));
  LUT3 #(.INIT(8'hE8)) lut_n4263 (.I0(x1548), .I1(x1549), .I2(x1550), .O(n4263));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4264 (.I0(x1539), .I1(x1540), .I2(x1541), .I3(n4258), .I4(n4259), .O(n4264));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4265 (.I0(x1545), .I1(x1546), .I2(x1547), .I3(n4263), .I4(n4264), .O(n4265));
  LUT3 #(.INIT(8'hE8)) lut_n4266 (.I0(x1554), .I1(x1555), .I2(x1556), .O(n4266));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4267 (.I0(x1545), .I1(x1546), .I2(x1547), .I3(n4263), .I4(n4264), .O(n4267));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4268 (.I0(x1551), .I1(x1552), .I2(x1553), .I3(n4266), .I4(n4267), .O(n4268));
  LUT3 #(.INIT(8'h96)) lut_n4269 (.I0(n4257), .I1(n4260), .I2(n4261), .O(n4269));
  LUT3 #(.INIT(8'hE8)) lut_n4270 (.I0(n4265), .I1(n4268), .I2(n4269), .O(n4270));
  LUT3 #(.INIT(8'h96)) lut_n4271 (.I0(n4235), .I1(n4243), .I2(n4244), .O(n4271));
  LUT3 #(.INIT(8'hE8)) lut_n4272 (.I0(n4262), .I1(n4270), .I2(n4271), .O(n4272));
  LUT3 #(.INIT(8'hE8)) lut_n4273 (.I0(x1560), .I1(x1561), .I2(x1562), .O(n4273));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4274 (.I0(x1551), .I1(x1552), .I2(x1553), .I3(n4266), .I4(n4267), .O(n4274));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4275 (.I0(x1557), .I1(x1558), .I2(x1559), .I3(n4273), .I4(n4274), .O(n4275));
  LUT3 #(.INIT(8'hE8)) lut_n4276 (.I0(x1566), .I1(x1567), .I2(x1568), .O(n4276));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4277 (.I0(x1557), .I1(x1558), .I2(x1559), .I3(n4273), .I4(n4274), .O(n4277));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4278 (.I0(x1563), .I1(x1564), .I2(x1565), .I3(n4276), .I4(n4277), .O(n4278));
  LUT3 #(.INIT(8'h96)) lut_n4279 (.I0(n4265), .I1(n4268), .I2(n4269), .O(n4279));
  LUT3 #(.INIT(8'hE8)) lut_n4280 (.I0(n4275), .I1(n4278), .I2(n4279), .O(n4280));
  LUT3 #(.INIT(8'hE8)) lut_n4281 (.I0(x1572), .I1(x1573), .I2(x1574), .O(n4281));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4282 (.I0(x1563), .I1(x1564), .I2(x1565), .I3(n4276), .I4(n4277), .O(n4282));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4283 (.I0(x1569), .I1(x1570), .I2(x1571), .I3(n4281), .I4(n4282), .O(n4283));
  LUT3 #(.INIT(8'hE8)) lut_n4284 (.I0(x1578), .I1(x1579), .I2(x1580), .O(n4284));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4285 (.I0(x1569), .I1(x1570), .I2(x1571), .I3(n4281), .I4(n4282), .O(n4285));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4286 (.I0(x1575), .I1(x1576), .I2(x1577), .I3(n4284), .I4(n4285), .O(n4286));
  LUT3 #(.INIT(8'h96)) lut_n4287 (.I0(n4275), .I1(n4278), .I2(n4279), .O(n4287));
  LUT3 #(.INIT(8'hE8)) lut_n4288 (.I0(n4283), .I1(n4286), .I2(n4287), .O(n4288));
  LUT3 #(.INIT(8'h96)) lut_n4289 (.I0(n4262), .I1(n4270), .I2(n4271), .O(n4289));
  LUT3 #(.INIT(8'hE8)) lut_n4290 (.I0(n4280), .I1(n4288), .I2(n4289), .O(n4290));
  LUT3 #(.INIT(8'h96)) lut_n4291 (.I0(n4227), .I1(n4245), .I2(n4246), .O(n4291));
  LUT3 #(.INIT(8'hE8)) lut_n4292 (.I0(n4272), .I1(n4290), .I2(n4291), .O(n4292));
  LUT3 #(.INIT(8'hE8)) lut_n4293 (.I0(x1584), .I1(x1585), .I2(x1586), .O(n4293));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4294 (.I0(x1575), .I1(x1576), .I2(x1577), .I3(n4284), .I4(n4285), .O(n4294));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4295 (.I0(x1581), .I1(x1582), .I2(x1583), .I3(n4293), .I4(n4294), .O(n4295));
  LUT3 #(.INIT(8'hE8)) lut_n4296 (.I0(x1590), .I1(x1591), .I2(x1592), .O(n4296));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4297 (.I0(x1581), .I1(x1582), .I2(x1583), .I3(n4293), .I4(n4294), .O(n4297));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4298 (.I0(x1587), .I1(x1588), .I2(x1589), .I3(n4296), .I4(n4297), .O(n4298));
  LUT3 #(.INIT(8'h96)) lut_n4299 (.I0(n4283), .I1(n4286), .I2(n4287), .O(n4299));
  LUT3 #(.INIT(8'hE8)) lut_n4300 (.I0(n4295), .I1(n4298), .I2(n4299), .O(n4300));
  LUT3 #(.INIT(8'hE8)) lut_n4301 (.I0(x1596), .I1(x1597), .I2(x1598), .O(n4301));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4302 (.I0(x1587), .I1(x1588), .I2(x1589), .I3(n4296), .I4(n4297), .O(n4302));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4303 (.I0(x1593), .I1(x1594), .I2(x1595), .I3(n4301), .I4(n4302), .O(n4303));
  LUT3 #(.INIT(8'hE8)) lut_n4304 (.I0(x1602), .I1(x1603), .I2(x1604), .O(n4304));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4305 (.I0(x1593), .I1(x1594), .I2(x1595), .I3(n4301), .I4(n4302), .O(n4305));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4306 (.I0(x1599), .I1(x1600), .I2(x1601), .I3(n4304), .I4(n4305), .O(n4306));
  LUT3 #(.INIT(8'h96)) lut_n4307 (.I0(n4295), .I1(n4298), .I2(n4299), .O(n4307));
  LUT3 #(.INIT(8'hE8)) lut_n4308 (.I0(n4303), .I1(n4306), .I2(n4307), .O(n4308));
  LUT3 #(.INIT(8'h96)) lut_n4309 (.I0(n4280), .I1(n4288), .I2(n4289), .O(n4309));
  LUT3 #(.INIT(8'hE8)) lut_n4310 (.I0(n4300), .I1(n4308), .I2(n4309), .O(n4310));
  LUT3 #(.INIT(8'hE8)) lut_n4311 (.I0(x1608), .I1(x1609), .I2(x1610), .O(n4311));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4312 (.I0(x1599), .I1(x1600), .I2(x1601), .I3(n4304), .I4(n4305), .O(n4312));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4313 (.I0(x1605), .I1(x1606), .I2(x1607), .I3(n4311), .I4(n4312), .O(n4313));
  LUT3 #(.INIT(8'hE8)) lut_n4314 (.I0(x1614), .I1(x1615), .I2(x1616), .O(n4314));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4315 (.I0(x1605), .I1(x1606), .I2(x1607), .I3(n4311), .I4(n4312), .O(n4315));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4316 (.I0(x1611), .I1(x1612), .I2(x1613), .I3(n4314), .I4(n4315), .O(n4316));
  LUT3 #(.INIT(8'h96)) lut_n4317 (.I0(n4303), .I1(n4306), .I2(n4307), .O(n4317));
  LUT3 #(.INIT(8'hE8)) lut_n4318 (.I0(n4313), .I1(n4316), .I2(n4317), .O(n4318));
  LUT3 #(.INIT(8'hE8)) lut_n4319 (.I0(x1620), .I1(x1621), .I2(x1622), .O(n4319));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4320 (.I0(x1611), .I1(x1612), .I2(x1613), .I3(n4314), .I4(n4315), .O(n4320));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4321 (.I0(x1617), .I1(x1618), .I2(x1619), .I3(n4319), .I4(n4320), .O(n4321));
  LUT3 #(.INIT(8'hE8)) lut_n4322 (.I0(x1626), .I1(x1627), .I2(x1628), .O(n4322));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4323 (.I0(x1617), .I1(x1618), .I2(x1619), .I3(n4319), .I4(n4320), .O(n4323));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4324 (.I0(x1623), .I1(x1624), .I2(x1625), .I3(n4322), .I4(n4323), .O(n4324));
  LUT3 #(.INIT(8'h96)) lut_n4325 (.I0(n4313), .I1(n4316), .I2(n4317), .O(n4325));
  LUT3 #(.INIT(8'hE8)) lut_n4326 (.I0(n4321), .I1(n4324), .I2(n4325), .O(n4326));
  LUT3 #(.INIT(8'h96)) lut_n4327 (.I0(n4300), .I1(n4308), .I2(n4309), .O(n4327));
  LUT3 #(.INIT(8'hE8)) lut_n4328 (.I0(n4318), .I1(n4326), .I2(n4327), .O(n4328));
  LUT3 #(.INIT(8'h96)) lut_n4329 (.I0(n4272), .I1(n4290), .I2(n4291), .O(n4329));
  LUT3 #(.INIT(8'hE8)) lut_n4330 (.I0(n4310), .I1(n4328), .I2(n4329), .O(n4330));
  LUT3 #(.INIT(8'h96)) lut_n4331 (.I0(n4209), .I1(n4247), .I2(n4248), .O(n4331));
  LUT3 #(.INIT(8'hE8)) lut_n4332 (.I0(n4292), .I1(n4330), .I2(n4331), .O(n4332));
  LUT3 #(.INIT(8'hE8)) lut_n4333 (.I0(x1632), .I1(x1633), .I2(x1634), .O(n4333));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4334 (.I0(x1623), .I1(x1624), .I2(x1625), .I3(n4322), .I4(n4323), .O(n4334));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4335 (.I0(x1629), .I1(x1630), .I2(x1631), .I3(n4333), .I4(n4334), .O(n4335));
  LUT3 #(.INIT(8'hE8)) lut_n4336 (.I0(x1638), .I1(x1639), .I2(x1640), .O(n4336));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4337 (.I0(x1629), .I1(x1630), .I2(x1631), .I3(n4333), .I4(n4334), .O(n4337));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4338 (.I0(x1635), .I1(x1636), .I2(x1637), .I3(n4336), .I4(n4337), .O(n4338));
  LUT3 #(.INIT(8'h96)) lut_n4339 (.I0(n4321), .I1(n4324), .I2(n4325), .O(n4339));
  LUT3 #(.INIT(8'hE8)) lut_n4340 (.I0(n4335), .I1(n4338), .I2(n4339), .O(n4340));
  LUT3 #(.INIT(8'hE8)) lut_n4341 (.I0(x1644), .I1(x1645), .I2(x1646), .O(n4341));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4342 (.I0(x1635), .I1(x1636), .I2(x1637), .I3(n4336), .I4(n4337), .O(n4342));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4343 (.I0(x1641), .I1(x1642), .I2(x1643), .I3(n4341), .I4(n4342), .O(n4343));
  LUT3 #(.INIT(8'hE8)) lut_n4344 (.I0(x1650), .I1(x1651), .I2(x1652), .O(n4344));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4345 (.I0(x1641), .I1(x1642), .I2(x1643), .I3(n4341), .I4(n4342), .O(n4345));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4346 (.I0(x1647), .I1(x1648), .I2(x1649), .I3(n4344), .I4(n4345), .O(n4346));
  LUT3 #(.INIT(8'h96)) lut_n4347 (.I0(n4335), .I1(n4338), .I2(n4339), .O(n4347));
  LUT3 #(.INIT(8'hE8)) lut_n4348 (.I0(n4343), .I1(n4346), .I2(n4347), .O(n4348));
  LUT3 #(.INIT(8'h96)) lut_n4349 (.I0(n4318), .I1(n4326), .I2(n4327), .O(n4349));
  LUT3 #(.INIT(8'hE8)) lut_n4350 (.I0(n4340), .I1(n4348), .I2(n4349), .O(n4350));
  LUT3 #(.INIT(8'hE8)) lut_n4351 (.I0(x1656), .I1(x1657), .I2(x1658), .O(n4351));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4352 (.I0(x1647), .I1(x1648), .I2(x1649), .I3(n4344), .I4(n4345), .O(n4352));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4353 (.I0(x1653), .I1(x1654), .I2(x1655), .I3(n4351), .I4(n4352), .O(n4353));
  LUT3 #(.INIT(8'hE8)) lut_n4354 (.I0(x1662), .I1(x1663), .I2(x1664), .O(n4354));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4355 (.I0(x1653), .I1(x1654), .I2(x1655), .I3(n4351), .I4(n4352), .O(n4355));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4356 (.I0(x1659), .I1(x1660), .I2(x1661), .I3(n4354), .I4(n4355), .O(n4356));
  LUT3 #(.INIT(8'h96)) lut_n4357 (.I0(n4343), .I1(n4346), .I2(n4347), .O(n4357));
  LUT3 #(.INIT(8'hE8)) lut_n4358 (.I0(n4353), .I1(n4356), .I2(n4357), .O(n4358));
  LUT3 #(.INIT(8'hE8)) lut_n4359 (.I0(x1668), .I1(x1669), .I2(x1670), .O(n4359));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4360 (.I0(x1659), .I1(x1660), .I2(x1661), .I3(n4354), .I4(n4355), .O(n4360));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4361 (.I0(x1665), .I1(x1666), .I2(x1667), .I3(n4359), .I4(n4360), .O(n4361));
  LUT3 #(.INIT(8'hE8)) lut_n4362 (.I0(x1674), .I1(x1675), .I2(x1676), .O(n4362));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4363 (.I0(x1665), .I1(x1666), .I2(x1667), .I3(n4359), .I4(n4360), .O(n4363));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4364 (.I0(x1671), .I1(x1672), .I2(x1673), .I3(n4362), .I4(n4363), .O(n4364));
  LUT3 #(.INIT(8'h96)) lut_n4365 (.I0(n4353), .I1(n4356), .I2(n4357), .O(n4365));
  LUT3 #(.INIT(8'hE8)) lut_n4366 (.I0(n4361), .I1(n4364), .I2(n4365), .O(n4366));
  LUT3 #(.INIT(8'h96)) lut_n4367 (.I0(n4340), .I1(n4348), .I2(n4349), .O(n4367));
  LUT3 #(.INIT(8'hE8)) lut_n4368 (.I0(n4358), .I1(n4366), .I2(n4367), .O(n4368));
  LUT3 #(.INIT(8'h96)) lut_n4369 (.I0(n4310), .I1(n4328), .I2(n4329), .O(n4369));
  LUT3 #(.INIT(8'hE8)) lut_n4370 (.I0(n4350), .I1(n4368), .I2(n4369), .O(n4370));
  LUT3 #(.INIT(8'hE8)) lut_n4371 (.I0(x1680), .I1(x1681), .I2(x1682), .O(n4371));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4372 (.I0(x1671), .I1(x1672), .I2(x1673), .I3(n4362), .I4(n4363), .O(n4372));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4373 (.I0(x1677), .I1(x1678), .I2(x1679), .I3(n4371), .I4(n4372), .O(n4373));
  LUT3 #(.INIT(8'hE8)) lut_n4374 (.I0(x1686), .I1(x1687), .I2(x1688), .O(n4374));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4375 (.I0(x1677), .I1(x1678), .I2(x1679), .I3(n4371), .I4(n4372), .O(n4375));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4376 (.I0(x1683), .I1(x1684), .I2(x1685), .I3(n4374), .I4(n4375), .O(n4376));
  LUT3 #(.INIT(8'h96)) lut_n4377 (.I0(n4361), .I1(n4364), .I2(n4365), .O(n4377));
  LUT3 #(.INIT(8'hE8)) lut_n4378 (.I0(n4373), .I1(n4376), .I2(n4377), .O(n4378));
  LUT3 #(.INIT(8'hE8)) lut_n4379 (.I0(x1692), .I1(x1693), .I2(x1694), .O(n4379));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4380 (.I0(x1683), .I1(x1684), .I2(x1685), .I3(n4374), .I4(n4375), .O(n4380));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4381 (.I0(x1689), .I1(x1690), .I2(x1691), .I3(n4379), .I4(n4380), .O(n4381));
  LUT3 #(.INIT(8'hE8)) lut_n4382 (.I0(x1698), .I1(x1699), .I2(x1700), .O(n4382));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4383 (.I0(x1689), .I1(x1690), .I2(x1691), .I3(n4379), .I4(n4380), .O(n4383));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4384 (.I0(x1695), .I1(x1696), .I2(x1697), .I3(n4382), .I4(n4383), .O(n4384));
  LUT3 #(.INIT(8'h96)) lut_n4385 (.I0(n4373), .I1(n4376), .I2(n4377), .O(n4385));
  LUT3 #(.INIT(8'hE8)) lut_n4386 (.I0(n4381), .I1(n4384), .I2(n4385), .O(n4386));
  LUT3 #(.INIT(8'h96)) lut_n4387 (.I0(n4358), .I1(n4366), .I2(n4367), .O(n4387));
  LUT3 #(.INIT(8'hE8)) lut_n4388 (.I0(n4378), .I1(n4386), .I2(n4387), .O(n4388));
  LUT3 #(.INIT(8'hE8)) lut_n4389 (.I0(x1704), .I1(x1705), .I2(x1706), .O(n4389));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4390 (.I0(x1695), .I1(x1696), .I2(x1697), .I3(n4382), .I4(n4383), .O(n4390));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4391 (.I0(x1701), .I1(x1702), .I2(x1703), .I3(n4389), .I4(n4390), .O(n4391));
  LUT3 #(.INIT(8'hE8)) lut_n4392 (.I0(x1710), .I1(x1711), .I2(x1712), .O(n4392));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4393 (.I0(x1701), .I1(x1702), .I2(x1703), .I3(n4389), .I4(n4390), .O(n4393));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4394 (.I0(x1707), .I1(x1708), .I2(x1709), .I3(n4392), .I4(n4393), .O(n4394));
  LUT3 #(.INIT(8'h96)) lut_n4395 (.I0(n4381), .I1(n4384), .I2(n4385), .O(n4395));
  LUT3 #(.INIT(8'hE8)) lut_n4396 (.I0(n4391), .I1(n4394), .I2(n4395), .O(n4396));
  LUT3 #(.INIT(8'hE8)) lut_n4397 (.I0(x1716), .I1(x1717), .I2(x1718), .O(n4397));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4398 (.I0(x1707), .I1(x1708), .I2(x1709), .I3(n4392), .I4(n4393), .O(n4398));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4399 (.I0(x1713), .I1(x1714), .I2(x1715), .I3(n4397), .I4(n4398), .O(n4399));
  LUT3 #(.INIT(8'hE8)) lut_n4400 (.I0(x1722), .I1(x1723), .I2(x1724), .O(n4400));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4401 (.I0(x1713), .I1(x1714), .I2(x1715), .I3(n4397), .I4(n4398), .O(n4401));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4402 (.I0(x1719), .I1(x1720), .I2(x1721), .I3(n4400), .I4(n4401), .O(n4402));
  LUT3 #(.INIT(8'h96)) lut_n4403 (.I0(n4391), .I1(n4394), .I2(n4395), .O(n4403));
  LUT3 #(.INIT(8'hE8)) lut_n4404 (.I0(n4399), .I1(n4402), .I2(n4403), .O(n4404));
  LUT3 #(.INIT(8'h96)) lut_n4405 (.I0(n4378), .I1(n4386), .I2(n4387), .O(n4405));
  LUT3 #(.INIT(8'hE8)) lut_n4406 (.I0(n4396), .I1(n4404), .I2(n4405), .O(n4406));
  LUT3 #(.INIT(8'h96)) lut_n4407 (.I0(n4350), .I1(n4368), .I2(n4369), .O(n4407));
  LUT3 #(.INIT(8'hE8)) lut_n4408 (.I0(n4388), .I1(n4406), .I2(n4407), .O(n4408));
  LUT3 #(.INIT(8'h96)) lut_n4409 (.I0(n4292), .I1(n4330), .I2(n4331), .O(n4409));
  LUT3 #(.INIT(8'hE8)) lut_n4410 (.I0(n4370), .I1(n4408), .I2(n4409), .O(n4410));
  LUT3 #(.INIT(8'h96)) lut_n4411 (.I0(n4171), .I1(n4249), .I2(n4250), .O(n4411));
  LUT3 #(.INIT(8'hE8)) lut_n4412 (.I0(n4332), .I1(n4410), .I2(n4411), .O(n4412));
  LUT3 #(.INIT(8'hE8)) lut_n4413 (.I0(x1728), .I1(x1729), .I2(x1730), .O(n4413));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4414 (.I0(x1719), .I1(x1720), .I2(x1721), .I3(n4400), .I4(n4401), .O(n4414));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4415 (.I0(x1725), .I1(x1726), .I2(x1727), .I3(n4413), .I4(n4414), .O(n4415));
  LUT3 #(.INIT(8'hE8)) lut_n4416 (.I0(x1734), .I1(x1735), .I2(x1736), .O(n4416));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4417 (.I0(x1725), .I1(x1726), .I2(x1727), .I3(n4413), .I4(n4414), .O(n4417));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4418 (.I0(x1731), .I1(x1732), .I2(x1733), .I3(n4416), .I4(n4417), .O(n4418));
  LUT3 #(.INIT(8'h96)) lut_n4419 (.I0(n4399), .I1(n4402), .I2(n4403), .O(n4419));
  LUT3 #(.INIT(8'hE8)) lut_n4420 (.I0(n4415), .I1(n4418), .I2(n4419), .O(n4420));
  LUT3 #(.INIT(8'hE8)) lut_n4421 (.I0(x1740), .I1(x1741), .I2(x1742), .O(n4421));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4422 (.I0(x1731), .I1(x1732), .I2(x1733), .I3(n4416), .I4(n4417), .O(n4422));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4423 (.I0(x1737), .I1(x1738), .I2(x1739), .I3(n4421), .I4(n4422), .O(n4423));
  LUT3 #(.INIT(8'hE8)) lut_n4424 (.I0(x1746), .I1(x1747), .I2(x1748), .O(n4424));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4425 (.I0(x1737), .I1(x1738), .I2(x1739), .I3(n4421), .I4(n4422), .O(n4425));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4426 (.I0(x1743), .I1(x1744), .I2(x1745), .I3(n4424), .I4(n4425), .O(n4426));
  LUT3 #(.INIT(8'h96)) lut_n4427 (.I0(n4415), .I1(n4418), .I2(n4419), .O(n4427));
  LUT3 #(.INIT(8'hE8)) lut_n4428 (.I0(n4423), .I1(n4426), .I2(n4427), .O(n4428));
  LUT3 #(.INIT(8'h96)) lut_n4429 (.I0(n4396), .I1(n4404), .I2(n4405), .O(n4429));
  LUT3 #(.INIT(8'hE8)) lut_n4430 (.I0(n4420), .I1(n4428), .I2(n4429), .O(n4430));
  LUT3 #(.INIT(8'hE8)) lut_n4431 (.I0(x1752), .I1(x1753), .I2(x1754), .O(n4431));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4432 (.I0(x1743), .I1(x1744), .I2(x1745), .I3(n4424), .I4(n4425), .O(n4432));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4433 (.I0(x1749), .I1(x1750), .I2(x1751), .I3(n4431), .I4(n4432), .O(n4433));
  LUT3 #(.INIT(8'hE8)) lut_n4434 (.I0(x1758), .I1(x1759), .I2(x1760), .O(n4434));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4435 (.I0(x1749), .I1(x1750), .I2(x1751), .I3(n4431), .I4(n4432), .O(n4435));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4436 (.I0(x1755), .I1(x1756), .I2(x1757), .I3(n4434), .I4(n4435), .O(n4436));
  LUT3 #(.INIT(8'h96)) lut_n4437 (.I0(n4423), .I1(n4426), .I2(n4427), .O(n4437));
  LUT3 #(.INIT(8'hE8)) lut_n4438 (.I0(n4433), .I1(n4436), .I2(n4437), .O(n4438));
  LUT3 #(.INIT(8'hE8)) lut_n4439 (.I0(x1764), .I1(x1765), .I2(x1766), .O(n4439));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4440 (.I0(x1755), .I1(x1756), .I2(x1757), .I3(n4434), .I4(n4435), .O(n4440));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4441 (.I0(x1761), .I1(x1762), .I2(x1763), .I3(n4439), .I4(n4440), .O(n4441));
  LUT3 #(.INIT(8'hE8)) lut_n4442 (.I0(x1770), .I1(x1771), .I2(x1772), .O(n4442));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4443 (.I0(x1761), .I1(x1762), .I2(x1763), .I3(n4439), .I4(n4440), .O(n4443));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4444 (.I0(x1767), .I1(x1768), .I2(x1769), .I3(n4442), .I4(n4443), .O(n4444));
  LUT3 #(.INIT(8'h96)) lut_n4445 (.I0(n4433), .I1(n4436), .I2(n4437), .O(n4445));
  LUT3 #(.INIT(8'hE8)) lut_n4446 (.I0(n4441), .I1(n4444), .I2(n4445), .O(n4446));
  LUT3 #(.INIT(8'h96)) lut_n4447 (.I0(n4420), .I1(n4428), .I2(n4429), .O(n4447));
  LUT3 #(.INIT(8'hE8)) lut_n4448 (.I0(n4438), .I1(n4446), .I2(n4447), .O(n4448));
  LUT3 #(.INIT(8'h96)) lut_n4449 (.I0(n4388), .I1(n4406), .I2(n4407), .O(n4449));
  LUT3 #(.INIT(8'hE8)) lut_n4450 (.I0(n4430), .I1(n4448), .I2(n4449), .O(n4450));
  LUT3 #(.INIT(8'hE8)) lut_n4451 (.I0(x1776), .I1(x1777), .I2(x1778), .O(n4451));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4452 (.I0(x1767), .I1(x1768), .I2(x1769), .I3(n4442), .I4(n4443), .O(n4452));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4453 (.I0(x1773), .I1(x1774), .I2(x1775), .I3(n4451), .I4(n4452), .O(n4453));
  LUT3 #(.INIT(8'hE8)) lut_n4454 (.I0(x1782), .I1(x1783), .I2(x1784), .O(n4454));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4455 (.I0(x1773), .I1(x1774), .I2(x1775), .I3(n4451), .I4(n4452), .O(n4455));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4456 (.I0(x1779), .I1(x1780), .I2(x1781), .I3(n4454), .I4(n4455), .O(n4456));
  LUT3 #(.INIT(8'h96)) lut_n4457 (.I0(n4441), .I1(n4444), .I2(n4445), .O(n4457));
  LUT3 #(.INIT(8'hE8)) lut_n4458 (.I0(n4453), .I1(n4456), .I2(n4457), .O(n4458));
  LUT3 #(.INIT(8'hE8)) lut_n4459 (.I0(x1788), .I1(x1789), .I2(x1790), .O(n4459));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4460 (.I0(x1779), .I1(x1780), .I2(x1781), .I3(n4454), .I4(n4455), .O(n4460));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4461 (.I0(x1785), .I1(x1786), .I2(x1787), .I3(n4459), .I4(n4460), .O(n4461));
  LUT3 #(.INIT(8'hE8)) lut_n4462 (.I0(x1794), .I1(x1795), .I2(x1796), .O(n4462));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4463 (.I0(x1785), .I1(x1786), .I2(x1787), .I3(n4459), .I4(n4460), .O(n4463));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4464 (.I0(x1791), .I1(x1792), .I2(x1793), .I3(n4462), .I4(n4463), .O(n4464));
  LUT3 #(.INIT(8'h96)) lut_n4465 (.I0(n4453), .I1(n4456), .I2(n4457), .O(n4465));
  LUT3 #(.INIT(8'hE8)) lut_n4466 (.I0(n4461), .I1(n4464), .I2(n4465), .O(n4466));
  LUT3 #(.INIT(8'h96)) lut_n4467 (.I0(n4438), .I1(n4446), .I2(n4447), .O(n4467));
  LUT3 #(.INIT(8'hE8)) lut_n4468 (.I0(n4458), .I1(n4466), .I2(n4467), .O(n4468));
  LUT3 #(.INIT(8'hE8)) lut_n4469 (.I0(x1800), .I1(x1801), .I2(x1802), .O(n4469));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4470 (.I0(x1791), .I1(x1792), .I2(x1793), .I3(n4462), .I4(n4463), .O(n4470));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4471 (.I0(x1797), .I1(x1798), .I2(x1799), .I3(n4469), .I4(n4470), .O(n4471));
  LUT3 #(.INIT(8'hE8)) lut_n4472 (.I0(x1806), .I1(x1807), .I2(x1808), .O(n4472));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4473 (.I0(x1797), .I1(x1798), .I2(x1799), .I3(n4469), .I4(n4470), .O(n4473));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4474 (.I0(x1803), .I1(x1804), .I2(x1805), .I3(n4472), .I4(n4473), .O(n4474));
  LUT3 #(.INIT(8'h96)) lut_n4475 (.I0(n4461), .I1(n4464), .I2(n4465), .O(n4475));
  LUT3 #(.INIT(8'hE8)) lut_n4476 (.I0(n4471), .I1(n4474), .I2(n4475), .O(n4476));
  LUT3 #(.INIT(8'hE8)) lut_n4477 (.I0(x1812), .I1(x1813), .I2(x1814), .O(n4477));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4478 (.I0(x1803), .I1(x1804), .I2(x1805), .I3(n4472), .I4(n4473), .O(n4478));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4479 (.I0(x1809), .I1(x1810), .I2(x1811), .I3(n4477), .I4(n4478), .O(n4479));
  LUT3 #(.INIT(8'hE8)) lut_n4480 (.I0(x1818), .I1(x1819), .I2(x1820), .O(n4480));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4481 (.I0(x1809), .I1(x1810), .I2(x1811), .I3(n4477), .I4(n4478), .O(n4481));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4482 (.I0(x1815), .I1(x1816), .I2(x1817), .I3(n4480), .I4(n4481), .O(n4482));
  LUT3 #(.INIT(8'h96)) lut_n4483 (.I0(n4471), .I1(n4474), .I2(n4475), .O(n4483));
  LUT3 #(.INIT(8'hE8)) lut_n4484 (.I0(n4479), .I1(n4482), .I2(n4483), .O(n4484));
  LUT3 #(.INIT(8'h96)) lut_n4485 (.I0(n4458), .I1(n4466), .I2(n4467), .O(n4485));
  LUT3 #(.INIT(8'hE8)) lut_n4486 (.I0(n4476), .I1(n4484), .I2(n4485), .O(n4486));
  LUT3 #(.INIT(8'h96)) lut_n4487 (.I0(n4430), .I1(n4448), .I2(n4449), .O(n4487));
  LUT3 #(.INIT(8'hE8)) lut_n4488 (.I0(n4468), .I1(n4486), .I2(n4487), .O(n4488));
  LUT3 #(.INIT(8'h96)) lut_n4489 (.I0(n4370), .I1(n4408), .I2(n4409), .O(n4489));
  LUT3 #(.INIT(8'hE8)) lut_n4490 (.I0(n4450), .I1(n4488), .I2(n4489), .O(n4490));
  LUT3 #(.INIT(8'hE8)) lut_n4491 (.I0(x1824), .I1(x1825), .I2(x1826), .O(n4491));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4492 (.I0(x1815), .I1(x1816), .I2(x1817), .I3(n4480), .I4(n4481), .O(n4492));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4493 (.I0(x1821), .I1(x1822), .I2(x1823), .I3(n4491), .I4(n4492), .O(n4493));
  LUT3 #(.INIT(8'hE8)) lut_n4494 (.I0(x1830), .I1(x1831), .I2(x1832), .O(n4494));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4495 (.I0(x1821), .I1(x1822), .I2(x1823), .I3(n4491), .I4(n4492), .O(n4495));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4496 (.I0(x1827), .I1(x1828), .I2(x1829), .I3(n4494), .I4(n4495), .O(n4496));
  LUT3 #(.INIT(8'h96)) lut_n4497 (.I0(n4479), .I1(n4482), .I2(n4483), .O(n4497));
  LUT3 #(.INIT(8'hE8)) lut_n4498 (.I0(n4493), .I1(n4496), .I2(n4497), .O(n4498));
  LUT3 #(.INIT(8'hE8)) lut_n4499 (.I0(x1836), .I1(x1837), .I2(x1838), .O(n4499));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4500 (.I0(x1827), .I1(x1828), .I2(x1829), .I3(n4494), .I4(n4495), .O(n4500));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4501 (.I0(x1833), .I1(x1834), .I2(x1835), .I3(n4499), .I4(n4500), .O(n4501));
  LUT3 #(.INIT(8'hE8)) lut_n4502 (.I0(x1842), .I1(x1843), .I2(x1844), .O(n4502));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4503 (.I0(x1833), .I1(x1834), .I2(x1835), .I3(n4499), .I4(n4500), .O(n4503));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4504 (.I0(x1839), .I1(x1840), .I2(x1841), .I3(n4502), .I4(n4503), .O(n4504));
  LUT3 #(.INIT(8'h96)) lut_n4505 (.I0(n4493), .I1(n4496), .I2(n4497), .O(n4505));
  LUT3 #(.INIT(8'hE8)) lut_n4506 (.I0(n4501), .I1(n4504), .I2(n4505), .O(n4506));
  LUT3 #(.INIT(8'h96)) lut_n4507 (.I0(n4476), .I1(n4484), .I2(n4485), .O(n4507));
  LUT3 #(.INIT(8'hE8)) lut_n4508 (.I0(n4498), .I1(n4506), .I2(n4507), .O(n4508));
  LUT3 #(.INIT(8'hE8)) lut_n4509 (.I0(x1848), .I1(x1849), .I2(x1850), .O(n4509));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4510 (.I0(x1839), .I1(x1840), .I2(x1841), .I3(n4502), .I4(n4503), .O(n4510));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4511 (.I0(x1845), .I1(x1846), .I2(x1847), .I3(n4509), .I4(n4510), .O(n4511));
  LUT3 #(.INIT(8'hE8)) lut_n4512 (.I0(x1854), .I1(x1855), .I2(x1856), .O(n4512));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4513 (.I0(x1845), .I1(x1846), .I2(x1847), .I3(n4509), .I4(n4510), .O(n4513));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4514 (.I0(x1851), .I1(x1852), .I2(x1853), .I3(n4512), .I4(n4513), .O(n4514));
  LUT3 #(.INIT(8'h96)) lut_n4515 (.I0(n4501), .I1(n4504), .I2(n4505), .O(n4515));
  LUT3 #(.INIT(8'hE8)) lut_n4516 (.I0(n4511), .I1(n4514), .I2(n4515), .O(n4516));
  LUT3 #(.INIT(8'hE8)) lut_n4517 (.I0(x1860), .I1(x1861), .I2(x1862), .O(n4517));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4518 (.I0(x1851), .I1(x1852), .I2(x1853), .I3(n4512), .I4(n4513), .O(n4518));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4519 (.I0(x1857), .I1(x1858), .I2(x1859), .I3(n4517), .I4(n4518), .O(n4519));
  LUT3 #(.INIT(8'hE8)) lut_n4520 (.I0(x1866), .I1(x1867), .I2(x1868), .O(n4520));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4521 (.I0(x1857), .I1(x1858), .I2(x1859), .I3(n4517), .I4(n4518), .O(n4521));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4522 (.I0(x1863), .I1(x1864), .I2(x1865), .I3(n4520), .I4(n4521), .O(n4522));
  LUT3 #(.INIT(8'h96)) lut_n4523 (.I0(n4511), .I1(n4514), .I2(n4515), .O(n4523));
  LUT3 #(.INIT(8'hE8)) lut_n4524 (.I0(n4519), .I1(n4522), .I2(n4523), .O(n4524));
  LUT3 #(.INIT(8'h96)) lut_n4525 (.I0(n4498), .I1(n4506), .I2(n4507), .O(n4525));
  LUT3 #(.INIT(8'hE8)) lut_n4526 (.I0(n4516), .I1(n4524), .I2(n4525), .O(n4526));
  LUT3 #(.INIT(8'h96)) lut_n4527 (.I0(n4468), .I1(n4486), .I2(n4487), .O(n4527));
  LUT3 #(.INIT(8'hE8)) lut_n4528 (.I0(n4508), .I1(n4526), .I2(n4527), .O(n4528));
  LUT3 #(.INIT(8'hE8)) lut_n4529 (.I0(x1872), .I1(x1873), .I2(x1874), .O(n4529));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4530 (.I0(x1863), .I1(x1864), .I2(x1865), .I3(n4520), .I4(n4521), .O(n4530));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4531 (.I0(x1869), .I1(x1870), .I2(x1871), .I3(n4529), .I4(n4530), .O(n4531));
  LUT3 #(.INIT(8'hE8)) lut_n4532 (.I0(x1878), .I1(x1879), .I2(x1880), .O(n4532));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4533 (.I0(x1869), .I1(x1870), .I2(x1871), .I3(n4529), .I4(n4530), .O(n4533));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4534 (.I0(x1875), .I1(x1876), .I2(x1877), .I3(n4532), .I4(n4533), .O(n4534));
  LUT3 #(.INIT(8'h96)) lut_n4535 (.I0(n4519), .I1(n4522), .I2(n4523), .O(n4535));
  LUT3 #(.INIT(8'hE8)) lut_n4536 (.I0(n4531), .I1(n4534), .I2(n4535), .O(n4536));
  LUT3 #(.INIT(8'hE8)) lut_n4537 (.I0(x1884), .I1(x1885), .I2(x1886), .O(n4537));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4538 (.I0(x1875), .I1(x1876), .I2(x1877), .I3(n4532), .I4(n4533), .O(n4538));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4539 (.I0(x1881), .I1(x1882), .I2(x1883), .I3(n4537), .I4(n4538), .O(n4539));
  LUT3 #(.INIT(8'hE8)) lut_n4540 (.I0(x1890), .I1(x1891), .I2(x1892), .O(n4540));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4541 (.I0(x1881), .I1(x1882), .I2(x1883), .I3(n4537), .I4(n4538), .O(n4541));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4542 (.I0(x1887), .I1(x1888), .I2(x1889), .I3(n4540), .I4(n4541), .O(n4542));
  LUT3 #(.INIT(8'h96)) lut_n4543 (.I0(n4531), .I1(n4534), .I2(n4535), .O(n4543));
  LUT3 #(.INIT(8'hE8)) lut_n4544 (.I0(n4539), .I1(n4542), .I2(n4543), .O(n4544));
  LUT3 #(.INIT(8'h96)) lut_n4545 (.I0(n4516), .I1(n4524), .I2(n4525), .O(n4545));
  LUT3 #(.INIT(8'hE8)) lut_n4546 (.I0(n4536), .I1(n4544), .I2(n4545), .O(n4546));
  LUT3 #(.INIT(8'hE8)) lut_n4547 (.I0(x1896), .I1(x1897), .I2(x1898), .O(n4547));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4548 (.I0(x1887), .I1(x1888), .I2(x1889), .I3(n4540), .I4(n4541), .O(n4548));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4549 (.I0(x1893), .I1(x1894), .I2(x1895), .I3(n4547), .I4(n4548), .O(n4549));
  LUT3 #(.INIT(8'hE8)) lut_n4550 (.I0(x1902), .I1(x1903), .I2(x1904), .O(n4550));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4551 (.I0(x1893), .I1(x1894), .I2(x1895), .I3(n4547), .I4(n4548), .O(n4551));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4552 (.I0(x1899), .I1(x1900), .I2(x1901), .I3(n4550), .I4(n4551), .O(n4552));
  LUT3 #(.INIT(8'h96)) lut_n4553 (.I0(n4539), .I1(n4542), .I2(n4543), .O(n4553));
  LUT3 #(.INIT(8'hE8)) lut_n4554 (.I0(n4549), .I1(n4552), .I2(n4553), .O(n4554));
  LUT3 #(.INIT(8'hE8)) lut_n4555 (.I0(x1908), .I1(x1909), .I2(x1910), .O(n4555));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4556 (.I0(x1899), .I1(x1900), .I2(x1901), .I3(n4550), .I4(n4551), .O(n4556));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4557 (.I0(x1905), .I1(x1906), .I2(x1907), .I3(n4555), .I4(n4556), .O(n4557));
  LUT3 #(.INIT(8'hE8)) lut_n4558 (.I0(x1914), .I1(x1915), .I2(x1916), .O(n4558));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4559 (.I0(x1905), .I1(x1906), .I2(x1907), .I3(n4555), .I4(n4556), .O(n4559));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4560 (.I0(x1911), .I1(x1912), .I2(x1913), .I3(n4558), .I4(n4559), .O(n4560));
  LUT3 #(.INIT(8'h96)) lut_n4561 (.I0(n4549), .I1(n4552), .I2(n4553), .O(n4561));
  LUT3 #(.INIT(8'hE8)) lut_n4562 (.I0(n4557), .I1(n4560), .I2(n4561), .O(n4562));
  LUT3 #(.INIT(8'h96)) lut_n4563 (.I0(n4536), .I1(n4544), .I2(n4545), .O(n4563));
  LUT3 #(.INIT(8'hE8)) lut_n4564 (.I0(n4554), .I1(n4562), .I2(n4563), .O(n4564));
  LUT3 #(.INIT(8'h96)) lut_n4565 (.I0(n4508), .I1(n4526), .I2(n4527), .O(n4565));
  LUT3 #(.INIT(8'hE8)) lut_n4566 (.I0(n4546), .I1(n4564), .I2(n4565), .O(n4566));
  LUT3 #(.INIT(8'h96)) lut_n4567 (.I0(n4450), .I1(n4488), .I2(n4489), .O(n4567));
  LUT3 #(.INIT(8'hE8)) lut_n4568 (.I0(n4528), .I1(n4566), .I2(n4567), .O(n4568));
  LUT3 #(.INIT(8'h96)) lut_n4569 (.I0(n4332), .I1(n4410), .I2(n4411), .O(n4569));
  LUT3 #(.INIT(8'hE8)) lut_n4570 (.I0(n4490), .I1(n4568), .I2(n4569), .O(n4570));
  LUT3 #(.INIT(8'h96)) lut_n4571 (.I0(n4093), .I1(n4251), .I2(n4252), .O(n4571));
  LUT3 #(.INIT(8'hE8)) lut_n4572 (.I0(n4412), .I1(n4570), .I2(n4571), .O(n4572));
  LUT3 #(.INIT(8'hE8)) lut_n4573 (.I0(x1920), .I1(x1921), .I2(x1922), .O(n4573));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4574 (.I0(x1911), .I1(x1912), .I2(x1913), .I3(n4558), .I4(n4559), .O(n4574));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4575 (.I0(x1917), .I1(x1918), .I2(x1919), .I3(n4573), .I4(n4574), .O(n4575));
  LUT3 #(.INIT(8'hE8)) lut_n4576 (.I0(x1926), .I1(x1927), .I2(x1928), .O(n4576));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4577 (.I0(x1917), .I1(x1918), .I2(x1919), .I3(n4573), .I4(n4574), .O(n4577));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4578 (.I0(x1923), .I1(x1924), .I2(x1925), .I3(n4576), .I4(n4577), .O(n4578));
  LUT3 #(.INIT(8'h96)) lut_n4579 (.I0(n4557), .I1(n4560), .I2(n4561), .O(n4579));
  LUT3 #(.INIT(8'hE8)) lut_n4580 (.I0(n4575), .I1(n4578), .I2(n4579), .O(n4580));
  LUT3 #(.INIT(8'hE8)) lut_n4581 (.I0(x1932), .I1(x1933), .I2(x1934), .O(n4581));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4582 (.I0(x1923), .I1(x1924), .I2(x1925), .I3(n4576), .I4(n4577), .O(n4582));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4583 (.I0(x1929), .I1(x1930), .I2(x1931), .I3(n4581), .I4(n4582), .O(n4583));
  LUT3 #(.INIT(8'hE8)) lut_n4584 (.I0(x1938), .I1(x1939), .I2(x1940), .O(n4584));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4585 (.I0(x1929), .I1(x1930), .I2(x1931), .I3(n4581), .I4(n4582), .O(n4585));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4586 (.I0(x1935), .I1(x1936), .I2(x1937), .I3(n4584), .I4(n4585), .O(n4586));
  LUT3 #(.INIT(8'h96)) lut_n4587 (.I0(n4575), .I1(n4578), .I2(n4579), .O(n4587));
  LUT3 #(.INIT(8'hE8)) lut_n4588 (.I0(n4583), .I1(n4586), .I2(n4587), .O(n4588));
  LUT3 #(.INIT(8'h96)) lut_n4589 (.I0(n4554), .I1(n4562), .I2(n4563), .O(n4589));
  LUT3 #(.INIT(8'hE8)) lut_n4590 (.I0(n4580), .I1(n4588), .I2(n4589), .O(n4590));
  LUT3 #(.INIT(8'hE8)) lut_n4591 (.I0(x1944), .I1(x1945), .I2(x1946), .O(n4591));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4592 (.I0(x1935), .I1(x1936), .I2(x1937), .I3(n4584), .I4(n4585), .O(n4592));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4593 (.I0(x1941), .I1(x1942), .I2(x1943), .I3(n4591), .I4(n4592), .O(n4593));
  LUT3 #(.INIT(8'hE8)) lut_n4594 (.I0(x1950), .I1(x1951), .I2(x1952), .O(n4594));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4595 (.I0(x1941), .I1(x1942), .I2(x1943), .I3(n4591), .I4(n4592), .O(n4595));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4596 (.I0(x1947), .I1(x1948), .I2(x1949), .I3(n4594), .I4(n4595), .O(n4596));
  LUT3 #(.INIT(8'h96)) lut_n4597 (.I0(n4583), .I1(n4586), .I2(n4587), .O(n4597));
  LUT3 #(.INIT(8'hE8)) lut_n4598 (.I0(n4593), .I1(n4596), .I2(n4597), .O(n4598));
  LUT3 #(.INIT(8'hE8)) lut_n4599 (.I0(x1956), .I1(x1957), .I2(x1958), .O(n4599));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4600 (.I0(x1947), .I1(x1948), .I2(x1949), .I3(n4594), .I4(n4595), .O(n4600));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4601 (.I0(x1953), .I1(x1954), .I2(x1955), .I3(n4599), .I4(n4600), .O(n4601));
  LUT3 #(.INIT(8'hE8)) lut_n4602 (.I0(x1962), .I1(x1963), .I2(x1964), .O(n4602));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4603 (.I0(x1953), .I1(x1954), .I2(x1955), .I3(n4599), .I4(n4600), .O(n4603));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4604 (.I0(x1959), .I1(x1960), .I2(x1961), .I3(n4602), .I4(n4603), .O(n4604));
  LUT3 #(.INIT(8'h96)) lut_n4605 (.I0(n4593), .I1(n4596), .I2(n4597), .O(n4605));
  LUT3 #(.INIT(8'hE8)) lut_n4606 (.I0(n4601), .I1(n4604), .I2(n4605), .O(n4606));
  LUT3 #(.INIT(8'h96)) lut_n4607 (.I0(n4580), .I1(n4588), .I2(n4589), .O(n4607));
  LUT3 #(.INIT(8'hE8)) lut_n4608 (.I0(n4598), .I1(n4606), .I2(n4607), .O(n4608));
  LUT3 #(.INIT(8'h96)) lut_n4609 (.I0(n4546), .I1(n4564), .I2(n4565), .O(n4609));
  LUT3 #(.INIT(8'hE8)) lut_n4610 (.I0(n4590), .I1(n4608), .I2(n4609), .O(n4610));
  LUT3 #(.INIT(8'hE8)) lut_n4611 (.I0(x1968), .I1(x1969), .I2(x1970), .O(n4611));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4612 (.I0(x1959), .I1(x1960), .I2(x1961), .I3(n4602), .I4(n4603), .O(n4612));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4613 (.I0(x1965), .I1(x1966), .I2(x1967), .I3(n4611), .I4(n4612), .O(n4613));
  LUT3 #(.INIT(8'hE8)) lut_n4614 (.I0(x1974), .I1(x1975), .I2(x1976), .O(n4614));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4615 (.I0(x1965), .I1(x1966), .I2(x1967), .I3(n4611), .I4(n4612), .O(n4615));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4616 (.I0(x1971), .I1(x1972), .I2(x1973), .I3(n4614), .I4(n4615), .O(n4616));
  LUT3 #(.INIT(8'h96)) lut_n4617 (.I0(n4601), .I1(n4604), .I2(n4605), .O(n4617));
  LUT3 #(.INIT(8'hE8)) lut_n4618 (.I0(n4613), .I1(n4616), .I2(n4617), .O(n4618));
  LUT3 #(.INIT(8'hE8)) lut_n4619 (.I0(x1980), .I1(x1981), .I2(x1982), .O(n4619));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4620 (.I0(x1971), .I1(x1972), .I2(x1973), .I3(n4614), .I4(n4615), .O(n4620));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4621 (.I0(x1977), .I1(x1978), .I2(x1979), .I3(n4619), .I4(n4620), .O(n4621));
  LUT3 #(.INIT(8'hE8)) lut_n4622 (.I0(x1986), .I1(x1987), .I2(x1988), .O(n4622));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4623 (.I0(x1977), .I1(x1978), .I2(x1979), .I3(n4619), .I4(n4620), .O(n4623));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4624 (.I0(x1983), .I1(x1984), .I2(x1985), .I3(n4622), .I4(n4623), .O(n4624));
  LUT3 #(.INIT(8'h96)) lut_n4625 (.I0(n4613), .I1(n4616), .I2(n4617), .O(n4625));
  LUT3 #(.INIT(8'hE8)) lut_n4626 (.I0(n4621), .I1(n4624), .I2(n4625), .O(n4626));
  LUT3 #(.INIT(8'h96)) lut_n4627 (.I0(n4598), .I1(n4606), .I2(n4607), .O(n4627));
  LUT3 #(.INIT(8'hE8)) lut_n4628 (.I0(n4618), .I1(n4626), .I2(n4627), .O(n4628));
  LUT3 #(.INIT(8'hE8)) lut_n4629 (.I0(x1992), .I1(x1993), .I2(x1994), .O(n4629));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4630 (.I0(x1983), .I1(x1984), .I2(x1985), .I3(n4622), .I4(n4623), .O(n4630));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4631 (.I0(x1989), .I1(x1990), .I2(x1991), .I3(n4629), .I4(n4630), .O(n4631));
  LUT3 #(.INIT(8'hE8)) lut_n4632 (.I0(x1998), .I1(x1999), .I2(x2000), .O(n4632));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4633 (.I0(x1989), .I1(x1990), .I2(x1991), .I3(n4629), .I4(n4630), .O(n4633));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4634 (.I0(x1995), .I1(x1996), .I2(x1997), .I3(n4632), .I4(n4633), .O(n4634));
  LUT3 #(.INIT(8'h96)) lut_n4635 (.I0(n4621), .I1(n4624), .I2(n4625), .O(n4635));
  LUT3 #(.INIT(8'hE8)) lut_n4636 (.I0(n4631), .I1(n4634), .I2(n4635), .O(n4636));
  LUT3 #(.INIT(8'hE8)) lut_n4637 (.I0(x2004), .I1(x2005), .I2(x2006), .O(n4637));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4638 (.I0(x1995), .I1(x1996), .I2(x1997), .I3(n4632), .I4(n4633), .O(n4638));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4639 (.I0(x2001), .I1(x2002), .I2(x2003), .I3(n4637), .I4(n4638), .O(n4639));
  LUT3 #(.INIT(8'hE8)) lut_n4640 (.I0(x2010), .I1(x2011), .I2(x2012), .O(n4640));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4641 (.I0(x2001), .I1(x2002), .I2(x2003), .I3(n4637), .I4(n4638), .O(n4641));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4642 (.I0(x2007), .I1(x2008), .I2(x2009), .I3(n4640), .I4(n4641), .O(n4642));
  LUT3 #(.INIT(8'h96)) lut_n4643 (.I0(n4631), .I1(n4634), .I2(n4635), .O(n4643));
  LUT3 #(.INIT(8'hE8)) lut_n4644 (.I0(n4639), .I1(n4642), .I2(n4643), .O(n4644));
  LUT3 #(.INIT(8'h96)) lut_n4645 (.I0(n4618), .I1(n4626), .I2(n4627), .O(n4645));
  LUT3 #(.INIT(8'hE8)) lut_n4646 (.I0(n4636), .I1(n4644), .I2(n4645), .O(n4646));
  LUT3 #(.INIT(8'h96)) lut_n4647 (.I0(n4590), .I1(n4608), .I2(n4609), .O(n4647));
  LUT3 #(.INIT(8'hE8)) lut_n4648 (.I0(n4628), .I1(n4646), .I2(n4647), .O(n4648));
  LUT3 #(.INIT(8'h96)) lut_n4649 (.I0(n4528), .I1(n4566), .I2(n4567), .O(n4649));
  LUT3 #(.INIT(8'hE8)) lut_n4650 (.I0(n4610), .I1(n4648), .I2(n4649), .O(n4650));
  LUT3 #(.INIT(8'hE8)) lut_n4651 (.I0(x2016), .I1(x2017), .I2(x2018), .O(n4651));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4652 (.I0(x2007), .I1(x2008), .I2(x2009), .I3(n4640), .I4(n4641), .O(n4652));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4653 (.I0(x2013), .I1(x2014), .I2(x2015), .I3(n4651), .I4(n4652), .O(n4653));
  LUT3 #(.INIT(8'hE8)) lut_n4654 (.I0(x2022), .I1(x2023), .I2(x2024), .O(n4654));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4655 (.I0(x2013), .I1(x2014), .I2(x2015), .I3(n4651), .I4(n4652), .O(n4655));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4656 (.I0(x2019), .I1(x2020), .I2(x2021), .I3(n4654), .I4(n4655), .O(n4656));
  LUT3 #(.INIT(8'h96)) lut_n4657 (.I0(n4639), .I1(n4642), .I2(n4643), .O(n4657));
  LUT3 #(.INIT(8'hE8)) lut_n4658 (.I0(n4653), .I1(n4656), .I2(n4657), .O(n4658));
  LUT3 #(.INIT(8'hE8)) lut_n4659 (.I0(x2028), .I1(x2029), .I2(x2030), .O(n4659));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4660 (.I0(x2019), .I1(x2020), .I2(x2021), .I3(n4654), .I4(n4655), .O(n4660));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4661 (.I0(x2025), .I1(x2026), .I2(x2027), .I3(n4659), .I4(n4660), .O(n4661));
  LUT3 #(.INIT(8'hE8)) lut_n4662 (.I0(x2034), .I1(x2035), .I2(x2036), .O(n4662));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4663 (.I0(x2025), .I1(x2026), .I2(x2027), .I3(n4659), .I4(n4660), .O(n4663));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4664 (.I0(x2031), .I1(x2032), .I2(x2033), .I3(n4662), .I4(n4663), .O(n4664));
  LUT3 #(.INIT(8'h96)) lut_n4665 (.I0(n4653), .I1(n4656), .I2(n4657), .O(n4665));
  LUT3 #(.INIT(8'hE8)) lut_n4666 (.I0(n4661), .I1(n4664), .I2(n4665), .O(n4666));
  LUT3 #(.INIT(8'h96)) lut_n4667 (.I0(n4636), .I1(n4644), .I2(n4645), .O(n4667));
  LUT3 #(.INIT(8'hE8)) lut_n4668 (.I0(n4658), .I1(n4666), .I2(n4667), .O(n4668));
  LUT3 #(.INIT(8'hE8)) lut_n4669 (.I0(x2040), .I1(x2041), .I2(x2042), .O(n4669));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4670 (.I0(x2031), .I1(x2032), .I2(x2033), .I3(n4662), .I4(n4663), .O(n4670));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4671 (.I0(x2037), .I1(x2038), .I2(x2039), .I3(n4669), .I4(n4670), .O(n4671));
  LUT3 #(.INIT(8'hE8)) lut_n4672 (.I0(x2046), .I1(x2047), .I2(x2048), .O(n4672));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4673 (.I0(x2037), .I1(x2038), .I2(x2039), .I3(n4669), .I4(n4670), .O(n4673));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4674 (.I0(x2043), .I1(x2044), .I2(x2045), .I3(n4672), .I4(n4673), .O(n4674));
  LUT3 #(.INIT(8'h96)) lut_n4675 (.I0(n4661), .I1(n4664), .I2(n4665), .O(n4675));
  LUT3 #(.INIT(8'hE8)) lut_n4676 (.I0(n4671), .I1(n4674), .I2(n4675), .O(n4676));
  LUT3 #(.INIT(8'hE8)) lut_n4677 (.I0(x2052), .I1(x2053), .I2(x2054), .O(n4677));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4678 (.I0(x2043), .I1(x2044), .I2(x2045), .I3(n4672), .I4(n4673), .O(n4678));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4679 (.I0(x2049), .I1(x2050), .I2(x2051), .I3(n4677), .I4(n4678), .O(n4679));
  LUT3 #(.INIT(8'hE8)) lut_n4680 (.I0(x2058), .I1(x2059), .I2(x2060), .O(n4680));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4681 (.I0(x2049), .I1(x2050), .I2(x2051), .I3(n4677), .I4(n4678), .O(n4681));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4682 (.I0(x2055), .I1(x2056), .I2(x2057), .I3(n4680), .I4(n4681), .O(n4682));
  LUT3 #(.INIT(8'h96)) lut_n4683 (.I0(n4671), .I1(n4674), .I2(n4675), .O(n4683));
  LUT3 #(.INIT(8'hE8)) lut_n4684 (.I0(n4679), .I1(n4682), .I2(n4683), .O(n4684));
  LUT3 #(.INIT(8'h96)) lut_n4685 (.I0(n4658), .I1(n4666), .I2(n4667), .O(n4685));
  LUT3 #(.INIT(8'hE8)) lut_n4686 (.I0(n4676), .I1(n4684), .I2(n4685), .O(n4686));
  LUT3 #(.INIT(8'h96)) lut_n4687 (.I0(n4628), .I1(n4646), .I2(n4647), .O(n4687));
  LUT3 #(.INIT(8'hE8)) lut_n4688 (.I0(n4668), .I1(n4686), .I2(n4687), .O(n4688));
  LUT3 #(.INIT(8'hE8)) lut_n4689 (.I0(x2064), .I1(x2065), .I2(x2066), .O(n4689));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4690 (.I0(x2055), .I1(x2056), .I2(x2057), .I3(n4680), .I4(n4681), .O(n4690));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4691 (.I0(x2061), .I1(x2062), .I2(x2063), .I3(n4689), .I4(n4690), .O(n4691));
  LUT3 #(.INIT(8'hE8)) lut_n4692 (.I0(x2070), .I1(x2071), .I2(x2072), .O(n4692));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4693 (.I0(x2061), .I1(x2062), .I2(x2063), .I3(n4689), .I4(n4690), .O(n4693));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4694 (.I0(x2067), .I1(x2068), .I2(x2069), .I3(n4692), .I4(n4693), .O(n4694));
  LUT3 #(.INIT(8'h96)) lut_n4695 (.I0(n4679), .I1(n4682), .I2(n4683), .O(n4695));
  LUT3 #(.INIT(8'hE8)) lut_n4696 (.I0(n4691), .I1(n4694), .I2(n4695), .O(n4696));
  LUT3 #(.INIT(8'hE8)) lut_n4697 (.I0(x2076), .I1(x2077), .I2(x2078), .O(n4697));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4698 (.I0(x2067), .I1(x2068), .I2(x2069), .I3(n4692), .I4(n4693), .O(n4698));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4699 (.I0(x2073), .I1(x2074), .I2(x2075), .I3(n4697), .I4(n4698), .O(n4699));
  LUT3 #(.INIT(8'hE8)) lut_n4700 (.I0(x2082), .I1(x2083), .I2(x2084), .O(n4700));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4701 (.I0(x2073), .I1(x2074), .I2(x2075), .I3(n4697), .I4(n4698), .O(n4701));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4702 (.I0(x2079), .I1(x2080), .I2(x2081), .I3(n4700), .I4(n4701), .O(n4702));
  LUT3 #(.INIT(8'h96)) lut_n4703 (.I0(n4691), .I1(n4694), .I2(n4695), .O(n4703));
  LUT3 #(.INIT(8'hE8)) lut_n4704 (.I0(n4699), .I1(n4702), .I2(n4703), .O(n4704));
  LUT3 #(.INIT(8'h96)) lut_n4705 (.I0(n4676), .I1(n4684), .I2(n4685), .O(n4705));
  LUT3 #(.INIT(8'hE8)) lut_n4706 (.I0(n4696), .I1(n4704), .I2(n4705), .O(n4706));
  LUT3 #(.INIT(8'hE8)) lut_n4707 (.I0(x2088), .I1(x2089), .I2(x2090), .O(n4707));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4708 (.I0(x2079), .I1(x2080), .I2(x2081), .I3(n4700), .I4(n4701), .O(n4708));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4709 (.I0(x2085), .I1(x2086), .I2(x2087), .I3(n4707), .I4(n4708), .O(n4709));
  LUT3 #(.INIT(8'hE8)) lut_n4710 (.I0(x2094), .I1(x2095), .I2(x2096), .O(n4710));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4711 (.I0(x2085), .I1(x2086), .I2(x2087), .I3(n4707), .I4(n4708), .O(n4711));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4712 (.I0(x2091), .I1(x2092), .I2(x2093), .I3(n4710), .I4(n4711), .O(n4712));
  LUT3 #(.INIT(8'h96)) lut_n4713 (.I0(n4699), .I1(n4702), .I2(n4703), .O(n4713));
  LUT3 #(.INIT(8'hE8)) lut_n4714 (.I0(n4709), .I1(n4712), .I2(n4713), .O(n4714));
  LUT3 #(.INIT(8'hE8)) lut_n4715 (.I0(x2100), .I1(x2101), .I2(x2102), .O(n4715));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4716 (.I0(x2091), .I1(x2092), .I2(x2093), .I3(n4710), .I4(n4711), .O(n4716));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4717 (.I0(x2097), .I1(x2098), .I2(x2099), .I3(n4715), .I4(n4716), .O(n4717));
  LUT3 #(.INIT(8'hE8)) lut_n4718 (.I0(x2106), .I1(x2107), .I2(x2108), .O(n4718));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4719 (.I0(x2097), .I1(x2098), .I2(x2099), .I3(n4715), .I4(n4716), .O(n4719));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4720 (.I0(x2103), .I1(x2104), .I2(x2105), .I3(n4718), .I4(n4719), .O(n4720));
  LUT3 #(.INIT(8'h96)) lut_n4721 (.I0(n4709), .I1(n4712), .I2(n4713), .O(n4721));
  LUT3 #(.INIT(8'hE8)) lut_n4722 (.I0(n4717), .I1(n4720), .I2(n4721), .O(n4722));
  LUT3 #(.INIT(8'h96)) lut_n4723 (.I0(n4696), .I1(n4704), .I2(n4705), .O(n4723));
  LUT3 #(.INIT(8'hE8)) lut_n4724 (.I0(n4714), .I1(n4722), .I2(n4723), .O(n4724));
  LUT3 #(.INIT(8'h96)) lut_n4725 (.I0(n4668), .I1(n4686), .I2(n4687), .O(n4725));
  LUT3 #(.INIT(8'hE8)) lut_n4726 (.I0(n4706), .I1(n4724), .I2(n4725), .O(n4726));
  LUT3 #(.INIT(8'h96)) lut_n4727 (.I0(n4610), .I1(n4648), .I2(n4649), .O(n4727));
  LUT3 #(.INIT(8'hE8)) lut_n4728 (.I0(n4688), .I1(n4726), .I2(n4727), .O(n4728));
  LUT3 #(.INIT(8'h96)) lut_n4729 (.I0(n4490), .I1(n4568), .I2(n4569), .O(n4729));
  LUT3 #(.INIT(8'hE8)) lut_n4730 (.I0(n4650), .I1(n4728), .I2(n4729), .O(n4730));
  LUT3 #(.INIT(8'hE8)) lut_n4731 (.I0(x2112), .I1(x2113), .I2(x2114), .O(n4731));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4732 (.I0(x2103), .I1(x2104), .I2(x2105), .I3(n4718), .I4(n4719), .O(n4732));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4733 (.I0(x2109), .I1(x2110), .I2(x2111), .I3(n4731), .I4(n4732), .O(n4733));
  LUT3 #(.INIT(8'hE8)) lut_n4734 (.I0(x2118), .I1(x2119), .I2(x2120), .O(n4734));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4735 (.I0(x2109), .I1(x2110), .I2(x2111), .I3(n4731), .I4(n4732), .O(n4735));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4736 (.I0(x2115), .I1(x2116), .I2(x2117), .I3(n4734), .I4(n4735), .O(n4736));
  LUT3 #(.INIT(8'h96)) lut_n4737 (.I0(n4717), .I1(n4720), .I2(n4721), .O(n4737));
  LUT3 #(.INIT(8'hE8)) lut_n4738 (.I0(n4733), .I1(n4736), .I2(n4737), .O(n4738));
  LUT3 #(.INIT(8'hE8)) lut_n4739 (.I0(x2124), .I1(x2125), .I2(x2126), .O(n4739));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4740 (.I0(x2115), .I1(x2116), .I2(x2117), .I3(n4734), .I4(n4735), .O(n4740));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4741 (.I0(x2121), .I1(x2122), .I2(x2123), .I3(n4739), .I4(n4740), .O(n4741));
  LUT3 #(.INIT(8'hE8)) lut_n4742 (.I0(x2130), .I1(x2131), .I2(x2132), .O(n4742));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4743 (.I0(x2121), .I1(x2122), .I2(x2123), .I3(n4739), .I4(n4740), .O(n4743));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4744 (.I0(x2127), .I1(x2128), .I2(x2129), .I3(n4742), .I4(n4743), .O(n4744));
  LUT3 #(.INIT(8'h96)) lut_n4745 (.I0(n4733), .I1(n4736), .I2(n4737), .O(n4745));
  LUT3 #(.INIT(8'hE8)) lut_n4746 (.I0(n4741), .I1(n4744), .I2(n4745), .O(n4746));
  LUT3 #(.INIT(8'h96)) lut_n4747 (.I0(n4714), .I1(n4722), .I2(n4723), .O(n4747));
  LUT3 #(.INIT(8'hE8)) lut_n4748 (.I0(n4738), .I1(n4746), .I2(n4747), .O(n4748));
  LUT3 #(.INIT(8'hE8)) lut_n4749 (.I0(x2136), .I1(x2137), .I2(x2138), .O(n4749));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4750 (.I0(x2127), .I1(x2128), .I2(x2129), .I3(n4742), .I4(n4743), .O(n4750));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4751 (.I0(x2133), .I1(x2134), .I2(x2135), .I3(n4749), .I4(n4750), .O(n4751));
  LUT3 #(.INIT(8'hE8)) lut_n4752 (.I0(x2142), .I1(x2143), .I2(x2144), .O(n4752));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4753 (.I0(x2133), .I1(x2134), .I2(x2135), .I3(n4749), .I4(n4750), .O(n4753));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4754 (.I0(x2139), .I1(x2140), .I2(x2141), .I3(n4752), .I4(n4753), .O(n4754));
  LUT3 #(.INIT(8'h96)) lut_n4755 (.I0(n4741), .I1(n4744), .I2(n4745), .O(n4755));
  LUT3 #(.INIT(8'hE8)) lut_n4756 (.I0(n4751), .I1(n4754), .I2(n4755), .O(n4756));
  LUT3 #(.INIT(8'hE8)) lut_n4757 (.I0(x2148), .I1(x2149), .I2(x2150), .O(n4757));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4758 (.I0(x2139), .I1(x2140), .I2(x2141), .I3(n4752), .I4(n4753), .O(n4758));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4759 (.I0(x2145), .I1(x2146), .I2(x2147), .I3(n4757), .I4(n4758), .O(n4759));
  LUT3 #(.INIT(8'hE8)) lut_n4760 (.I0(x2154), .I1(x2155), .I2(x2156), .O(n4760));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4761 (.I0(x2145), .I1(x2146), .I2(x2147), .I3(n4757), .I4(n4758), .O(n4761));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4762 (.I0(x2151), .I1(x2152), .I2(x2153), .I3(n4760), .I4(n4761), .O(n4762));
  LUT3 #(.INIT(8'h96)) lut_n4763 (.I0(n4751), .I1(n4754), .I2(n4755), .O(n4763));
  LUT3 #(.INIT(8'hE8)) lut_n4764 (.I0(n4759), .I1(n4762), .I2(n4763), .O(n4764));
  LUT3 #(.INIT(8'h96)) lut_n4765 (.I0(n4738), .I1(n4746), .I2(n4747), .O(n4765));
  LUT3 #(.INIT(8'hE8)) lut_n4766 (.I0(n4756), .I1(n4764), .I2(n4765), .O(n4766));
  LUT3 #(.INIT(8'h96)) lut_n4767 (.I0(n4706), .I1(n4724), .I2(n4725), .O(n4767));
  LUT3 #(.INIT(8'hE8)) lut_n4768 (.I0(n4748), .I1(n4766), .I2(n4767), .O(n4768));
  LUT3 #(.INIT(8'hE8)) lut_n4769 (.I0(x2160), .I1(x2161), .I2(x2162), .O(n4769));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4770 (.I0(x2151), .I1(x2152), .I2(x2153), .I3(n4760), .I4(n4761), .O(n4770));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4771 (.I0(x2157), .I1(x2158), .I2(x2159), .I3(n4769), .I4(n4770), .O(n4771));
  LUT3 #(.INIT(8'hE8)) lut_n4772 (.I0(x2166), .I1(x2167), .I2(x2168), .O(n4772));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4773 (.I0(x2157), .I1(x2158), .I2(x2159), .I3(n4769), .I4(n4770), .O(n4773));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4774 (.I0(x2163), .I1(x2164), .I2(x2165), .I3(n4772), .I4(n4773), .O(n4774));
  LUT3 #(.INIT(8'h96)) lut_n4775 (.I0(n4759), .I1(n4762), .I2(n4763), .O(n4775));
  LUT3 #(.INIT(8'hE8)) lut_n4776 (.I0(n4771), .I1(n4774), .I2(n4775), .O(n4776));
  LUT3 #(.INIT(8'hE8)) lut_n4777 (.I0(x2172), .I1(x2173), .I2(x2174), .O(n4777));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4778 (.I0(x2163), .I1(x2164), .I2(x2165), .I3(n4772), .I4(n4773), .O(n4778));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4779 (.I0(x2169), .I1(x2170), .I2(x2171), .I3(n4777), .I4(n4778), .O(n4779));
  LUT3 #(.INIT(8'hE8)) lut_n4780 (.I0(x2178), .I1(x2179), .I2(x2180), .O(n4780));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4781 (.I0(x2169), .I1(x2170), .I2(x2171), .I3(n4777), .I4(n4778), .O(n4781));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4782 (.I0(x2175), .I1(x2176), .I2(x2177), .I3(n4780), .I4(n4781), .O(n4782));
  LUT3 #(.INIT(8'h96)) lut_n4783 (.I0(n4771), .I1(n4774), .I2(n4775), .O(n4783));
  LUT3 #(.INIT(8'hE8)) lut_n4784 (.I0(n4779), .I1(n4782), .I2(n4783), .O(n4784));
  LUT3 #(.INIT(8'h96)) lut_n4785 (.I0(n4756), .I1(n4764), .I2(n4765), .O(n4785));
  LUT3 #(.INIT(8'hE8)) lut_n4786 (.I0(n4776), .I1(n4784), .I2(n4785), .O(n4786));
  LUT3 #(.INIT(8'hE8)) lut_n4787 (.I0(x2184), .I1(x2185), .I2(x2186), .O(n4787));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4788 (.I0(x2175), .I1(x2176), .I2(x2177), .I3(n4780), .I4(n4781), .O(n4788));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4789 (.I0(x2181), .I1(x2182), .I2(x2183), .I3(n4787), .I4(n4788), .O(n4789));
  LUT3 #(.INIT(8'hE8)) lut_n4790 (.I0(x2190), .I1(x2191), .I2(x2192), .O(n4790));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4791 (.I0(x2181), .I1(x2182), .I2(x2183), .I3(n4787), .I4(n4788), .O(n4791));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4792 (.I0(x2187), .I1(x2188), .I2(x2189), .I3(n4790), .I4(n4791), .O(n4792));
  LUT3 #(.INIT(8'h96)) lut_n4793 (.I0(n4779), .I1(n4782), .I2(n4783), .O(n4793));
  LUT3 #(.INIT(8'hE8)) lut_n4794 (.I0(n4789), .I1(n4792), .I2(n4793), .O(n4794));
  LUT3 #(.INIT(8'hE8)) lut_n4795 (.I0(x2196), .I1(x2197), .I2(x2198), .O(n4795));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4796 (.I0(x2187), .I1(x2188), .I2(x2189), .I3(n4790), .I4(n4791), .O(n4796));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4797 (.I0(x2193), .I1(x2194), .I2(x2195), .I3(n4795), .I4(n4796), .O(n4797));
  LUT3 #(.INIT(8'hE8)) lut_n4798 (.I0(x2202), .I1(x2203), .I2(x2204), .O(n4798));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4799 (.I0(x2193), .I1(x2194), .I2(x2195), .I3(n4795), .I4(n4796), .O(n4799));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4800 (.I0(x2199), .I1(x2200), .I2(x2201), .I3(n4798), .I4(n4799), .O(n4800));
  LUT3 #(.INIT(8'h96)) lut_n4801 (.I0(n4789), .I1(n4792), .I2(n4793), .O(n4801));
  LUT3 #(.INIT(8'hE8)) lut_n4802 (.I0(n4797), .I1(n4800), .I2(n4801), .O(n4802));
  LUT3 #(.INIT(8'h96)) lut_n4803 (.I0(n4776), .I1(n4784), .I2(n4785), .O(n4803));
  LUT3 #(.INIT(8'hE8)) lut_n4804 (.I0(n4794), .I1(n4802), .I2(n4803), .O(n4804));
  LUT3 #(.INIT(8'h96)) lut_n4805 (.I0(n4748), .I1(n4766), .I2(n4767), .O(n4805));
  LUT3 #(.INIT(8'hE8)) lut_n4806 (.I0(n4786), .I1(n4804), .I2(n4805), .O(n4806));
  LUT3 #(.INIT(8'h96)) lut_n4807 (.I0(n4688), .I1(n4726), .I2(n4727), .O(n4807));
  LUT3 #(.INIT(8'hE8)) lut_n4808 (.I0(n4768), .I1(n4806), .I2(n4807), .O(n4808));
  LUT3 #(.INIT(8'hE8)) lut_n4809 (.I0(x2208), .I1(x2209), .I2(x2210), .O(n4809));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4810 (.I0(x2199), .I1(x2200), .I2(x2201), .I3(n4798), .I4(n4799), .O(n4810));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4811 (.I0(x2205), .I1(x2206), .I2(x2207), .I3(n4809), .I4(n4810), .O(n4811));
  LUT3 #(.INIT(8'hE8)) lut_n4812 (.I0(x2214), .I1(x2215), .I2(x2216), .O(n4812));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4813 (.I0(x2205), .I1(x2206), .I2(x2207), .I3(n4809), .I4(n4810), .O(n4813));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4814 (.I0(x2211), .I1(x2212), .I2(x2213), .I3(n4812), .I4(n4813), .O(n4814));
  LUT3 #(.INIT(8'h96)) lut_n4815 (.I0(n4797), .I1(n4800), .I2(n4801), .O(n4815));
  LUT3 #(.INIT(8'hE8)) lut_n4816 (.I0(n4811), .I1(n4814), .I2(n4815), .O(n4816));
  LUT3 #(.INIT(8'hE8)) lut_n4817 (.I0(x2220), .I1(x2221), .I2(x2222), .O(n4817));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4818 (.I0(x2211), .I1(x2212), .I2(x2213), .I3(n4812), .I4(n4813), .O(n4818));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4819 (.I0(x2217), .I1(x2218), .I2(x2219), .I3(n4817), .I4(n4818), .O(n4819));
  LUT3 #(.INIT(8'hE8)) lut_n4820 (.I0(x2226), .I1(x2227), .I2(x2228), .O(n4820));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4821 (.I0(x2217), .I1(x2218), .I2(x2219), .I3(n4817), .I4(n4818), .O(n4821));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4822 (.I0(x2223), .I1(x2224), .I2(x2225), .I3(n4820), .I4(n4821), .O(n4822));
  LUT3 #(.INIT(8'h96)) lut_n4823 (.I0(n4811), .I1(n4814), .I2(n4815), .O(n4823));
  LUT3 #(.INIT(8'hE8)) lut_n4824 (.I0(n4819), .I1(n4822), .I2(n4823), .O(n4824));
  LUT3 #(.INIT(8'h96)) lut_n4825 (.I0(n4794), .I1(n4802), .I2(n4803), .O(n4825));
  LUT3 #(.INIT(8'hE8)) lut_n4826 (.I0(n4816), .I1(n4824), .I2(n4825), .O(n4826));
  LUT3 #(.INIT(8'hE8)) lut_n4827 (.I0(x2232), .I1(x2233), .I2(x2234), .O(n4827));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4828 (.I0(x2223), .I1(x2224), .I2(x2225), .I3(n4820), .I4(n4821), .O(n4828));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4829 (.I0(x2229), .I1(x2230), .I2(x2231), .I3(n4827), .I4(n4828), .O(n4829));
  LUT3 #(.INIT(8'hE8)) lut_n4830 (.I0(x2238), .I1(x2239), .I2(x2240), .O(n4830));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4831 (.I0(x2229), .I1(x2230), .I2(x2231), .I3(n4827), .I4(n4828), .O(n4831));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4832 (.I0(x2235), .I1(x2236), .I2(x2237), .I3(n4830), .I4(n4831), .O(n4832));
  LUT3 #(.INIT(8'h96)) lut_n4833 (.I0(n4819), .I1(n4822), .I2(n4823), .O(n4833));
  LUT3 #(.INIT(8'hE8)) lut_n4834 (.I0(n4829), .I1(n4832), .I2(n4833), .O(n4834));
  LUT3 #(.INIT(8'hE8)) lut_n4835 (.I0(x2244), .I1(x2245), .I2(x2246), .O(n4835));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4836 (.I0(x2235), .I1(x2236), .I2(x2237), .I3(n4830), .I4(n4831), .O(n4836));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4837 (.I0(x2241), .I1(x2242), .I2(x2243), .I3(n4835), .I4(n4836), .O(n4837));
  LUT3 #(.INIT(8'hE8)) lut_n4838 (.I0(x2250), .I1(x2251), .I2(x2252), .O(n4838));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4839 (.I0(x2241), .I1(x2242), .I2(x2243), .I3(n4835), .I4(n4836), .O(n4839));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4840 (.I0(x2247), .I1(x2248), .I2(x2249), .I3(n4838), .I4(n4839), .O(n4840));
  LUT3 #(.INIT(8'h96)) lut_n4841 (.I0(n4829), .I1(n4832), .I2(n4833), .O(n4841));
  LUT3 #(.INIT(8'hE8)) lut_n4842 (.I0(n4837), .I1(n4840), .I2(n4841), .O(n4842));
  LUT3 #(.INIT(8'h96)) lut_n4843 (.I0(n4816), .I1(n4824), .I2(n4825), .O(n4843));
  LUT3 #(.INIT(8'hE8)) lut_n4844 (.I0(n4834), .I1(n4842), .I2(n4843), .O(n4844));
  LUT3 #(.INIT(8'h96)) lut_n4845 (.I0(n4786), .I1(n4804), .I2(n4805), .O(n4845));
  LUT3 #(.INIT(8'hE8)) lut_n4846 (.I0(n4826), .I1(n4844), .I2(n4845), .O(n4846));
  LUT3 #(.INIT(8'hE8)) lut_n4847 (.I0(x2256), .I1(x2257), .I2(x2258), .O(n4847));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4848 (.I0(x2247), .I1(x2248), .I2(x2249), .I3(n4838), .I4(n4839), .O(n4848));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4849 (.I0(x2253), .I1(x2254), .I2(x2255), .I3(n4847), .I4(n4848), .O(n4849));
  LUT3 #(.INIT(8'hE8)) lut_n4850 (.I0(x2262), .I1(x2263), .I2(x2264), .O(n4850));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4851 (.I0(x2253), .I1(x2254), .I2(x2255), .I3(n4847), .I4(n4848), .O(n4851));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4852 (.I0(x2259), .I1(x2260), .I2(x2261), .I3(n4850), .I4(n4851), .O(n4852));
  LUT3 #(.INIT(8'h96)) lut_n4853 (.I0(n4837), .I1(n4840), .I2(n4841), .O(n4853));
  LUT3 #(.INIT(8'hE8)) lut_n4854 (.I0(n4849), .I1(n4852), .I2(n4853), .O(n4854));
  LUT3 #(.INIT(8'hE8)) lut_n4855 (.I0(x2268), .I1(x2269), .I2(x2270), .O(n4855));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4856 (.I0(x2259), .I1(x2260), .I2(x2261), .I3(n4850), .I4(n4851), .O(n4856));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4857 (.I0(x2265), .I1(x2266), .I2(x2267), .I3(n4855), .I4(n4856), .O(n4857));
  LUT3 #(.INIT(8'hE8)) lut_n4858 (.I0(x2274), .I1(x2275), .I2(x2276), .O(n4858));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4859 (.I0(x2265), .I1(x2266), .I2(x2267), .I3(n4855), .I4(n4856), .O(n4859));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4860 (.I0(x2271), .I1(x2272), .I2(x2273), .I3(n4858), .I4(n4859), .O(n4860));
  LUT3 #(.INIT(8'h96)) lut_n4861 (.I0(n4849), .I1(n4852), .I2(n4853), .O(n4861));
  LUT3 #(.INIT(8'hE8)) lut_n4862 (.I0(n4857), .I1(n4860), .I2(n4861), .O(n4862));
  LUT3 #(.INIT(8'h96)) lut_n4863 (.I0(n4834), .I1(n4842), .I2(n4843), .O(n4863));
  LUT3 #(.INIT(8'hE8)) lut_n4864 (.I0(n4854), .I1(n4862), .I2(n4863), .O(n4864));
  LUT3 #(.INIT(8'hE8)) lut_n4865 (.I0(x2280), .I1(x2281), .I2(x2282), .O(n4865));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4866 (.I0(x2271), .I1(x2272), .I2(x2273), .I3(n4858), .I4(n4859), .O(n4866));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4867 (.I0(x2277), .I1(x2278), .I2(x2279), .I3(n4865), .I4(n4866), .O(n4867));
  LUT3 #(.INIT(8'hE8)) lut_n4868 (.I0(x2286), .I1(x2287), .I2(x2288), .O(n4868));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4869 (.I0(x2277), .I1(x2278), .I2(x2279), .I3(n4865), .I4(n4866), .O(n4869));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4870 (.I0(x2283), .I1(x2284), .I2(x2285), .I3(n4868), .I4(n4869), .O(n4870));
  LUT3 #(.INIT(8'h96)) lut_n4871 (.I0(n4857), .I1(n4860), .I2(n4861), .O(n4871));
  LUT3 #(.INIT(8'hE8)) lut_n4872 (.I0(n4867), .I1(n4870), .I2(n4871), .O(n4872));
  LUT3 #(.INIT(8'hE8)) lut_n4873 (.I0(x2292), .I1(x2293), .I2(x2294), .O(n4873));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4874 (.I0(x2283), .I1(x2284), .I2(x2285), .I3(n4868), .I4(n4869), .O(n4874));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4875 (.I0(x2289), .I1(x2290), .I2(x2291), .I3(n4873), .I4(n4874), .O(n4875));
  LUT3 #(.INIT(8'hE8)) lut_n4876 (.I0(x2298), .I1(x2299), .I2(x2300), .O(n4876));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4877 (.I0(x2289), .I1(x2290), .I2(x2291), .I3(n4873), .I4(n4874), .O(n4877));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4878 (.I0(x2295), .I1(x2296), .I2(x2297), .I3(n4876), .I4(n4877), .O(n4878));
  LUT3 #(.INIT(8'h96)) lut_n4879 (.I0(n4867), .I1(n4870), .I2(n4871), .O(n4879));
  LUT3 #(.INIT(8'hE8)) lut_n4880 (.I0(n4875), .I1(n4878), .I2(n4879), .O(n4880));
  LUT3 #(.INIT(8'h96)) lut_n4881 (.I0(n4854), .I1(n4862), .I2(n4863), .O(n4881));
  LUT3 #(.INIT(8'hE8)) lut_n4882 (.I0(n4872), .I1(n4880), .I2(n4881), .O(n4882));
  LUT3 #(.INIT(8'h96)) lut_n4883 (.I0(n4826), .I1(n4844), .I2(n4845), .O(n4883));
  LUT3 #(.INIT(8'hE8)) lut_n4884 (.I0(n4864), .I1(n4882), .I2(n4883), .O(n4884));
  LUT3 #(.INIT(8'h96)) lut_n4885 (.I0(n4768), .I1(n4806), .I2(n4807), .O(n4885));
  LUT3 #(.INIT(8'hE8)) lut_n4886 (.I0(n4846), .I1(n4884), .I2(n4885), .O(n4886));
  LUT3 #(.INIT(8'h96)) lut_n4887 (.I0(n4650), .I1(n4728), .I2(n4729), .O(n4887));
  LUT3 #(.INIT(8'hE8)) lut_n4888 (.I0(n4808), .I1(n4886), .I2(n4887), .O(n4888));
  LUT3 #(.INIT(8'h96)) lut_n4889 (.I0(n4412), .I1(n4570), .I2(n4571), .O(n4889));
  LUT3 #(.INIT(8'hE8)) lut_n4890 (.I0(n4730), .I1(n4888), .I2(n4889), .O(n4890));
  LUT3 #(.INIT(8'h96)) lut_n4891 (.I0(n3617), .I1(n3935), .I2(n4253), .O(n4891));
  LUT3 #(.INIT(8'hE8)) lut_n4892 (.I0(n4572), .I1(n4890), .I2(n4891), .O(n4892));
  LUT3 #(.INIT(8'hE8)) lut_n4893 (.I0(x2304), .I1(x2305), .I2(x2306), .O(n4893));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4894 (.I0(x2295), .I1(x2296), .I2(x2297), .I3(n4876), .I4(n4877), .O(n4894));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4895 (.I0(x2301), .I1(x2302), .I2(x2303), .I3(n4893), .I4(n4894), .O(n4895));
  LUT3 #(.INIT(8'hE8)) lut_n4896 (.I0(x2310), .I1(x2311), .I2(x2312), .O(n4896));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4897 (.I0(x2301), .I1(x2302), .I2(x2303), .I3(n4893), .I4(n4894), .O(n4897));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4898 (.I0(x2307), .I1(x2308), .I2(x2309), .I3(n4896), .I4(n4897), .O(n4898));
  LUT3 #(.INIT(8'h96)) lut_n4899 (.I0(n4875), .I1(n4878), .I2(n4879), .O(n4899));
  LUT3 #(.INIT(8'hE8)) lut_n4900 (.I0(n4895), .I1(n4898), .I2(n4899), .O(n4900));
  LUT3 #(.INIT(8'hE8)) lut_n4901 (.I0(x2316), .I1(x2317), .I2(x2318), .O(n4901));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4902 (.I0(x2307), .I1(x2308), .I2(x2309), .I3(n4896), .I4(n4897), .O(n4902));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4903 (.I0(x2313), .I1(x2314), .I2(x2315), .I3(n4901), .I4(n4902), .O(n4903));
  LUT3 #(.INIT(8'hE8)) lut_n4904 (.I0(x2322), .I1(x2323), .I2(x2324), .O(n4904));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4905 (.I0(x2313), .I1(x2314), .I2(x2315), .I3(n4901), .I4(n4902), .O(n4905));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4906 (.I0(x2319), .I1(x2320), .I2(x2321), .I3(n4904), .I4(n4905), .O(n4906));
  LUT3 #(.INIT(8'h96)) lut_n4907 (.I0(n4895), .I1(n4898), .I2(n4899), .O(n4907));
  LUT3 #(.INIT(8'hE8)) lut_n4908 (.I0(n4903), .I1(n4906), .I2(n4907), .O(n4908));
  LUT3 #(.INIT(8'h96)) lut_n4909 (.I0(n4872), .I1(n4880), .I2(n4881), .O(n4909));
  LUT3 #(.INIT(8'hE8)) lut_n4910 (.I0(n4900), .I1(n4908), .I2(n4909), .O(n4910));
  LUT3 #(.INIT(8'hE8)) lut_n4911 (.I0(x2328), .I1(x2329), .I2(x2330), .O(n4911));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4912 (.I0(x2319), .I1(x2320), .I2(x2321), .I3(n4904), .I4(n4905), .O(n4912));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4913 (.I0(x2325), .I1(x2326), .I2(x2327), .I3(n4911), .I4(n4912), .O(n4913));
  LUT3 #(.INIT(8'hE8)) lut_n4914 (.I0(x2334), .I1(x2335), .I2(x2336), .O(n4914));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4915 (.I0(x2325), .I1(x2326), .I2(x2327), .I3(n4911), .I4(n4912), .O(n4915));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4916 (.I0(x2331), .I1(x2332), .I2(x2333), .I3(n4914), .I4(n4915), .O(n4916));
  LUT3 #(.INIT(8'h96)) lut_n4917 (.I0(n4903), .I1(n4906), .I2(n4907), .O(n4917));
  LUT3 #(.INIT(8'hE8)) lut_n4918 (.I0(n4913), .I1(n4916), .I2(n4917), .O(n4918));
  LUT3 #(.INIT(8'hE8)) lut_n4919 (.I0(x2340), .I1(x2341), .I2(x2342), .O(n4919));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4920 (.I0(x2331), .I1(x2332), .I2(x2333), .I3(n4914), .I4(n4915), .O(n4920));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4921 (.I0(x2337), .I1(x2338), .I2(x2339), .I3(n4919), .I4(n4920), .O(n4921));
  LUT3 #(.INIT(8'hE8)) lut_n4922 (.I0(x2346), .I1(x2347), .I2(x2348), .O(n4922));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4923 (.I0(x2337), .I1(x2338), .I2(x2339), .I3(n4919), .I4(n4920), .O(n4923));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4924 (.I0(x2343), .I1(x2344), .I2(x2345), .I3(n4922), .I4(n4923), .O(n4924));
  LUT3 #(.INIT(8'h96)) lut_n4925 (.I0(n4913), .I1(n4916), .I2(n4917), .O(n4925));
  LUT3 #(.INIT(8'hE8)) lut_n4926 (.I0(n4921), .I1(n4924), .I2(n4925), .O(n4926));
  LUT3 #(.INIT(8'h96)) lut_n4927 (.I0(n4900), .I1(n4908), .I2(n4909), .O(n4927));
  LUT3 #(.INIT(8'hE8)) lut_n4928 (.I0(n4918), .I1(n4926), .I2(n4927), .O(n4928));
  LUT3 #(.INIT(8'h96)) lut_n4929 (.I0(n4864), .I1(n4882), .I2(n4883), .O(n4929));
  LUT3 #(.INIT(8'hE8)) lut_n4930 (.I0(n4910), .I1(n4928), .I2(n4929), .O(n4930));
  LUT3 #(.INIT(8'hE8)) lut_n4931 (.I0(x2352), .I1(x2353), .I2(x2354), .O(n4931));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4932 (.I0(x2343), .I1(x2344), .I2(x2345), .I3(n4922), .I4(n4923), .O(n4932));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4933 (.I0(x2349), .I1(x2350), .I2(x2351), .I3(n4931), .I4(n4932), .O(n4933));
  LUT3 #(.INIT(8'hE8)) lut_n4934 (.I0(x2358), .I1(x2359), .I2(x2360), .O(n4934));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4935 (.I0(x2349), .I1(x2350), .I2(x2351), .I3(n4931), .I4(n4932), .O(n4935));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4936 (.I0(x2355), .I1(x2356), .I2(x2357), .I3(n4934), .I4(n4935), .O(n4936));
  LUT3 #(.INIT(8'h96)) lut_n4937 (.I0(n4921), .I1(n4924), .I2(n4925), .O(n4937));
  LUT3 #(.INIT(8'hE8)) lut_n4938 (.I0(n4933), .I1(n4936), .I2(n4937), .O(n4938));
  LUT3 #(.INIT(8'hE8)) lut_n4939 (.I0(x2364), .I1(x2365), .I2(x2366), .O(n4939));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4940 (.I0(x2355), .I1(x2356), .I2(x2357), .I3(n4934), .I4(n4935), .O(n4940));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4941 (.I0(x2361), .I1(x2362), .I2(x2363), .I3(n4939), .I4(n4940), .O(n4941));
  LUT3 #(.INIT(8'hE8)) lut_n4942 (.I0(x2370), .I1(x2371), .I2(x2372), .O(n4942));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4943 (.I0(x2361), .I1(x2362), .I2(x2363), .I3(n4939), .I4(n4940), .O(n4943));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4944 (.I0(x2367), .I1(x2368), .I2(x2369), .I3(n4942), .I4(n4943), .O(n4944));
  LUT3 #(.INIT(8'h96)) lut_n4945 (.I0(n4933), .I1(n4936), .I2(n4937), .O(n4945));
  LUT3 #(.INIT(8'hE8)) lut_n4946 (.I0(n4941), .I1(n4944), .I2(n4945), .O(n4946));
  LUT3 #(.INIT(8'h96)) lut_n4947 (.I0(n4918), .I1(n4926), .I2(n4927), .O(n4947));
  LUT3 #(.INIT(8'hE8)) lut_n4948 (.I0(n4938), .I1(n4946), .I2(n4947), .O(n4948));
  LUT3 #(.INIT(8'hE8)) lut_n4949 (.I0(x2376), .I1(x2377), .I2(x2378), .O(n4949));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4950 (.I0(x2367), .I1(x2368), .I2(x2369), .I3(n4942), .I4(n4943), .O(n4950));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4951 (.I0(x2373), .I1(x2374), .I2(x2375), .I3(n4949), .I4(n4950), .O(n4951));
  LUT3 #(.INIT(8'hE8)) lut_n4952 (.I0(x2382), .I1(x2383), .I2(x2384), .O(n4952));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4953 (.I0(x2373), .I1(x2374), .I2(x2375), .I3(n4949), .I4(n4950), .O(n4953));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4954 (.I0(x2379), .I1(x2380), .I2(x2381), .I3(n4952), .I4(n4953), .O(n4954));
  LUT3 #(.INIT(8'h96)) lut_n4955 (.I0(n4941), .I1(n4944), .I2(n4945), .O(n4955));
  LUT3 #(.INIT(8'hE8)) lut_n4956 (.I0(n4951), .I1(n4954), .I2(n4955), .O(n4956));
  LUT3 #(.INIT(8'hE8)) lut_n4957 (.I0(x2388), .I1(x2389), .I2(x2390), .O(n4957));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4958 (.I0(x2379), .I1(x2380), .I2(x2381), .I3(n4952), .I4(n4953), .O(n4958));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4959 (.I0(x2385), .I1(x2386), .I2(x2387), .I3(n4957), .I4(n4958), .O(n4959));
  LUT3 #(.INIT(8'hE8)) lut_n4960 (.I0(x2394), .I1(x2395), .I2(x2396), .O(n4960));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4961 (.I0(x2385), .I1(x2386), .I2(x2387), .I3(n4957), .I4(n4958), .O(n4961));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4962 (.I0(x2391), .I1(x2392), .I2(x2393), .I3(n4960), .I4(n4961), .O(n4962));
  LUT3 #(.INIT(8'h96)) lut_n4963 (.I0(n4951), .I1(n4954), .I2(n4955), .O(n4963));
  LUT3 #(.INIT(8'hE8)) lut_n4964 (.I0(n4959), .I1(n4962), .I2(n4963), .O(n4964));
  LUT3 #(.INIT(8'h96)) lut_n4965 (.I0(n4938), .I1(n4946), .I2(n4947), .O(n4965));
  LUT3 #(.INIT(8'hE8)) lut_n4966 (.I0(n4956), .I1(n4964), .I2(n4965), .O(n4966));
  LUT3 #(.INIT(8'h96)) lut_n4967 (.I0(n4910), .I1(n4928), .I2(n4929), .O(n4967));
  LUT3 #(.INIT(8'hE8)) lut_n4968 (.I0(n4948), .I1(n4966), .I2(n4967), .O(n4968));
  LUT3 #(.INIT(8'h96)) lut_n4969 (.I0(n4846), .I1(n4884), .I2(n4885), .O(n4969));
  LUT3 #(.INIT(8'hE8)) lut_n4970 (.I0(n4930), .I1(n4968), .I2(n4969), .O(n4970));
  LUT3 #(.INIT(8'hE8)) lut_n4971 (.I0(x2400), .I1(x2401), .I2(x2402), .O(n4971));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4972 (.I0(x2391), .I1(x2392), .I2(x2393), .I3(n4960), .I4(n4961), .O(n4972));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4973 (.I0(x2397), .I1(x2398), .I2(x2399), .I3(n4971), .I4(n4972), .O(n4973));
  LUT3 #(.INIT(8'hE8)) lut_n4974 (.I0(x2406), .I1(x2407), .I2(x2408), .O(n4974));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4975 (.I0(x2397), .I1(x2398), .I2(x2399), .I3(n4971), .I4(n4972), .O(n4975));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4976 (.I0(x2403), .I1(x2404), .I2(x2405), .I3(n4974), .I4(n4975), .O(n4976));
  LUT3 #(.INIT(8'h96)) lut_n4977 (.I0(n4959), .I1(n4962), .I2(n4963), .O(n4977));
  LUT3 #(.INIT(8'hE8)) lut_n4978 (.I0(n4973), .I1(n4976), .I2(n4977), .O(n4978));
  LUT3 #(.INIT(8'hE8)) lut_n4979 (.I0(x2412), .I1(x2413), .I2(x2414), .O(n4979));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4980 (.I0(x2403), .I1(x2404), .I2(x2405), .I3(n4974), .I4(n4975), .O(n4980));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4981 (.I0(x2409), .I1(x2410), .I2(x2411), .I3(n4979), .I4(n4980), .O(n4981));
  LUT3 #(.INIT(8'hE8)) lut_n4982 (.I0(x2418), .I1(x2419), .I2(x2420), .O(n4982));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4983 (.I0(x2409), .I1(x2410), .I2(x2411), .I3(n4979), .I4(n4980), .O(n4983));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4984 (.I0(x2415), .I1(x2416), .I2(x2417), .I3(n4982), .I4(n4983), .O(n4984));
  LUT3 #(.INIT(8'h96)) lut_n4985 (.I0(n4973), .I1(n4976), .I2(n4977), .O(n4985));
  LUT3 #(.INIT(8'hE8)) lut_n4986 (.I0(n4981), .I1(n4984), .I2(n4985), .O(n4986));
  LUT3 #(.INIT(8'h96)) lut_n4987 (.I0(n4956), .I1(n4964), .I2(n4965), .O(n4987));
  LUT3 #(.INIT(8'hE8)) lut_n4988 (.I0(n4978), .I1(n4986), .I2(n4987), .O(n4988));
  LUT3 #(.INIT(8'hE8)) lut_n4989 (.I0(x2424), .I1(x2425), .I2(x2426), .O(n4989));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4990 (.I0(x2415), .I1(x2416), .I2(x2417), .I3(n4982), .I4(n4983), .O(n4990));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4991 (.I0(x2421), .I1(x2422), .I2(x2423), .I3(n4989), .I4(n4990), .O(n4991));
  LUT3 #(.INIT(8'hE8)) lut_n4992 (.I0(x2430), .I1(x2431), .I2(x2432), .O(n4992));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4993 (.I0(x2421), .I1(x2422), .I2(x2423), .I3(n4989), .I4(n4990), .O(n4993));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4994 (.I0(x2427), .I1(x2428), .I2(x2429), .I3(n4992), .I4(n4993), .O(n4994));
  LUT3 #(.INIT(8'h96)) lut_n4995 (.I0(n4981), .I1(n4984), .I2(n4985), .O(n4995));
  LUT3 #(.INIT(8'hE8)) lut_n4996 (.I0(n4991), .I1(n4994), .I2(n4995), .O(n4996));
  LUT3 #(.INIT(8'hE8)) lut_n4997 (.I0(x2436), .I1(x2437), .I2(x2438), .O(n4997));
  LUT5 #(.INIT(32'hE81717E8)) lut_n4998 (.I0(x2427), .I1(x2428), .I2(x2429), .I3(n4992), .I4(n4993), .O(n4998));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n4999 (.I0(x2433), .I1(x2434), .I2(x2435), .I3(n4997), .I4(n4998), .O(n4999));
  LUT3 #(.INIT(8'hE8)) lut_n5000 (.I0(x2442), .I1(x2443), .I2(x2444), .O(n5000));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5001 (.I0(x2433), .I1(x2434), .I2(x2435), .I3(n4997), .I4(n4998), .O(n5001));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5002 (.I0(x2439), .I1(x2440), .I2(x2441), .I3(n5000), .I4(n5001), .O(n5002));
  LUT3 #(.INIT(8'h96)) lut_n5003 (.I0(n4991), .I1(n4994), .I2(n4995), .O(n5003));
  LUT3 #(.INIT(8'hE8)) lut_n5004 (.I0(n4999), .I1(n5002), .I2(n5003), .O(n5004));
  LUT3 #(.INIT(8'h96)) lut_n5005 (.I0(n4978), .I1(n4986), .I2(n4987), .O(n5005));
  LUT3 #(.INIT(8'hE8)) lut_n5006 (.I0(n4996), .I1(n5004), .I2(n5005), .O(n5006));
  LUT3 #(.INIT(8'h96)) lut_n5007 (.I0(n4948), .I1(n4966), .I2(n4967), .O(n5007));
  LUT3 #(.INIT(8'hE8)) lut_n5008 (.I0(n4988), .I1(n5006), .I2(n5007), .O(n5008));
  LUT3 #(.INIT(8'hE8)) lut_n5009 (.I0(x2448), .I1(x2449), .I2(x2450), .O(n5009));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5010 (.I0(x2439), .I1(x2440), .I2(x2441), .I3(n5000), .I4(n5001), .O(n5010));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5011 (.I0(x2445), .I1(x2446), .I2(x2447), .I3(n5009), .I4(n5010), .O(n5011));
  LUT3 #(.INIT(8'hE8)) lut_n5012 (.I0(x2454), .I1(x2455), .I2(x2456), .O(n5012));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5013 (.I0(x2445), .I1(x2446), .I2(x2447), .I3(n5009), .I4(n5010), .O(n5013));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5014 (.I0(x2451), .I1(x2452), .I2(x2453), .I3(n5012), .I4(n5013), .O(n5014));
  LUT3 #(.INIT(8'h96)) lut_n5015 (.I0(n4999), .I1(n5002), .I2(n5003), .O(n5015));
  LUT3 #(.INIT(8'hE8)) lut_n5016 (.I0(n5011), .I1(n5014), .I2(n5015), .O(n5016));
  LUT3 #(.INIT(8'hE8)) lut_n5017 (.I0(x2460), .I1(x2461), .I2(x2462), .O(n5017));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5018 (.I0(x2451), .I1(x2452), .I2(x2453), .I3(n5012), .I4(n5013), .O(n5018));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5019 (.I0(x2457), .I1(x2458), .I2(x2459), .I3(n5017), .I4(n5018), .O(n5019));
  LUT3 #(.INIT(8'hE8)) lut_n5020 (.I0(x2466), .I1(x2467), .I2(x2468), .O(n5020));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5021 (.I0(x2457), .I1(x2458), .I2(x2459), .I3(n5017), .I4(n5018), .O(n5021));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5022 (.I0(x2463), .I1(x2464), .I2(x2465), .I3(n5020), .I4(n5021), .O(n5022));
  LUT3 #(.INIT(8'h96)) lut_n5023 (.I0(n5011), .I1(n5014), .I2(n5015), .O(n5023));
  LUT3 #(.INIT(8'hE8)) lut_n5024 (.I0(n5019), .I1(n5022), .I2(n5023), .O(n5024));
  LUT3 #(.INIT(8'h96)) lut_n5025 (.I0(n4996), .I1(n5004), .I2(n5005), .O(n5025));
  LUT3 #(.INIT(8'hE8)) lut_n5026 (.I0(n5016), .I1(n5024), .I2(n5025), .O(n5026));
  LUT3 #(.INIT(8'hE8)) lut_n5027 (.I0(x2472), .I1(x2473), .I2(x2474), .O(n5027));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5028 (.I0(x2463), .I1(x2464), .I2(x2465), .I3(n5020), .I4(n5021), .O(n5028));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5029 (.I0(x2469), .I1(x2470), .I2(x2471), .I3(n5027), .I4(n5028), .O(n5029));
  LUT3 #(.INIT(8'hE8)) lut_n5030 (.I0(x2478), .I1(x2479), .I2(x2480), .O(n5030));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5031 (.I0(x2469), .I1(x2470), .I2(x2471), .I3(n5027), .I4(n5028), .O(n5031));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5032 (.I0(x2475), .I1(x2476), .I2(x2477), .I3(n5030), .I4(n5031), .O(n5032));
  LUT3 #(.INIT(8'h96)) lut_n5033 (.I0(n5019), .I1(n5022), .I2(n5023), .O(n5033));
  LUT3 #(.INIT(8'hE8)) lut_n5034 (.I0(n5029), .I1(n5032), .I2(n5033), .O(n5034));
  LUT3 #(.INIT(8'hE8)) lut_n5035 (.I0(x2484), .I1(x2485), .I2(x2486), .O(n5035));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5036 (.I0(x2475), .I1(x2476), .I2(x2477), .I3(n5030), .I4(n5031), .O(n5036));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5037 (.I0(x2481), .I1(x2482), .I2(x2483), .I3(n5035), .I4(n5036), .O(n5037));
  LUT3 #(.INIT(8'hE8)) lut_n5038 (.I0(x2490), .I1(x2491), .I2(x2492), .O(n5038));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5039 (.I0(x2481), .I1(x2482), .I2(x2483), .I3(n5035), .I4(n5036), .O(n5039));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5040 (.I0(x2487), .I1(x2488), .I2(x2489), .I3(n5038), .I4(n5039), .O(n5040));
  LUT3 #(.INIT(8'h96)) lut_n5041 (.I0(n5029), .I1(n5032), .I2(n5033), .O(n5041));
  LUT3 #(.INIT(8'hE8)) lut_n5042 (.I0(n5037), .I1(n5040), .I2(n5041), .O(n5042));
  LUT3 #(.INIT(8'h96)) lut_n5043 (.I0(n5016), .I1(n5024), .I2(n5025), .O(n5043));
  LUT3 #(.INIT(8'hE8)) lut_n5044 (.I0(n5034), .I1(n5042), .I2(n5043), .O(n5044));
  LUT3 #(.INIT(8'h96)) lut_n5045 (.I0(n4988), .I1(n5006), .I2(n5007), .O(n5045));
  LUT3 #(.INIT(8'hE8)) lut_n5046 (.I0(n5026), .I1(n5044), .I2(n5045), .O(n5046));
  LUT3 #(.INIT(8'h96)) lut_n5047 (.I0(n4930), .I1(n4968), .I2(n4969), .O(n5047));
  LUT3 #(.INIT(8'hE8)) lut_n5048 (.I0(n5008), .I1(n5046), .I2(n5047), .O(n5048));
  LUT3 #(.INIT(8'h96)) lut_n5049 (.I0(n4808), .I1(n4886), .I2(n4887), .O(n5049));
  LUT3 #(.INIT(8'hE8)) lut_n5050 (.I0(n4970), .I1(n5048), .I2(n5049), .O(n5050));
  LUT3 #(.INIT(8'hE8)) lut_n5051 (.I0(x2496), .I1(x2497), .I2(x2498), .O(n5051));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5052 (.I0(x2487), .I1(x2488), .I2(x2489), .I3(n5038), .I4(n5039), .O(n5052));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5053 (.I0(x2493), .I1(x2494), .I2(x2495), .I3(n5051), .I4(n5052), .O(n5053));
  LUT3 #(.INIT(8'hE8)) lut_n5054 (.I0(x2502), .I1(x2503), .I2(x2504), .O(n5054));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5055 (.I0(x2493), .I1(x2494), .I2(x2495), .I3(n5051), .I4(n5052), .O(n5055));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5056 (.I0(x2499), .I1(x2500), .I2(x2501), .I3(n5054), .I4(n5055), .O(n5056));
  LUT3 #(.INIT(8'h96)) lut_n5057 (.I0(n5037), .I1(n5040), .I2(n5041), .O(n5057));
  LUT3 #(.INIT(8'hE8)) lut_n5058 (.I0(n5053), .I1(n5056), .I2(n5057), .O(n5058));
  LUT3 #(.INIT(8'hE8)) lut_n5059 (.I0(x2508), .I1(x2509), .I2(x2510), .O(n5059));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5060 (.I0(x2499), .I1(x2500), .I2(x2501), .I3(n5054), .I4(n5055), .O(n5060));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5061 (.I0(x2505), .I1(x2506), .I2(x2507), .I3(n5059), .I4(n5060), .O(n5061));
  LUT3 #(.INIT(8'hE8)) lut_n5062 (.I0(x2514), .I1(x2515), .I2(x2516), .O(n5062));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5063 (.I0(x2505), .I1(x2506), .I2(x2507), .I3(n5059), .I4(n5060), .O(n5063));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5064 (.I0(x2511), .I1(x2512), .I2(x2513), .I3(n5062), .I4(n5063), .O(n5064));
  LUT3 #(.INIT(8'h96)) lut_n5065 (.I0(n5053), .I1(n5056), .I2(n5057), .O(n5065));
  LUT3 #(.INIT(8'hE8)) lut_n5066 (.I0(n5061), .I1(n5064), .I2(n5065), .O(n5066));
  LUT3 #(.INIT(8'h96)) lut_n5067 (.I0(n5034), .I1(n5042), .I2(n5043), .O(n5067));
  LUT3 #(.INIT(8'hE8)) lut_n5068 (.I0(n5058), .I1(n5066), .I2(n5067), .O(n5068));
  LUT3 #(.INIT(8'hE8)) lut_n5069 (.I0(x2520), .I1(x2521), .I2(x2522), .O(n5069));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5070 (.I0(x2511), .I1(x2512), .I2(x2513), .I3(n5062), .I4(n5063), .O(n5070));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5071 (.I0(x2517), .I1(x2518), .I2(x2519), .I3(n5069), .I4(n5070), .O(n5071));
  LUT3 #(.INIT(8'hE8)) lut_n5072 (.I0(x2526), .I1(x2527), .I2(x2528), .O(n5072));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5073 (.I0(x2517), .I1(x2518), .I2(x2519), .I3(n5069), .I4(n5070), .O(n5073));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5074 (.I0(x2523), .I1(x2524), .I2(x2525), .I3(n5072), .I4(n5073), .O(n5074));
  LUT3 #(.INIT(8'h96)) lut_n5075 (.I0(n5061), .I1(n5064), .I2(n5065), .O(n5075));
  LUT3 #(.INIT(8'hE8)) lut_n5076 (.I0(n5071), .I1(n5074), .I2(n5075), .O(n5076));
  LUT3 #(.INIT(8'hE8)) lut_n5077 (.I0(x2532), .I1(x2533), .I2(x2534), .O(n5077));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5078 (.I0(x2523), .I1(x2524), .I2(x2525), .I3(n5072), .I4(n5073), .O(n5078));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5079 (.I0(x2529), .I1(x2530), .I2(x2531), .I3(n5077), .I4(n5078), .O(n5079));
  LUT3 #(.INIT(8'hE8)) lut_n5080 (.I0(x2538), .I1(x2539), .I2(x2540), .O(n5080));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5081 (.I0(x2529), .I1(x2530), .I2(x2531), .I3(n5077), .I4(n5078), .O(n5081));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5082 (.I0(x2535), .I1(x2536), .I2(x2537), .I3(n5080), .I4(n5081), .O(n5082));
  LUT3 #(.INIT(8'h96)) lut_n5083 (.I0(n5071), .I1(n5074), .I2(n5075), .O(n5083));
  LUT3 #(.INIT(8'hE8)) lut_n5084 (.I0(n5079), .I1(n5082), .I2(n5083), .O(n5084));
  LUT3 #(.INIT(8'h96)) lut_n5085 (.I0(n5058), .I1(n5066), .I2(n5067), .O(n5085));
  LUT3 #(.INIT(8'hE8)) lut_n5086 (.I0(n5076), .I1(n5084), .I2(n5085), .O(n5086));
  LUT3 #(.INIT(8'h96)) lut_n5087 (.I0(n5026), .I1(n5044), .I2(n5045), .O(n5087));
  LUT3 #(.INIT(8'hE8)) lut_n5088 (.I0(n5068), .I1(n5086), .I2(n5087), .O(n5088));
  LUT3 #(.INIT(8'hE8)) lut_n5089 (.I0(x2544), .I1(x2545), .I2(x2546), .O(n5089));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5090 (.I0(x2535), .I1(x2536), .I2(x2537), .I3(n5080), .I4(n5081), .O(n5090));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5091 (.I0(x2541), .I1(x2542), .I2(x2543), .I3(n5089), .I4(n5090), .O(n5091));
  LUT3 #(.INIT(8'hE8)) lut_n5092 (.I0(x2550), .I1(x2551), .I2(x2552), .O(n5092));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5093 (.I0(x2541), .I1(x2542), .I2(x2543), .I3(n5089), .I4(n5090), .O(n5093));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5094 (.I0(x2547), .I1(x2548), .I2(x2549), .I3(n5092), .I4(n5093), .O(n5094));
  LUT3 #(.INIT(8'h96)) lut_n5095 (.I0(n5079), .I1(n5082), .I2(n5083), .O(n5095));
  LUT3 #(.INIT(8'hE8)) lut_n5096 (.I0(n5091), .I1(n5094), .I2(n5095), .O(n5096));
  LUT3 #(.INIT(8'hE8)) lut_n5097 (.I0(x2556), .I1(x2557), .I2(x2558), .O(n5097));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5098 (.I0(x2547), .I1(x2548), .I2(x2549), .I3(n5092), .I4(n5093), .O(n5098));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5099 (.I0(x2553), .I1(x2554), .I2(x2555), .I3(n5097), .I4(n5098), .O(n5099));
  LUT3 #(.INIT(8'hE8)) lut_n5100 (.I0(x2562), .I1(x2563), .I2(x2564), .O(n5100));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5101 (.I0(x2553), .I1(x2554), .I2(x2555), .I3(n5097), .I4(n5098), .O(n5101));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5102 (.I0(x2559), .I1(x2560), .I2(x2561), .I3(n5100), .I4(n5101), .O(n5102));
  LUT3 #(.INIT(8'h96)) lut_n5103 (.I0(n5091), .I1(n5094), .I2(n5095), .O(n5103));
  LUT3 #(.INIT(8'hE8)) lut_n5104 (.I0(n5099), .I1(n5102), .I2(n5103), .O(n5104));
  LUT3 #(.INIT(8'h96)) lut_n5105 (.I0(n5076), .I1(n5084), .I2(n5085), .O(n5105));
  LUT3 #(.INIT(8'hE8)) lut_n5106 (.I0(n5096), .I1(n5104), .I2(n5105), .O(n5106));
  LUT3 #(.INIT(8'hE8)) lut_n5107 (.I0(x2568), .I1(x2569), .I2(x2570), .O(n5107));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5108 (.I0(x2559), .I1(x2560), .I2(x2561), .I3(n5100), .I4(n5101), .O(n5108));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5109 (.I0(x2565), .I1(x2566), .I2(x2567), .I3(n5107), .I4(n5108), .O(n5109));
  LUT3 #(.INIT(8'hE8)) lut_n5110 (.I0(x2574), .I1(x2575), .I2(x2576), .O(n5110));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5111 (.I0(x2565), .I1(x2566), .I2(x2567), .I3(n5107), .I4(n5108), .O(n5111));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5112 (.I0(x2571), .I1(x2572), .I2(x2573), .I3(n5110), .I4(n5111), .O(n5112));
  LUT3 #(.INIT(8'h96)) lut_n5113 (.I0(n5099), .I1(n5102), .I2(n5103), .O(n5113));
  LUT3 #(.INIT(8'hE8)) lut_n5114 (.I0(n5109), .I1(n5112), .I2(n5113), .O(n5114));
  LUT3 #(.INIT(8'hE8)) lut_n5115 (.I0(x2580), .I1(x2581), .I2(x2582), .O(n5115));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5116 (.I0(x2571), .I1(x2572), .I2(x2573), .I3(n5110), .I4(n5111), .O(n5116));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5117 (.I0(x2577), .I1(x2578), .I2(x2579), .I3(n5115), .I4(n5116), .O(n5117));
  LUT3 #(.INIT(8'hE8)) lut_n5118 (.I0(x2586), .I1(x2587), .I2(x2588), .O(n5118));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5119 (.I0(x2577), .I1(x2578), .I2(x2579), .I3(n5115), .I4(n5116), .O(n5119));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5120 (.I0(x2583), .I1(x2584), .I2(x2585), .I3(n5118), .I4(n5119), .O(n5120));
  LUT3 #(.INIT(8'h96)) lut_n5121 (.I0(n5109), .I1(n5112), .I2(n5113), .O(n5121));
  LUT3 #(.INIT(8'hE8)) lut_n5122 (.I0(n5117), .I1(n5120), .I2(n5121), .O(n5122));
  LUT3 #(.INIT(8'h96)) lut_n5123 (.I0(n5096), .I1(n5104), .I2(n5105), .O(n5123));
  LUT3 #(.INIT(8'hE8)) lut_n5124 (.I0(n5114), .I1(n5122), .I2(n5123), .O(n5124));
  LUT3 #(.INIT(8'h96)) lut_n5125 (.I0(n5068), .I1(n5086), .I2(n5087), .O(n5125));
  LUT3 #(.INIT(8'hE8)) lut_n5126 (.I0(n5106), .I1(n5124), .I2(n5125), .O(n5126));
  LUT3 #(.INIT(8'h96)) lut_n5127 (.I0(n5008), .I1(n5046), .I2(n5047), .O(n5127));
  LUT3 #(.INIT(8'hE8)) lut_n5128 (.I0(n5088), .I1(n5126), .I2(n5127), .O(n5128));
  LUT3 #(.INIT(8'hE8)) lut_n5129 (.I0(x2592), .I1(x2593), .I2(x2594), .O(n5129));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5130 (.I0(x2583), .I1(x2584), .I2(x2585), .I3(n5118), .I4(n5119), .O(n5130));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5131 (.I0(x2589), .I1(x2590), .I2(x2591), .I3(n5129), .I4(n5130), .O(n5131));
  LUT3 #(.INIT(8'hE8)) lut_n5132 (.I0(x2598), .I1(x2599), .I2(x2600), .O(n5132));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5133 (.I0(x2589), .I1(x2590), .I2(x2591), .I3(n5129), .I4(n5130), .O(n5133));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5134 (.I0(x2595), .I1(x2596), .I2(x2597), .I3(n5132), .I4(n5133), .O(n5134));
  LUT3 #(.INIT(8'h96)) lut_n5135 (.I0(n5117), .I1(n5120), .I2(n5121), .O(n5135));
  LUT3 #(.INIT(8'hE8)) lut_n5136 (.I0(n5131), .I1(n5134), .I2(n5135), .O(n5136));
  LUT3 #(.INIT(8'hE8)) lut_n5137 (.I0(x2604), .I1(x2605), .I2(x2606), .O(n5137));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5138 (.I0(x2595), .I1(x2596), .I2(x2597), .I3(n5132), .I4(n5133), .O(n5138));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5139 (.I0(x2601), .I1(x2602), .I2(x2603), .I3(n5137), .I4(n5138), .O(n5139));
  LUT3 #(.INIT(8'hE8)) lut_n5140 (.I0(x2610), .I1(x2611), .I2(x2612), .O(n5140));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5141 (.I0(x2601), .I1(x2602), .I2(x2603), .I3(n5137), .I4(n5138), .O(n5141));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5142 (.I0(x2607), .I1(x2608), .I2(x2609), .I3(n5140), .I4(n5141), .O(n5142));
  LUT3 #(.INIT(8'h96)) lut_n5143 (.I0(n5131), .I1(n5134), .I2(n5135), .O(n5143));
  LUT3 #(.INIT(8'hE8)) lut_n5144 (.I0(n5139), .I1(n5142), .I2(n5143), .O(n5144));
  LUT3 #(.INIT(8'h96)) lut_n5145 (.I0(n5114), .I1(n5122), .I2(n5123), .O(n5145));
  LUT3 #(.INIT(8'hE8)) lut_n5146 (.I0(n5136), .I1(n5144), .I2(n5145), .O(n5146));
  LUT3 #(.INIT(8'hE8)) lut_n5147 (.I0(x2616), .I1(x2617), .I2(x2618), .O(n5147));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5148 (.I0(x2607), .I1(x2608), .I2(x2609), .I3(n5140), .I4(n5141), .O(n5148));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5149 (.I0(x2613), .I1(x2614), .I2(x2615), .I3(n5147), .I4(n5148), .O(n5149));
  LUT3 #(.INIT(8'hE8)) lut_n5150 (.I0(x2622), .I1(x2623), .I2(x2624), .O(n5150));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5151 (.I0(x2613), .I1(x2614), .I2(x2615), .I3(n5147), .I4(n5148), .O(n5151));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5152 (.I0(x2619), .I1(x2620), .I2(x2621), .I3(n5150), .I4(n5151), .O(n5152));
  LUT3 #(.INIT(8'h96)) lut_n5153 (.I0(n5139), .I1(n5142), .I2(n5143), .O(n5153));
  LUT3 #(.INIT(8'hE8)) lut_n5154 (.I0(n5149), .I1(n5152), .I2(n5153), .O(n5154));
  LUT3 #(.INIT(8'hE8)) lut_n5155 (.I0(x2628), .I1(x2629), .I2(x2630), .O(n5155));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5156 (.I0(x2619), .I1(x2620), .I2(x2621), .I3(n5150), .I4(n5151), .O(n5156));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5157 (.I0(x2625), .I1(x2626), .I2(x2627), .I3(n5155), .I4(n5156), .O(n5157));
  LUT3 #(.INIT(8'hE8)) lut_n5158 (.I0(x2634), .I1(x2635), .I2(x2636), .O(n5158));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5159 (.I0(x2625), .I1(x2626), .I2(x2627), .I3(n5155), .I4(n5156), .O(n5159));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5160 (.I0(x2631), .I1(x2632), .I2(x2633), .I3(n5158), .I4(n5159), .O(n5160));
  LUT3 #(.INIT(8'h96)) lut_n5161 (.I0(n5149), .I1(n5152), .I2(n5153), .O(n5161));
  LUT3 #(.INIT(8'hE8)) lut_n5162 (.I0(n5157), .I1(n5160), .I2(n5161), .O(n5162));
  LUT3 #(.INIT(8'h96)) lut_n5163 (.I0(n5136), .I1(n5144), .I2(n5145), .O(n5163));
  LUT3 #(.INIT(8'hE8)) lut_n5164 (.I0(n5154), .I1(n5162), .I2(n5163), .O(n5164));
  LUT3 #(.INIT(8'h96)) lut_n5165 (.I0(n5106), .I1(n5124), .I2(n5125), .O(n5165));
  LUT3 #(.INIT(8'hE8)) lut_n5166 (.I0(n5146), .I1(n5164), .I2(n5165), .O(n5166));
  LUT3 #(.INIT(8'hE8)) lut_n5167 (.I0(x2640), .I1(x2641), .I2(x2642), .O(n5167));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5168 (.I0(x2631), .I1(x2632), .I2(x2633), .I3(n5158), .I4(n5159), .O(n5168));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5169 (.I0(x2637), .I1(x2638), .I2(x2639), .I3(n5167), .I4(n5168), .O(n5169));
  LUT3 #(.INIT(8'hE8)) lut_n5170 (.I0(x2646), .I1(x2647), .I2(x2648), .O(n5170));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5171 (.I0(x2637), .I1(x2638), .I2(x2639), .I3(n5167), .I4(n5168), .O(n5171));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5172 (.I0(x2643), .I1(x2644), .I2(x2645), .I3(n5170), .I4(n5171), .O(n5172));
  LUT3 #(.INIT(8'h96)) lut_n5173 (.I0(n5157), .I1(n5160), .I2(n5161), .O(n5173));
  LUT3 #(.INIT(8'hE8)) lut_n5174 (.I0(n5169), .I1(n5172), .I2(n5173), .O(n5174));
  LUT3 #(.INIT(8'hE8)) lut_n5175 (.I0(x2652), .I1(x2653), .I2(x2654), .O(n5175));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5176 (.I0(x2643), .I1(x2644), .I2(x2645), .I3(n5170), .I4(n5171), .O(n5176));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5177 (.I0(x2649), .I1(x2650), .I2(x2651), .I3(n5175), .I4(n5176), .O(n5177));
  LUT3 #(.INIT(8'hE8)) lut_n5178 (.I0(x2658), .I1(x2659), .I2(x2660), .O(n5178));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5179 (.I0(x2649), .I1(x2650), .I2(x2651), .I3(n5175), .I4(n5176), .O(n5179));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5180 (.I0(x2655), .I1(x2656), .I2(x2657), .I3(n5178), .I4(n5179), .O(n5180));
  LUT3 #(.INIT(8'h96)) lut_n5181 (.I0(n5169), .I1(n5172), .I2(n5173), .O(n5181));
  LUT3 #(.INIT(8'hE8)) lut_n5182 (.I0(n5177), .I1(n5180), .I2(n5181), .O(n5182));
  LUT3 #(.INIT(8'h96)) lut_n5183 (.I0(n5154), .I1(n5162), .I2(n5163), .O(n5183));
  LUT3 #(.INIT(8'hE8)) lut_n5184 (.I0(n5174), .I1(n5182), .I2(n5183), .O(n5184));
  LUT3 #(.INIT(8'hE8)) lut_n5185 (.I0(x2664), .I1(x2665), .I2(x2666), .O(n5185));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5186 (.I0(x2655), .I1(x2656), .I2(x2657), .I3(n5178), .I4(n5179), .O(n5186));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5187 (.I0(x2661), .I1(x2662), .I2(x2663), .I3(n5185), .I4(n5186), .O(n5187));
  LUT3 #(.INIT(8'hE8)) lut_n5188 (.I0(x2670), .I1(x2671), .I2(x2672), .O(n5188));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5189 (.I0(x2661), .I1(x2662), .I2(x2663), .I3(n5185), .I4(n5186), .O(n5189));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5190 (.I0(x2667), .I1(x2668), .I2(x2669), .I3(n5188), .I4(n5189), .O(n5190));
  LUT3 #(.INIT(8'h96)) lut_n5191 (.I0(n5177), .I1(n5180), .I2(n5181), .O(n5191));
  LUT3 #(.INIT(8'hE8)) lut_n5192 (.I0(n5187), .I1(n5190), .I2(n5191), .O(n5192));
  LUT3 #(.INIT(8'hE8)) lut_n5193 (.I0(x2676), .I1(x2677), .I2(x2678), .O(n5193));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5194 (.I0(x2667), .I1(x2668), .I2(x2669), .I3(n5188), .I4(n5189), .O(n5194));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5195 (.I0(x2673), .I1(x2674), .I2(x2675), .I3(n5193), .I4(n5194), .O(n5195));
  LUT3 #(.INIT(8'hE8)) lut_n5196 (.I0(x2682), .I1(x2683), .I2(x2684), .O(n5196));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5197 (.I0(x2673), .I1(x2674), .I2(x2675), .I3(n5193), .I4(n5194), .O(n5197));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5198 (.I0(x2679), .I1(x2680), .I2(x2681), .I3(n5196), .I4(n5197), .O(n5198));
  LUT3 #(.INIT(8'h96)) lut_n5199 (.I0(n5187), .I1(n5190), .I2(n5191), .O(n5199));
  LUT3 #(.INIT(8'hE8)) lut_n5200 (.I0(n5195), .I1(n5198), .I2(n5199), .O(n5200));
  LUT3 #(.INIT(8'h96)) lut_n5201 (.I0(n5174), .I1(n5182), .I2(n5183), .O(n5201));
  LUT3 #(.INIT(8'hE8)) lut_n5202 (.I0(n5192), .I1(n5200), .I2(n5201), .O(n5202));
  LUT3 #(.INIT(8'h96)) lut_n5203 (.I0(n5146), .I1(n5164), .I2(n5165), .O(n5203));
  LUT3 #(.INIT(8'hE8)) lut_n5204 (.I0(n5184), .I1(n5202), .I2(n5203), .O(n5204));
  LUT3 #(.INIT(8'h96)) lut_n5205 (.I0(n5088), .I1(n5126), .I2(n5127), .O(n5205));
  LUT3 #(.INIT(8'hE8)) lut_n5206 (.I0(n5166), .I1(n5204), .I2(n5205), .O(n5206));
  LUT3 #(.INIT(8'h96)) lut_n5207 (.I0(n4970), .I1(n5048), .I2(n5049), .O(n5207));
  LUT3 #(.INIT(8'hE8)) lut_n5208 (.I0(n5128), .I1(n5206), .I2(n5207), .O(n5208));
  LUT3 #(.INIT(8'h96)) lut_n5209 (.I0(n4730), .I1(n4888), .I2(n4889), .O(n5209));
  LUT3 #(.INIT(8'hE8)) lut_n5210 (.I0(n5050), .I1(n5208), .I2(n5209), .O(n5210));
  LUT3 #(.INIT(8'hE8)) lut_n5211 (.I0(x2688), .I1(x2689), .I2(x2690), .O(n5211));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5212 (.I0(x2679), .I1(x2680), .I2(x2681), .I3(n5196), .I4(n5197), .O(n5212));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5213 (.I0(x2685), .I1(x2686), .I2(x2687), .I3(n5211), .I4(n5212), .O(n5213));
  LUT3 #(.INIT(8'hE8)) lut_n5214 (.I0(x2694), .I1(x2695), .I2(x2696), .O(n5214));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5215 (.I0(x2685), .I1(x2686), .I2(x2687), .I3(n5211), .I4(n5212), .O(n5215));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5216 (.I0(x2691), .I1(x2692), .I2(x2693), .I3(n5214), .I4(n5215), .O(n5216));
  LUT3 #(.INIT(8'h96)) lut_n5217 (.I0(n5195), .I1(n5198), .I2(n5199), .O(n5217));
  LUT3 #(.INIT(8'hE8)) lut_n5218 (.I0(n5213), .I1(n5216), .I2(n5217), .O(n5218));
  LUT3 #(.INIT(8'hE8)) lut_n5219 (.I0(x2700), .I1(x2701), .I2(x2702), .O(n5219));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5220 (.I0(x2691), .I1(x2692), .I2(x2693), .I3(n5214), .I4(n5215), .O(n5220));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5221 (.I0(x2697), .I1(x2698), .I2(x2699), .I3(n5219), .I4(n5220), .O(n5221));
  LUT3 #(.INIT(8'hE8)) lut_n5222 (.I0(x2706), .I1(x2707), .I2(x2708), .O(n5222));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5223 (.I0(x2697), .I1(x2698), .I2(x2699), .I3(n5219), .I4(n5220), .O(n5223));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5224 (.I0(x2703), .I1(x2704), .I2(x2705), .I3(n5222), .I4(n5223), .O(n5224));
  LUT3 #(.INIT(8'h96)) lut_n5225 (.I0(n5213), .I1(n5216), .I2(n5217), .O(n5225));
  LUT3 #(.INIT(8'hE8)) lut_n5226 (.I0(n5221), .I1(n5224), .I2(n5225), .O(n5226));
  LUT3 #(.INIT(8'h96)) lut_n5227 (.I0(n5192), .I1(n5200), .I2(n5201), .O(n5227));
  LUT3 #(.INIT(8'hE8)) lut_n5228 (.I0(n5218), .I1(n5226), .I2(n5227), .O(n5228));
  LUT3 #(.INIT(8'hE8)) lut_n5229 (.I0(x2712), .I1(x2713), .I2(x2714), .O(n5229));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5230 (.I0(x2703), .I1(x2704), .I2(x2705), .I3(n5222), .I4(n5223), .O(n5230));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5231 (.I0(x2709), .I1(x2710), .I2(x2711), .I3(n5229), .I4(n5230), .O(n5231));
  LUT3 #(.INIT(8'hE8)) lut_n5232 (.I0(x2718), .I1(x2719), .I2(x2720), .O(n5232));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5233 (.I0(x2709), .I1(x2710), .I2(x2711), .I3(n5229), .I4(n5230), .O(n5233));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5234 (.I0(x2715), .I1(x2716), .I2(x2717), .I3(n5232), .I4(n5233), .O(n5234));
  LUT3 #(.INIT(8'h96)) lut_n5235 (.I0(n5221), .I1(n5224), .I2(n5225), .O(n5235));
  LUT3 #(.INIT(8'hE8)) lut_n5236 (.I0(n5231), .I1(n5234), .I2(n5235), .O(n5236));
  LUT3 #(.INIT(8'hE8)) lut_n5237 (.I0(x2724), .I1(x2725), .I2(x2726), .O(n5237));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5238 (.I0(x2715), .I1(x2716), .I2(x2717), .I3(n5232), .I4(n5233), .O(n5238));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5239 (.I0(x2721), .I1(x2722), .I2(x2723), .I3(n5237), .I4(n5238), .O(n5239));
  LUT3 #(.INIT(8'hE8)) lut_n5240 (.I0(x2730), .I1(x2731), .I2(x2732), .O(n5240));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5241 (.I0(x2721), .I1(x2722), .I2(x2723), .I3(n5237), .I4(n5238), .O(n5241));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5242 (.I0(x2727), .I1(x2728), .I2(x2729), .I3(n5240), .I4(n5241), .O(n5242));
  LUT3 #(.INIT(8'h96)) lut_n5243 (.I0(n5231), .I1(n5234), .I2(n5235), .O(n5243));
  LUT3 #(.INIT(8'hE8)) lut_n5244 (.I0(n5239), .I1(n5242), .I2(n5243), .O(n5244));
  LUT3 #(.INIT(8'h96)) lut_n5245 (.I0(n5218), .I1(n5226), .I2(n5227), .O(n5245));
  LUT3 #(.INIT(8'hE8)) lut_n5246 (.I0(n5236), .I1(n5244), .I2(n5245), .O(n5246));
  LUT3 #(.INIT(8'h96)) lut_n5247 (.I0(n5184), .I1(n5202), .I2(n5203), .O(n5247));
  LUT3 #(.INIT(8'hE8)) lut_n5248 (.I0(n5228), .I1(n5246), .I2(n5247), .O(n5248));
  LUT3 #(.INIT(8'hE8)) lut_n5249 (.I0(x2736), .I1(x2737), .I2(x2738), .O(n5249));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5250 (.I0(x2727), .I1(x2728), .I2(x2729), .I3(n5240), .I4(n5241), .O(n5250));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5251 (.I0(x2733), .I1(x2734), .I2(x2735), .I3(n5249), .I4(n5250), .O(n5251));
  LUT3 #(.INIT(8'hE8)) lut_n5252 (.I0(x2742), .I1(x2743), .I2(x2744), .O(n5252));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5253 (.I0(x2733), .I1(x2734), .I2(x2735), .I3(n5249), .I4(n5250), .O(n5253));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5254 (.I0(x2739), .I1(x2740), .I2(x2741), .I3(n5252), .I4(n5253), .O(n5254));
  LUT3 #(.INIT(8'h96)) lut_n5255 (.I0(n5239), .I1(n5242), .I2(n5243), .O(n5255));
  LUT3 #(.INIT(8'hE8)) lut_n5256 (.I0(n5251), .I1(n5254), .I2(n5255), .O(n5256));
  LUT3 #(.INIT(8'hE8)) lut_n5257 (.I0(x2748), .I1(x2749), .I2(x2750), .O(n5257));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5258 (.I0(x2739), .I1(x2740), .I2(x2741), .I3(n5252), .I4(n5253), .O(n5258));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5259 (.I0(x2745), .I1(x2746), .I2(x2747), .I3(n5257), .I4(n5258), .O(n5259));
  LUT3 #(.INIT(8'hE8)) lut_n5260 (.I0(x2754), .I1(x2755), .I2(x2756), .O(n5260));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5261 (.I0(x2745), .I1(x2746), .I2(x2747), .I3(n5257), .I4(n5258), .O(n5261));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5262 (.I0(x2751), .I1(x2752), .I2(x2753), .I3(n5260), .I4(n5261), .O(n5262));
  LUT3 #(.INIT(8'h96)) lut_n5263 (.I0(n5251), .I1(n5254), .I2(n5255), .O(n5263));
  LUT3 #(.INIT(8'hE8)) lut_n5264 (.I0(n5259), .I1(n5262), .I2(n5263), .O(n5264));
  LUT3 #(.INIT(8'h96)) lut_n5265 (.I0(n5236), .I1(n5244), .I2(n5245), .O(n5265));
  LUT3 #(.INIT(8'hE8)) lut_n5266 (.I0(n5256), .I1(n5264), .I2(n5265), .O(n5266));
  LUT3 #(.INIT(8'hE8)) lut_n5267 (.I0(x2760), .I1(x2761), .I2(x2762), .O(n5267));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5268 (.I0(x2751), .I1(x2752), .I2(x2753), .I3(n5260), .I4(n5261), .O(n5268));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5269 (.I0(x2757), .I1(x2758), .I2(x2759), .I3(n5267), .I4(n5268), .O(n5269));
  LUT3 #(.INIT(8'hE8)) lut_n5270 (.I0(x2766), .I1(x2767), .I2(x2768), .O(n5270));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5271 (.I0(x2757), .I1(x2758), .I2(x2759), .I3(n5267), .I4(n5268), .O(n5271));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5272 (.I0(x2763), .I1(x2764), .I2(x2765), .I3(n5270), .I4(n5271), .O(n5272));
  LUT3 #(.INIT(8'h96)) lut_n5273 (.I0(n5259), .I1(n5262), .I2(n5263), .O(n5273));
  LUT3 #(.INIT(8'hE8)) lut_n5274 (.I0(n5269), .I1(n5272), .I2(n5273), .O(n5274));
  LUT3 #(.INIT(8'hE8)) lut_n5275 (.I0(x2772), .I1(x2773), .I2(x2774), .O(n5275));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5276 (.I0(x2763), .I1(x2764), .I2(x2765), .I3(n5270), .I4(n5271), .O(n5276));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5277 (.I0(x2769), .I1(x2770), .I2(x2771), .I3(n5275), .I4(n5276), .O(n5277));
  LUT3 #(.INIT(8'hE8)) lut_n5278 (.I0(x2778), .I1(x2779), .I2(x2780), .O(n5278));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5279 (.I0(x2769), .I1(x2770), .I2(x2771), .I3(n5275), .I4(n5276), .O(n5279));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5280 (.I0(x2775), .I1(x2776), .I2(x2777), .I3(n5278), .I4(n5279), .O(n5280));
  LUT3 #(.INIT(8'h96)) lut_n5281 (.I0(n5269), .I1(n5272), .I2(n5273), .O(n5281));
  LUT3 #(.INIT(8'hE8)) lut_n5282 (.I0(n5277), .I1(n5280), .I2(n5281), .O(n5282));
  LUT3 #(.INIT(8'h96)) lut_n5283 (.I0(n5256), .I1(n5264), .I2(n5265), .O(n5283));
  LUT3 #(.INIT(8'hE8)) lut_n5284 (.I0(n5274), .I1(n5282), .I2(n5283), .O(n5284));
  LUT3 #(.INIT(8'h96)) lut_n5285 (.I0(n5228), .I1(n5246), .I2(n5247), .O(n5285));
  LUT3 #(.INIT(8'hE8)) lut_n5286 (.I0(n5266), .I1(n5284), .I2(n5285), .O(n5286));
  LUT3 #(.INIT(8'h96)) lut_n5287 (.I0(n5166), .I1(n5204), .I2(n5205), .O(n5287));
  LUT3 #(.INIT(8'hE8)) lut_n5288 (.I0(n5248), .I1(n5286), .I2(n5287), .O(n5288));
  LUT3 #(.INIT(8'hE8)) lut_n5289 (.I0(x2784), .I1(x2785), .I2(x2786), .O(n5289));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5290 (.I0(x2775), .I1(x2776), .I2(x2777), .I3(n5278), .I4(n5279), .O(n5290));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5291 (.I0(x2781), .I1(x2782), .I2(x2783), .I3(n5289), .I4(n5290), .O(n5291));
  LUT3 #(.INIT(8'hE8)) lut_n5292 (.I0(x2790), .I1(x2791), .I2(x2792), .O(n5292));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5293 (.I0(x2781), .I1(x2782), .I2(x2783), .I3(n5289), .I4(n5290), .O(n5293));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5294 (.I0(x2787), .I1(x2788), .I2(x2789), .I3(n5292), .I4(n5293), .O(n5294));
  LUT3 #(.INIT(8'h96)) lut_n5295 (.I0(n5277), .I1(n5280), .I2(n5281), .O(n5295));
  LUT3 #(.INIT(8'hE8)) lut_n5296 (.I0(n5291), .I1(n5294), .I2(n5295), .O(n5296));
  LUT3 #(.INIT(8'hE8)) lut_n5297 (.I0(x2796), .I1(x2797), .I2(x2798), .O(n5297));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5298 (.I0(x2787), .I1(x2788), .I2(x2789), .I3(n5292), .I4(n5293), .O(n5298));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5299 (.I0(x2793), .I1(x2794), .I2(x2795), .I3(n5297), .I4(n5298), .O(n5299));
  LUT3 #(.INIT(8'hE8)) lut_n5300 (.I0(x2802), .I1(x2803), .I2(x2804), .O(n5300));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5301 (.I0(x2793), .I1(x2794), .I2(x2795), .I3(n5297), .I4(n5298), .O(n5301));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5302 (.I0(x2799), .I1(x2800), .I2(x2801), .I3(n5300), .I4(n5301), .O(n5302));
  LUT3 #(.INIT(8'h96)) lut_n5303 (.I0(n5291), .I1(n5294), .I2(n5295), .O(n5303));
  LUT3 #(.INIT(8'hE8)) lut_n5304 (.I0(n5299), .I1(n5302), .I2(n5303), .O(n5304));
  LUT3 #(.INIT(8'h96)) lut_n5305 (.I0(n5274), .I1(n5282), .I2(n5283), .O(n5305));
  LUT3 #(.INIT(8'hE8)) lut_n5306 (.I0(n5296), .I1(n5304), .I2(n5305), .O(n5306));
  LUT3 #(.INIT(8'hE8)) lut_n5307 (.I0(x2808), .I1(x2809), .I2(x2810), .O(n5307));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5308 (.I0(x2799), .I1(x2800), .I2(x2801), .I3(n5300), .I4(n5301), .O(n5308));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5309 (.I0(x2805), .I1(x2806), .I2(x2807), .I3(n5307), .I4(n5308), .O(n5309));
  LUT3 #(.INIT(8'hE8)) lut_n5310 (.I0(x2814), .I1(x2815), .I2(x2816), .O(n5310));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5311 (.I0(x2805), .I1(x2806), .I2(x2807), .I3(n5307), .I4(n5308), .O(n5311));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5312 (.I0(x2811), .I1(x2812), .I2(x2813), .I3(n5310), .I4(n5311), .O(n5312));
  LUT3 #(.INIT(8'h96)) lut_n5313 (.I0(n5299), .I1(n5302), .I2(n5303), .O(n5313));
  LUT3 #(.INIT(8'hE8)) lut_n5314 (.I0(n5309), .I1(n5312), .I2(n5313), .O(n5314));
  LUT3 #(.INIT(8'hE8)) lut_n5315 (.I0(x2820), .I1(x2821), .I2(x2822), .O(n5315));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5316 (.I0(x2811), .I1(x2812), .I2(x2813), .I3(n5310), .I4(n5311), .O(n5316));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5317 (.I0(x2817), .I1(x2818), .I2(x2819), .I3(n5315), .I4(n5316), .O(n5317));
  LUT3 #(.INIT(8'hE8)) lut_n5318 (.I0(x2826), .I1(x2827), .I2(x2828), .O(n5318));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5319 (.I0(x2817), .I1(x2818), .I2(x2819), .I3(n5315), .I4(n5316), .O(n5319));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5320 (.I0(x2823), .I1(x2824), .I2(x2825), .I3(n5318), .I4(n5319), .O(n5320));
  LUT3 #(.INIT(8'h96)) lut_n5321 (.I0(n5309), .I1(n5312), .I2(n5313), .O(n5321));
  LUT3 #(.INIT(8'hE8)) lut_n5322 (.I0(n5317), .I1(n5320), .I2(n5321), .O(n5322));
  LUT3 #(.INIT(8'h96)) lut_n5323 (.I0(n5296), .I1(n5304), .I2(n5305), .O(n5323));
  LUT3 #(.INIT(8'hE8)) lut_n5324 (.I0(n5314), .I1(n5322), .I2(n5323), .O(n5324));
  LUT3 #(.INIT(8'h96)) lut_n5325 (.I0(n5266), .I1(n5284), .I2(n5285), .O(n5325));
  LUT3 #(.INIT(8'hE8)) lut_n5326 (.I0(n5306), .I1(n5324), .I2(n5325), .O(n5326));
  LUT3 #(.INIT(8'hE8)) lut_n5327 (.I0(x2832), .I1(x2833), .I2(x2834), .O(n5327));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5328 (.I0(x2823), .I1(x2824), .I2(x2825), .I3(n5318), .I4(n5319), .O(n5328));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5329 (.I0(x2829), .I1(x2830), .I2(x2831), .I3(n5327), .I4(n5328), .O(n5329));
  LUT3 #(.INIT(8'hE8)) lut_n5330 (.I0(x2838), .I1(x2839), .I2(x2840), .O(n5330));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5331 (.I0(x2829), .I1(x2830), .I2(x2831), .I3(n5327), .I4(n5328), .O(n5331));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5332 (.I0(x2835), .I1(x2836), .I2(x2837), .I3(n5330), .I4(n5331), .O(n5332));
  LUT3 #(.INIT(8'h96)) lut_n5333 (.I0(n5317), .I1(n5320), .I2(n5321), .O(n5333));
  LUT3 #(.INIT(8'hE8)) lut_n5334 (.I0(n5329), .I1(n5332), .I2(n5333), .O(n5334));
  LUT3 #(.INIT(8'hE8)) lut_n5335 (.I0(x2844), .I1(x2845), .I2(x2846), .O(n5335));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5336 (.I0(x2835), .I1(x2836), .I2(x2837), .I3(n5330), .I4(n5331), .O(n5336));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5337 (.I0(x2841), .I1(x2842), .I2(x2843), .I3(n5335), .I4(n5336), .O(n5337));
  LUT3 #(.INIT(8'hE8)) lut_n5338 (.I0(x2850), .I1(x2851), .I2(x2852), .O(n5338));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5339 (.I0(x2841), .I1(x2842), .I2(x2843), .I3(n5335), .I4(n5336), .O(n5339));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5340 (.I0(x2847), .I1(x2848), .I2(x2849), .I3(n5338), .I4(n5339), .O(n5340));
  LUT3 #(.INIT(8'h96)) lut_n5341 (.I0(n5329), .I1(n5332), .I2(n5333), .O(n5341));
  LUT3 #(.INIT(8'hE8)) lut_n5342 (.I0(n5337), .I1(n5340), .I2(n5341), .O(n5342));
  LUT3 #(.INIT(8'h96)) lut_n5343 (.I0(n5314), .I1(n5322), .I2(n5323), .O(n5343));
  LUT3 #(.INIT(8'hE8)) lut_n5344 (.I0(n5334), .I1(n5342), .I2(n5343), .O(n5344));
  LUT3 #(.INIT(8'hE8)) lut_n5345 (.I0(x2856), .I1(x2857), .I2(x2858), .O(n5345));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5346 (.I0(x2847), .I1(x2848), .I2(x2849), .I3(n5338), .I4(n5339), .O(n5346));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5347 (.I0(x2853), .I1(x2854), .I2(x2855), .I3(n5345), .I4(n5346), .O(n5347));
  LUT3 #(.INIT(8'hE8)) lut_n5348 (.I0(x2862), .I1(x2863), .I2(x2864), .O(n5348));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5349 (.I0(x2853), .I1(x2854), .I2(x2855), .I3(n5345), .I4(n5346), .O(n5349));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5350 (.I0(x2859), .I1(x2860), .I2(x2861), .I3(n5348), .I4(n5349), .O(n5350));
  LUT3 #(.INIT(8'h96)) lut_n5351 (.I0(n5337), .I1(n5340), .I2(n5341), .O(n5351));
  LUT3 #(.INIT(8'hE8)) lut_n5352 (.I0(n5347), .I1(n5350), .I2(n5351), .O(n5352));
  LUT3 #(.INIT(8'hE8)) lut_n5353 (.I0(x2868), .I1(x2869), .I2(x2870), .O(n5353));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5354 (.I0(x2859), .I1(x2860), .I2(x2861), .I3(n5348), .I4(n5349), .O(n5354));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5355 (.I0(x2865), .I1(x2866), .I2(x2867), .I3(n5353), .I4(n5354), .O(n5355));
  LUT3 #(.INIT(8'hE8)) lut_n5356 (.I0(x2874), .I1(x2875), .I2(x2876), .O(n5356));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5357 (.I0(x2865), .I1(x2866), .I2(x2867), .I3(n5353), .I4(n5354), .O(n5357));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5358 (.I0(x2871), .I1(x2872), .I2(x2873), .I3(n5356), .I4(n5357), .O(n5358));
  LUT3 #(.INIT(8'h96)) lut_n5359 (.I0(n5347), .I1(n5350), .I2(n5351), .O(n5359));
  LUT3 #(.INIT(8'hE8)) lut_n5360 (.I0(n5355), .I1(n5358), .I2(n5359), .O(n5360));
  LUT3 #(.INIT(8'h96)) lut_n5361 (.I0(n5334), .I1(n5342), .I2(n5343), .O(n5361));
  LUT3 #(.INIT(8'hE8)) lut_n5362 (.I0(n5352), .I1(n5360), .I2(n5361), .O(n5362));
  LUT3 #(.INIT(8'h96)) lut_n5363 (.I0(n5306), .I1(n5324), .I2(n5325), .O(n5363));
  LUT3 #(.INIT(8'hE8)) lut_n5364 (.I0(n5344), .I1(n5362), .I2(n5363), .O(n5364));
  LUT3 #(.INIT(8'h96)) lut_n5365 (.I0(n5248), .I1(n5286), .I2(n5287), .O(n5365));
  LUT3 #(.INIT(8'hE8)) lut_n5366 (.I0(n5326), .I1(n5364), .I2(n5365), .O(n5366));
  LUT3 #(.INIT(8'h96)) lut_n5367 (.I0(n5128), .I1(n5206), .I2(n5207), .O(n5367));
  LUT3 #(.INIT(8'hE8)) lut_n5368 (.I0(n5288), .I1(n5366), .I2(n5367), .O(n5368));
  LUT3 #(.INIT(8'hE8)) lut_n5369 (.I0(x2880), .I1(x2881), .I2(x2882), .O(n5369));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5370 (.I0(x2871), .I1(x2872), .I2(x2873), .I3(n5356), .I4(n5357), .O(n5370));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5371 (.I0(x2877), .I1(x2878), .I2(x2879), .I3(n5369), .I4(n5370), .O(n5371));
  LUT3 #(.INIT(8'hE8)) lut_n5372 (.I0(x2886), .I1(x2887), .I2(x2888), .O(n5372));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5373 (.I0(x2877), .I1(x2878), .I2(x2879), .I3(n5369), .I4(n5370), .O(n5373));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5374 (.I0(x2883), .I1(x2884), .I2(x2885), .I3(n5372), .I4(n5373), .O(n5374));
  LUT3 #(.INIT(8'h96)) lut_n5375 (.I0(n5355), .I1(n5358), .I2(n5359), .O(n5375));
  LUT3 #(.INIT(8'hE8)) lut_n5376 (.I0(n5371), .I1(n5374), .I2(n5375), .O(n5376));
  LUT3 #(.INIT(8'hE8)) lut_n5377 (.I0(x2892), .I1(x2893), .I2(x2894), .O(n5377));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5378 (.I0(x2883), .I1(x2884), .I2(x2885), .I3(n5372), .I4(n5373), .O(n5378));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5379 (.I0(x2889), .I1(x2890), .I2(x2891), .I3(n5377), .I4(n5378), .O(n5379));
  LUT3 #(.INIT(8'hE8)) lut_n5380 (.I0(x2898), .I1(x2899), .I2(x2900), .O(n5380));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5381 (.I0(x2889), .I1(x2890), .I2(x2891), .I3(n5377), .I4(n5378), .O(n5381));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5382 (.I0(x2895), .I1(x2896), .I2(x2897), .I3(n5380), .I4(n5381), .O(n5382));
  LUT3 #(.INIT(8'h96)) lut_n5383 (.I0(n5371), .I1(n5374), .I2(n5375), .O(n5383));
  LUT3 #(.INIT(8'hE8)) lut_n5384 (.I0(n5379), .I1(n5382), .I2(n5383), .O(n5384));
  LUT3 #(.INIT(8'h96)) lut_n5385 (.I0(n5352), .I1(n5360), .I2(n5361), .O(n5385));
  LUT3 #(.INIT(8'hE8)) lut_n5386 (.I0(n5376), .I1(n5384), .I2(n5385), .O(n5386));
  LUT3 #(.INIT(8'hE8)) lut_n5387 (.I0(x2904), .I1(x2905), .I2(x2906), .O(n5387));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5388 (.I0(x2895), .I1(x2896), .I2(x2897), .I3(n5380), .I4(n5381), .O(n5388));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5389 (.I0(x2901), .I1(x2902), .I2(x2903), .I3(n5387), .I4(n5388), .O(n5389));
  LUT3 #(.INIT(8'hE8)) lut_n5390 (.I0(x2910), .I1(x2911), .I2(x2912), .O(n5390));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5391 (.I0(x2901), .I1(x2902), .I2(x2903), .I3(n5387), .I4(n5388), .O(n5391));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5392 (.I0(x2907), .I1(x2908), .I2(x2909), .I3(n5390), .I4(n5391), .O(n5392));
  LUT3 #(.INIT(8'h96)) lut_n5393 (.I0(n5379), .I1(n5382), .I2(n5383), .O(n5393));
  LUT3 #(.INIT(8'hE8)) lut_n5394 (.I0(n5389), .I1(n5392), .I2(n5393), .O(n5394));
  LUT3 #(.INIT(8'hE8)) lut_n5395 (.I0(x2916), .I1(x2917), .I2(x2918), .O(n5395));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5396 (.I0(x2907), .I1(x2908), .I2(x2909), .I3(n5390), .I4(n5391), .O(n5396));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5397 (.I0(x2913), .I1(x2914), .I2(x2915), .I3(n5395), .I4(n5396), .O(n5397));
  LUT3 #(.INIT(8'hE8)) lut_n5398 (.I0(x2922), .I1(x2923), .I2(x2924), .O(n5398));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5399 (.I0(x2913), .I1(x2914), .I2(x2915), .I3(n5395), .I4(n5396), .O(n5399));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5400 (.I0(x2919), .I1(x2920), .I2(x2921), .I3(n5398), .I4(n5399), .O(n5400));
  LUT3 #(.INIT(8'h96)) lut_n5401 (.I0(n5389), .I1(n5392), .I2(n5393), .O(n5401));
  LUT3 #(.INIT(8'hE8)) lut_n5402 (.I0(n5397), .I1(n5400), .I2(n5401), .O(n5402));
  LUT3 #(.INIT(8'h96)) lut_n5403 (.I0(n5376), .I1(n5384), .I2(n5385), .O(n5403));
  LUT3 #(.INIT(8'hE8)) lut_n5404 (.I0(n5394), .I1(n5402), .I2(n5403), .O(n5404));
  LUT3 #(.INIT(8'h96)) lut_n5405 (.I0(n5344), .I1(n5362), .I2(n5363), .O(n5405));
  LUT3 #(.INIT(8'hE8)) lut_n5406 (.I0(n5386), .I1(n5404), .I2(n5405), .O(n5406));
  LUT3 #(.INIT(8'hE8)) lut_n5407 (.I0(x2928), .I1(x2929), .I2(x2930), .O(n5407));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5408 (.I0(x2919), .I1(x2920), .I2(x2921), .I3(n5398), .I4(n5399), .O(n5408));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5409 (.I0(x2925), .I1(x2926), .I2(x2927), .I3(n5407), .I4(n5408), .O(n5409));
  LUT3 #(.INIT(8'hE8)) lut_n5410 (.I0(x2934), .I1(x2935), .I2(x2936), .O(n5410));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5411 (.I0(x2925), .I1(x2926), .I2(x2927), .I3(n5407), .I4(n5408), .O(n5411));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5412 (.I0(x2931), .I1(x2932), .I2(x2933), .I3(n5410), .I4(n5411), .O(n5412));
  LUT3 #(.INIT(8'h96)) lut_n5413 (.I0(n5397), .I1(n5400), .I2(n5401), .O(n5413));
  LUT3 #(.INIT(8'hE8)) lut_n5414 (.I0(n5409), .I1(n5412), .I2(n5413), .O(n5414));
  LUT3 #(.INIT(8'hE8)) lut_n5415 (.I0(x2940), .I1(x2941), .I2(x2942), .O(n5415));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5416 (.I0(x2931), .I1(x2932), .I2(x2933), .I3(n5410), .I4(n5411), .O(n5416));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5417 (.I0(x2937), .I1(x2938), .I2(x2939), .I3(n5415), .I4(n5416), .O(n5417));
  LUT3 #(.INIT(8'hE8)) lut_n5418 (.I0(x2946), .I1(x2947), .I2(x2948), .O(n5418));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5419 (.I0(x2937), .I1(x2938), .I2(x2939), .I3(n5415), .I4(n5416), .O(n5419));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5420 (.I0(x2943), .I1(x2944), .I2(x2945), .I3(n5418), .I4(n5419), .O(n5420));
  LUT3 #(.INIT(8'h96)) lut_n5421 (.I0(n5409), .I1(n5412), .I2(n5413), .O(n5421));
  LUT3 #(.INIT(8'hE8)) lut_n5422 (.I0(n5417), .I1(n5420), .I2(n5421), .O(n5422));
  LUT3 #(.INIT(8'h96)) lut_n5423 (.I0(n5394), .I1(n5402), .I2(n5403), .O(n5423));
  LUT3 #(.INIT(8'hE8)) lut_n5424 (.I0(n5414), .I1(n5422), .I2(n5423), .O(n5424));
  LUT3 #(.INIT(8'hE8)) lut_n5425 (.I0(x2952), .I1(x2953), .I2(x2954), .O(n5425));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5426 (.I0(x2943), .I1(x2944), .I2(x2945), .I3(n5418), .I4(n5419), .O(n5426));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5427 (.I0(x2949), .I1(x2950), .I2(x2951), .I3(n5425), .I4(n5426), .O(n5427));
  LUT3 #(.INIT(8'hE8)) lut_n5428 (.I0(x2958), .I1(x2959), .I2(x2960), .O(n5428));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5429 (.I0(x2949), .I1(x2950), .I2(x2951), .I3(n5425), .I4(n5426), .O(n5429));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5430 (.I0(x2955), .I1(x2956), .I2(x2957), .I3(n5428), .I4(n5429), .O(n5430));
  LUT3 #(.INIT(8'h96)) lut_n5431 (.I0(n5417), .I1(n5420), .I2(n5421), .O(n5431));
  LUT3 #(.INIT(8'hE8)) lut_n5432 (.I0(n5427), .I1(n5430), .I2(n5431), .O(n5432));
  LUT3 #(.INIT(8'hE8)) lut_n5433 (.I0(x2964), .I1(x2965), .I2(x2966), .O(n5433));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5434 (.I0(x2955), .I1(x2956), .I2(x2957), .I3(n5428), .I4(n5429), .O(n5434));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5435 (.I0(x2961), .I1(x2962), .I2(x2963), .I3(n5433), .I4(n5434), .O(n5435));
  LUT3 #(.INIT(8'hE8)) lut_n5436 (.I0(x2970), .I1(x2971), .I2(x2972), .O(n5436));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5437 (.I0(x2961), .I1(x2962), .I2(x2963), .I3(n5433), .I4(n5434), .O(n5437));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5438 (.I0(x2967), .I1(x2968), .I2(x2969), .I3(n5436), .I4(n5437), .O(n5438));
  LUT3 #(.INIT(8'h96)) lut_n5439 (.I0(n5427), .I1(n5430), .I2(n5431), .O(n5439));
  LUT3 #(.INIT(8'hE8)) lut_n5440 (.I0(n5435), .I1(n5438), .I2(n5439), .O(n5440));
  LUT3 #(.INIT(8'h96)) lut_n5441 (.I0(n5414), .I1(n5422), .I2(n5423), .O(n5441));
  LUT3 #(.INIT(8'hE8)) lut_n5442 (.I0(n5432), .I1(n5440), .I2(n5441), .O(n5442));
  LUT3 #(.INIT(8'h96)) lut_n5443 (.I0(n5386), .I1(n5404), .I2(n5405), .O(n5443));
  LUT3 #(.INIT(8'hE8)) lut_n5444 (.I0(n5424), .I1(n5442), .I2(n5443), .O(n5444));
  LUT3 #(.INIT(8'h96)) lut_n5445 (.I0(n5326), .I1(n5364), .I2(n5365), .O(n5445));
  LUT3 #(.INIT(8'hE8)) lut_n5446 (.I0(n5406), .I1(n5444), .I2(n5445), .O(n5446));
  LUT3 #(.INIT(8'hE8)) lut_n5447 (.I0(x2976), .I1(x2977), .I2(x2978), .O(n5447));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5448 (.I0(x2967), .I1(x2968), .I2(x2969), .I3(n5436), .I4(n5437), .O(n5448));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5449 (.I0(x2973), .I1(x2974), .I2(x2975), .I3(n5447), .I4(n5448), .O(n5449));
  LUT3 #(.INIT(8'hE8)) lut_n5450 (.I0(x2982), .I1(x2983), .I2(x2984), .O(n5450));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5451 (.I0(x2973), .I1(x2974), .I2(x2975), .I3(n5447), .I4(n5448), .O(n5451));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5452 (.I0(x2979), .I1(x2980), .I2(x2981), .I3(n5450), .I4(n5451), .O(n5452));
  LUT3 #(.INIT(8'h96)) lut_n5453 (.I0(n5435), .I1(n5438), .I2(n5439), .O(n5453));
  LUT3 #(.INIT(8'hE8)) lut_n5454 (.I0(n5449), .I1(n5452), .I2(n5453), .O(n5454));
  LUT3 #(.INIT(8'hE8)) lut_n5455 (.I0(x2988), .I1(x2989), .I2(x2990), .O(n5455));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5456 (.I0(x2979), .I1(x2980), .I2(x2981), .I3(n5450), .I4(n5451), .O(n5456));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5457 (.I0(x2985), .I1(x2986), .I2(x2987), .I3(n5455), .I4(n5456), .O(n5457));
  LUT3 #(.INIT(8'hE8)) lut_n5458 (.I0(x2994), .I1(x2995), .I2(x2996), .O(n5458));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5459 (.I0(x2985), .I1(x2986), .I2(x2987), .I3(n5455), .I4(n5456), .O(n5459));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5460 (.I0(x2991), .I1(x2992), .I2(x2993), .I3(n5458), .I4(n5459), .O(n5460));
  LUT3 #(.INIT(8'h96)) lut_n5461 (.I0(n5449), .I1(n5452), .I2(n5453), .O(n5461));
  LUT3 #(.INIT(8'hE8)) lut_n5462 (.I0(n5457), .I1(n5460), .I2(n5461), .O(n5462));
  LUT3 #(.INIT(8'h96)) lut_n5463 (.I0(n5432), .I1(n5440), .I2(n5441), .O(n5463));
  LUT3 #(.INIT(8'hE8)) lut_n5464 (.I0(n5454), .I1(n5462), .I2(n5463), .O(n5464));
  LUT3 #(.INIT(8'h96)) lut_n5465 (.I0(x0), .I1(x1), .I2(x2), .O(n5465));
  LUT3 #(.INIT(8'h96)) lut_n5466 (.I0(x6), .I1(x7), .I2(x8), .O(n5466));
  LUT5 #(.INIT(32'hFF969600)) lut_n5467 (.I0(x3), .I1(x4), .I2(x5), .I3(n5465), .I4(n5466), .O(n5467));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5468 (.I0(x2991), .I1(x2992), .I2(x2993), .I3(n5458), .I4(n5459), .O(n5468));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5469 (.I0(x2997), .I1(x2998), .I2(x2999), .I3(n5467), .I4(n5468), .O(n5469));
  LUT3 #(.INIT(8'h96)) lut_n5470 (.I0(x12), .I1(x13), .I2(x14), .O(n5470));
  LUT5 #(.INIT(32'h96696996)) lut_n5471 (.I0(x3), .I1(x4), .I2(x5), .I3(n5465), .I4(n5466), .O(n5471));
  LUT5 #(.INIT(32'hFF969600)) lut_n5472 (.I0(x9), .I1(x10), .I2(x11), .I3(n5470), .I4(n5471), .O(n5472));
  LUT3 #(.INIT(8'h96)) lut_n5473 (.I0(x18), .I1(x19), .I2(x20), .O(n5473));
  LUT5 #(.INIT(32'h96696996)) lut_n5474 (.I0(x9), .I1(x10), .I2(x11), .I3(n5470), .I4(n5471), .O(n5474));
  LUT5 #(.INIT(32'hFF969600)) lut_n5475 (.I0(x15), .I1(x16), .I2(x17), .I3(n5473), .I4(n5474), .O(n5475));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5476 (.I0(x2997), .I1(x2998), .I2(x2999), .I3(n5467), .I4(n5468), .O(n5476));
  LUT3 #(.INIT(8'hE8)) lut_n5477 (.I0(n5472), .I1(n5475), .I2(n5476), .O(n5477));
  LUT3 #(.INIT(8'h96)) lut_n5478 (.I0(n5457), .I1(n5460), .I2(n5461), .O(n5478));
  LUT3 #(.INIT(8'hE8)) lut_n5479 (.I0(n5469), .I1(n5477), .I2(n5478), .O(n5479));
  LUT3 #(.INIT(8'h96)) lut_n5480 (.I0(x24), .I1(x25), .I2(x26), .O(n5480));
  LUT5 #(.INIT(32'h96696996)) lut_n5481 (.I0(x15), .I1(x16), .I2(x17), .I3(n5473), .I4(n5474), .O(n5481));
  LUT5 #(.INIT(32'hFF969600)) lut_n5482 (.I0(x21), .I1(x22), .I2(x23), .I3(n5480), .I4(n5481), .O(n5482));
  LUT3 #(.INIT(8'h96)) lut_n5483 (.I0(x27), .I1(x28), .I2(x29), .O(n5483));
  LUT5 #(.INIT(32'h96696996)) lut_n5484 (.I0(x21), .I1(x22), .I2(x23), .I3(n5480), .I4(n5481), .O(n5484));
  LUT5 #(.INIT(32'hFF969600)) lut_n5485 (.I0(x30), .I1(x31), .I2(x32), .I3(n5483), .I4(n5484), .O(n5485));
  LUT3 #(.INIT(8'h96)) lut_n5486 (.I0(n5472), .I1(n5475), .I2(n5476), .O(n5486));
  LUT3 #(.INIT(8'hE8)) lut_n5487 (.I0(n5482), .I1(n5485), .I2(n5486), .O(n5487));
  LUT3 #(.INIT(8'h96)) lut_n5488 (.I0(x36), .I1(x37), .I2(x38), .O(n5488));
  LUT5 #(.INIT(32'h96696996)) lut_n5489 (.I0(x30), .I1(x31), .I2(x32), .I3(n5483), .I4(n5484), .O(n5489));
  LUT5 #(.INIT(32'hFF969600)) lut_n5490 (.I0(x33), .I1(x34), .I2(x35), .I3(n5488), .I4(n5489), .O(n5490));
  LUT3 #(.INIT(8'h96)) lut_n5491 (.I0(x42), .I1(x43), .I2(x44), .O(n5491));
  LUT5 #(.INIT(32'h96696996)) lut_n5492 (.I0(x33), .I1(x34), .I2(x35), .I3(n5488), .I4(n5489), .O(n5492));
  LUT5 #(.INIT(32'hFF969600)) lut_n5493 (.I0(x39), .I1(x40), .I2(x41), .I3(n5491), .I4(n5492), .O(n5493));
  LUT3 #(.INIT(8'h96)) lut_n5494 (.I0(n5482), .I1(n5485), .I2(n5486), .O(n5494));
  LUT3 #(.INIT(8'hE8)) lut_n5495 (.I0(n5490), .I1(n5493), .I2(n5494), .O(n5495));
  LUT3 #(.INIT(8'h96)) lut_n5496 (.I0(n5469), .I1(n5477), .I2(n5478), .O(n5496));
  LUT3 #(.INIT(8'hE8)) lut_n5497 (.I0(n5487), .I1(n5495), .I2(n5496), .O(n5497));
  LUT3 #(.INIT(8'h96)) lut_n5498 (.I0(n5454), .I1(n5462), .I2(n5463), .O(n5498));
  LUT3 #(.INIT(8'hE8)) lut_n5499 (.I0(n5479), .I1(n5497), .I2(n5498), .O(n5499));
  LUT3 #(.INIT(8'h96)) lut_n5500 (.I0(n5424), .I1(n5442), .I2(n5443), .O(n5500));
  LUT3 #(.INIT(8'hE8)) lut_n5501 (.I0(n5464), .I1(n5499), .I2(n5500), .O(n5501));
  LUT3 #(.INIT(8'h96)) lut_n5502 (.I0(x48), .I1(x49), .I2(x50), .O(n5502));
  LUT5 #(.INIT(32'h96696996)) lut_n5503 (.I0(x39), .I1(x40), .I2(x41), .I3(n5491), .I4(n5492), .O(n5503));
  LUT5 #(.INIT(32'hFF969600)) lut_n5504 (.I0(x45), .I1(x46), .I2(x47), .I3(n5502), .I4(n5503), .O(n5504));
  LUT3 #(.INIT(8'h96)) lut_n5505 (.I0(x54), .I1(x55), .I2(x56), .O(n5505));
  LUT5 #(.INIT(32'h96696996)) lut_n5506 (.I0(x45), .I1(x46), .I2(x47), .I3(n5502), .I4(n5503), .O(n5506));
  LUT5 #(.INIT(32'hFF969600)) lut_n5507 (.I0(x51), .I1(x52), .I2(x53), .I3(n5505), .I4(n5506), .O(n5507));
  LUT3 #(.INIT(8'h96)) lut_n5508 (.I0(n5490), .I1(n5493), .I2(n5494), .O(n5508));
  LUT3 #(.INIT(8'hE8)) lut_n5509 (.I0(n5504), .I1(n5507), .I2(n5508), .O(n5509));
  LUT3 #(.INIT(8'h96)) lut_n5510 (.I0(x60), .I1(x61), .I2(x62), .O(n5510));
  LUT5 #(.INIT(32'h96696996)) lut_n5511 (.I0(x51), .I1(x52), .I2(x53), .I3(n5505), .I4(n5506), .O(n5511));
  LUT5 #(.INIT(32'hFF969600)) lut_n5512 (.I0(x57), .I1(x58), .I2(x59), .I3(n5510), .I4(n5511), .O(n5512));
  LUT3 #(.INIT(8'h96)) lut_n5513 (.I0(x66), .I1(x67), .I2(x68), .O(n5513));
  LUT5 #(.INIT(32'h96696996)) lut_n5514 (.I0(x57), .I1(x58), .I2(x59), .I3(n5510), .I4(n5511), .O(n5514));
  LUT5 #(.INIT(32'hFF969600)) lut_n5515 (.I0(x63), .I1(x64), .I2(x65), .I3(n5513), .I4(n5514), .O(n5515));
  LUT3 #(.INIT(8'h96)) lut_n5516 (.I0(n5504), .I1(n5507), .I2(n5508), .O(n5516));
  LUT3 #(.INIT(8'hE8)) lut_n5517 (.I0(n5512), .I1(n5515), .I2(n5516), .O(n5517));
  LUT3 #(.INIT(8'h96)) lut_n5518 (.I0(n5487), .I1(n5495), .I2(n5496), .O(n5518));
  LUT3 #(.INIT(8'hE8)) lut_n5519 (.I0(n5509), .I1(n5517), .I2(n5518), .O(n5519));
  LUT3 #(.INIT(8'h96)) lut_n5520 (.I0(x72), .I1(x73), .I2(x74), .O(n5520));
  LUT5 #(.INIT(32'h96696996)) lut_n5521 (.I0(x63), .I1(x64), .I2(x65), .I3(n5513), .I4(n5514), .O(n5521));
  LUT5 #(.INIT(32'hFF969600)) lut_n5522 (.I0(x69), .I1(x70), .I2(x71), .I3(n5520), .I4(n5521), .O(n5522));
  LUT3 #(.INIT(8'h96)) lut_n5523 (.I0(x78), .I1(x79), .I2(x80), .O(n5523));
  LUT5 #(.INIT(32'h96696996)) lut_n5524 (.I0(x69), .I1(x70), .I2(x71), .I3(n5520), .I4(n5521), .O(n5524));
  LUT5 #(.INIT(32'hFF969600)) lut_n5525 (.I0(x75), .I1(x76), .I2(x77), .I3(n5523), .I4(n5524), .O(n5525));
  LUT3 #(.INIT(8'h96)) lut_n5526 (.I0(n5512), .I1(n5515), .I2(n5516), .O(n5526));
  LUT3 #(.INIT(8'hE8)) lut_n5527 (.I0(n5522), .I1(n5525), .I2(n5526), .O(n5527));
  LUT3 #(.INIT(8'h96)) lut_n5528 (.I0(x84), .I1(x85), .I2(x86), .O(n5528));
  LUT5 #(.INIT(32'h96696996)) lut_n5529 (.I0(x75), .I1(x76), .I2(x77), .I3(n5523), .I4(n5524), .O(n5529));
  LUT5 #(.INIT(32'hFF969600)) lut_n5530 (.I0(x81), .I1(x82), .I2(x83), .I3(n5528), .I4(n5529), .O(n5530));
  LUT3 #(.INIT(8'h96)) lut_n5531 (.I0(x90), .I1(x91), .I2(x92), .O(n5531));
  LUT5 #(.INIT(32'h96696996)) lut_n5532 (.I0(x81), .I1(x82), .I2(x83), .I3(n5528), .I4(n5529), .O(n5532));
  LUT5 #(.INIT(32'hFF969600)) lut_n5533 (.I0(x87), .I1(x88), .I2(x89), .I3(n5531), .I4(n5532), .O(n5533));
  LUT3 #(.INIT(8'h96)) lut_n5534 (.I0(n5522), .I1(n5525), .I2(n5526), .O(n5534));
  LUT3 #(.INIT(8'hE8)) lut_n5535 (.I0(n5530), .I1(n5533), .I2(n5534), .O(n5535));
  LUT3 #(.INIT(8'h96)) lut_n5536 (.I0(n5509), .I1(n5517), .I2(n5518), .O(n5536));
  LUT3 #(.INIT(8'hE8)) lut_n5537 (.I0(n5527), .I1(n5535), .I2(n5536), .O(n5537));
  LUT3 #(.INIT(8'h96)) lut_n5538 (.I0(n5479), .I1(n5497), .I2(n5498), .O(n5538));
  LUT3 #(.INIT(8'hE8)) lut_n5539 (.I0(n5519), .I1(n5537), .I2(n5538), .O(n5539));
  LUT3 #(.INIT(8'h96)) lut_n5540 (.I0(x96), .I1(x97), .I2(x98), .O(n5540));
  LUT5 #(.INIT(32'h96696996)) lut_n5541 (.I0(x87), .I1(x88), .I2(x89), .I3(n5531), .I4(n5532), .O(n5541));
  LUT5 #(.INIT(32'hFF969600)) lut_n5542 (.I0(x93), .I1(x94), .I2(x95), .I3(n5540), .I4(n5541), .O(n5542));
  LUT3 #(.INIT(8'h96)) lut_n5543 (.I0(x102), .I1(x103), .I2(x104), .O(n5543));
  LUT5 #(.INIT(32'h96696996)) lut_n5544 (.I0(x93), .I1(x94), .I2(x95), .I3(n5540), .I4(n5541), .O(n5544));
  LUT5 #(.INIT(32'hFF969600)) lut_n5545 (.I0(x99), .I1(x100), .I2(x101), .I3(n5543), .I4(n5544), .O(n5545));
  LUT3 #(.INIT(8'h96)) lut_n5546 (.I0(n5530), .I1(n5533), .I2(n5534), .O(n5546));
  LUT3 #(.INIT(8'hE8)) lut_n5547 (.I0(n5542), .I1(n5545), .I2(n5546), .O(n5547));
  LUT3 #(.INIT(8'h96)) lut_n5548 (.I0(x108), .I1(x109), .I2(x110), .O(n5548));
  LUT5 #(.INIT(32'h96696996)) lut_n5549 (.I0(x99), .I1(x100), .I2(x101), .I3(n5543), .I4(n5544), .O(n5549));
  LUT5 #(.INIT(32'hFF969600)) lut_n5550 (.I0(x105), .I1(x106), .I2(x107), .I3(n5548), .I4(n5549), .O(n5550));
  LUT3 #(.INIT(8'h96)) lut_n5551 (.I0(x114), .I1(x115), .I2(x116), .O(n5551));
  LUT5 #(.INIT(32'h96696996)) lut_n5552 (.I0(x105), .I1(x106), .I2(x107), .I3(n5548), .I4(n5549), .O(n5552));
  LUT5 #(.INIT(32'hFF969600)) lut_n5553 (.I0(x111), .I1(x112), .I2(x113), .I3(n5551), .I4(n5552), .O(n5553));
  LUT3 #(.INIT(8'h96)) lut_n5554 (.I0(n5542), .I1(n5545), .I2(n5546), .O(n5554));
  LUT3 #(.INIT(8'hE8)) lut_n5555 (.I0(n5550), .I1(n5553), .I2(n5554), .O(n5555));
  LUT3 #(.INIT(8'h96)) lut_n5556 (.I0(n5527), .I1(n5535), .I2(n5536), .O(n5556));
  LUT3 #(.INIT(8'hE8)) lut_n5557 (.I0(n5547), .I1(n5555), .I2(n5556), .O(n5557));
  LUT3 #(.INIT(8'h96)) lut_n5558 (.I0(x120), .I1(x121), .I2(x122), .O(n5558));
  LUT5 #(.INIT(32'h96696996)) lut_n5559 (.I0(x111), .I1(x112), .I2(x113), .I3(n5551), .I4(n5552), .O(n5559));
  LUT5 #(.INIT(32'hFF969600)) lut_n5560 (.I0(x117), .I1(x118), .I2(x119), .I3(n5558), .I4(n5559), .O(n5560));
  LUT3 #(.INIT(8'h96)) lut_n5561 (.I0(x126), .I1(x127), .I2(x128), .O(n5561));
  LUT5 #(.INIT(32'h96696996)) lut_n5562 (.I0(x117), .I1(x118), .I2(x119), .I3(n5558), .I4(n5559), .O(n5562));
  LUT5 #(.INIT(32'hFF969600)) lut_n5563 (.I0(x123), .I1(x124), .I2(x125), .I3(n5561), .I4(n5562), .O(n5563));
  LUT3 #(.INIT(8'h96)) lut_n5564 (.I0(n5550), .I1(n5553), .I2(n5554), .O(n5564));
  LUT3 #(.INIT(8'hE8)) lut_n5565 (.I0(n5560), .I1(n5563), .I2(n5564), .O(n5565));
  LUT3 #(.INIT(8'h96)) lut_n5566 (.I0(x132), .I1(x133), .I2(x134), .O(n5566));
  LUT5 #(.INIT(32'h96696996)) lut_n5567 (.I0(x123), .I1(x124), .I2(x125), .I3(n5561), .I4(n5562), .O(n5567));
  LUT5 #(.INIT(32'hFF969600)) lut_n5568 (.I0(x129), .I1(x130), .I2(x131), .I3(n5566), .I4(n5567), .O(n5568));
  LUT3 #(.INIT(8'h96)) lut_n5569 (.I0(x138), .I1(x139), .I2(x140), .O(n5569));
  LUT5 #(.INIT(32'h96696996)) lut_n5570 (.I0(x129), .I1(x130), .I2(x131), .I3(n5566), .I4(n5567), .O(n5570));
  LUT5 #(.INIT(32'hFF969600)) lut_n5571 (.I0(x135), .I1(x136), .I2(x137), .I3(n5569), .I4(n5570), .O(n5571));
  LUT3 #(.INIT(8'h96)) lut_n5572 (.I0(n5560), .I1(n5563), .I2(n5564), .O(n5572));
  LUT3 #(.INIT(8'hE8)) lut_n5573 (.I0(n5568), .I1(n5571), .I2(n5572), .O(n5573));
  LUT3 #(.INIT(8'h96)) lut_n5574 (.I0(n5547), .I1(n5555), .I2(n5556), .O(n5574));
  LUT3 #(.INIT(8'hE8)) lut_n5575 (.I0(n5565), .I1(n5573), .I2(n5574), .O(n5575));
  LUT3 #(.INIT(8'h96)) lut_n5576 (.I0(n5519), .I1(n5537), .I2(n5538), .O(n5576));
  LUT3 #(.INIT(8'hE8)) lut_n5577 (.I0(n5557), .I1(n5575), .I2(n5576), .O(n5577));
  LUT3 #(.INIT(8'h96)) lut_n5578 (.I0(n5464), .I1(n5499), .I2(n5500), .O(n5578));
  LUT3 #(.INIT(8'hE8)) lut_n5579 (.I0(n5539), .I1(n5577), .I2(n5578), .O(n5579));
  LUT3 #(.INIT(8'h96)) lut_n5580 (.I0(n5406), .I1(n5444), .I2(n5445), .O(n5580));
  LUT3 #(.INIT(8'hE8)) lut_n5581 (.I0(n5501), .I1(n5579), .I2(n5580), .O(n5581));
  LUT3 #(.INIT(8'h96)) lut_n5582 (.I0(n5288), .I1(n5366), .I2(n5367), .O(n5582));
  LUT3 #(.INIT(8'hE8)) lut_n5583 (.I0(n5446), .I1(n5581), .I2(n5582), .O(n5583));
  LUT3 #(.INIT(8'h96)) lut_n5584 (.I0(n5050), .I1(n5208), .I2(n5209), .O(n5584));
  LUT3 #(.INIT(8'hE8)) lut_n5585 (.I0(n5368), .I1(n5583), .I2(n5584), .O(n5585));
  LUT3 #(.INIT(8'h96)) lut_n5586 (.I0(n4572), .I1(n4890), .I2(n4891), .O(n5586));
  LUT3 #(.INIT(8'hE8)) lut_n5587 (.I0(n5210), .I1(n5585), .I2(n5586), .O(n5587));
  LUT3 #(.INIT(8'hE8)) lut_n5588 (.I0(n4254), .I1(n4892), .I2(n5587), .O(n5588));
  LUT3 #(.INIT(8'h96)) lut_n5589 (.I0(x144), .I1(x145), .I2(x146), .O(n5589));
  LUT5 #(.INIT(32'h96696996)) lut_n5590 (.I0(x135), .I1(x136), .I2(x137), .I3(n5569), .I4(n5570), .O(n5590));
  LUT5 #(.INIT(32'hFF969600)) lut_n5591 (.I0(x141), .I1(x142), .I2(x143), .I3(n5589), .I4(n5590), .O(n5591));
  LUT3 #(.INIT(8'h96)) lut_n5592 (.I0(x150), .I1(x151), .I2(x152), .O(n5592));
  LUT5 #(.INIT(32'h96696996)) lut_n5593 (.I0(x141), .I1(x142), .I2(x143), .I3(n5589), .I4(n5590), .O(n5593));
  LUT5 #(.INIT(32'hFF969600)) lut_n5594 (.I0(x147), .I1(x148), .I2(x149), .I3(n5592), .I4(n5593), .O(n5594));
  LUT3 #(.INIT(8'h96)) lut_n5595 (.I0(n5568), .I1(n5571), .I2(n5572), .O(n5595));
  LUT3 #(.INIT(8'hE8)) lut_n5596 (.I0(n5591), .I1(n5594), .I2(n5595), .O(n5596));
  LUT3 #(.INIT(8'h96)) lut_n5597 (.I0(x156), .I1(x157), .I2(x158), .O(n5597));
  LUT5 #(.INIT(32'h96696996)) lut_n5598 (.I0(x147), .I1(x148), .I2(x149), .I3(n5592), .I4(n5593), .O(n5598));
  LUT5 #(.INIT(32'hFF969600)) lut_n5599 (.I0(x153), .I1(x154), .I2(x155), .I3(n5597), .I4(n5598), .O(n5599));
  LUT3 #(.INIT(8'h96)) lut_n5600 (.I0(x162), .I1(x163), .I2(x164), .O(n5600));
  LUT5 #(.INIT(32'h96696996)) lut_n5601 (.I0(x153), .I1(x154), .I2(x155), .I3(n5597), .I4(n5598), .O(n5601));
  LUT5 #(.INIT(32'hFF969600)) lut_n5602 (.I0(x159), .I1(x160), .I2(x161), .I3(n5600), .I4(n5601), .O(n5602));
  LUT3 #(.INIT(8'h96)) lut_n5603 (.I0(n5591), .I1(n5594), .I2(n5595), .O(n5603));
  LUT3 #(.INIT(8'hE8)) lut_n5604 (.I0(n5599), .I1(n5602), .I2(n5603), .O(n5604));
  LUT3 #(.INIT(8'h96)) lut_n5605 (.I0(n5565), .I1(n5573), .I2(n5574), .O(n5605));
  LUT3 #(.INIT(8'hE8)) lut_n5606 (.I0(n5596), .I1(n5604), .I2(n5605), .O(n5606));
  LUT3 #(.INIT(8'h96)) lut_n5607 (.I0(x168), .I1(x169), .I2(x170), .O(n5607));
  LUT5 #(.INIT(32'h96696996)) lut_n5608 (.I0(x159), .I1(x160), .I2(x161), .I3(n5600), .I4(n5601), .O(n5608));
  LUT5 #(.INIT(32'hFF969600)) lut_n5609 (.I0(x165), .I1(x166), .I2(x167), .I3(n5607), .I4(n5608), .O(n5609));
  LUT3 #(.INIT(8'h96)) lut_n5610 (.I0(x174), .I1(x175), .I2(x176), .O(n5610));
  LUT5 #(.INIT(32'h96696996)) lut_n5611 (.I0(x165), .I1(x166), .I2(x167), .I3(n5607), .I4(n5608), .O(n5611));
  LUT5 #(.INIT(32'hFF969600)) lut_n5612 (.I0(x171), .I1(x172), .I2(x173), .I3(n5610), .I4(n5611), .O(n5612));
  LUT3 #(.INIT(8'h96)) lut_n5613 (.I0(n5599), .I1(n5602), .I2(n5603), .O(n5613));
  LUT3 #(.INIT(8'hE8)) lut_n5614 (.I0(n5609), .I1(n5612), .I2(n5613), .O(n5614));
  LUT3 #(.INIT(8'h96)) lut_n5615 (.I0(x180), .I1(x181), .I2(x182), .O(n5615));
  LUT5 #(.INIT(32'h96696996)) lut_n5616 (.I0(x171), .I1(x172), .I2(x173), .I3(n5610), .I4(n5611), .O(n5616));
  LUT5 #(.INIT(32'hFF969600)) lut_n5617 (.I0(x177), .I1(x178), .I2(x179), .I3(n5615), .I4(n5616), .O(n5617));
  LUT3 #(.INIT(8'h96)) lut_n5618 (.I0(x186), .I1(x187), .I2(x188), .O(n5618));
  LUT5 #(.INIT(32'h96696996)) lut_n5619 (.I0(x177), .I1(x178), .I2(x179), .I3(n5615), .I4(n5616), .O(n5619));
  LUT5 #(.INIT(32'hFF969600)) lut_n5620 (.I0(x183), .I1(x184), .I2(x185), .I3(n5618), .I4(n5619), .O(n5620));
  LUT3 #(.INIT(8'h96)) lut_n5621 (.I0(n5609), .I1(n5612), .I2(n5613), .O(n5621));
  LUT3 #(.INIT(8'hE8)) lut_n5622 (.I0(n5617), .I1(n5620), .I2(n5621), .O(n5622));
  LUT3 #(.INIT(8'h96)) lut_n5623 (.I0(n5596), .I1(n5604), .I2(n5605), .O(n5623));
  LUT3 #(.INIT(8'hE8)) lut_n5624 (.I0(n5614), .I1(n5622), .I2(n5623), .O(n5624));
  LUT3 #(.INIT(8'h96)) lut_n5625 (.I0(n5557), .I1(n5575), .I2(n5576), .O(n5625));
  LUT3 #(.INIT(8'hE8)) lut_n5626 (.I0(n5606), .I1(n5624), .I2(n5625), .O(n5626));
  LUT3 #(.INIT(8'h96)) lut_n5627 (.I0(x192), .I1(x193), .I2(x194), .O(n5627));
  LUT5 #(.INIT(32'h96696996)) lut_n5628 (.I0(x183), .I1(x184), .I2(x185), .I3(n5618), .I4(n5619), .O(n5628));
  LUT5 #(.INIT(32'hFF969600)) lut_n5629 (.I0(x189), .I1(x190), .I2(x191), .I3(n5627), .I4(n5628), .O(n5629));
  LUT3 #(.INIT(8'h96)) lut_n5630 (.I0(x198), .I1(x199), .I2(x200), .O(n5630));
  LUT5 #(.INIT(32'h96696996)) lut_n5631 (.I0(x189), .I1(x190), .I2(x191), .I3(n5627), .I4(n5628), .O(n5631));
  LUT5 #(.INIT(32'hFF969600)) lut_n5632 (.I0(x195), .I1(x196), .I2(x197), .I3(n5630), .I4(n5631), .O(n5632));
  LUT3 #(.INIT(8'h96)) lut_n5633 (.I0(n5617), .I1(n5620), .I2(n5621), .O(n5633));
  LUT3 #(.INIT(8'hE8)) lut_n5634 (.I0(n5629), .I1(n5632), .I2(n5633), .O(n5634));
  LUT3 #(.INIT(8'h96)) lut_n5635 (.I0(x204), .I1(x205), .I2(x206), .O(n5635));
  LUT5 #(.INIT(32'h96696996)) lut_n5636 (.I0(x195), .I1(x196), .I2(x197), .I3(n5630), .I4(n5631), .O(n5636));
  LUT5 #(.INIT(32'hFF969600)) lut_n5637 (.I0(x201), .I1(x202), .I2(x203), .I3(n5635), .I4(n5636), .O(n5637));
  LUT3 #(.INIT(8'h96)) lut_n5638 (.I0(x210), .I1(x211), .I2(x212), .O(n5638));
  LUT5 #(.INIT(32'h96696996)) lut_n5639 (.I0(x201), .I1(x202), .I2(x203), .I3(n5635), .I4(n5636), .O(n5639));
  LUT5 #(.INIT(32'hFF969600)) lut_n5640 (.I0(x207), .I1(x208), .I2(x209), .I3(n5638), .I4(n5639), .O(n5640));
  LUT3 #(.INIT(8'h96)) lut_n5641 (.I0(n5629), .I1(n5632), .I2(n5633), .O(n5641));
  LUT3 #(.INIT(8'hE8)) lut_n5642 (.I0(n5637), .I1(n5640), .I2(n5641), .O(n5642));
  LUT3 #(.INIT(8'h96)) lut_n5643 (.I0(n5614), .I1(n5622), .I2(n5623), .O(n5643));
  LUT3 #(.INIT(8'hE8)) lut_n5644 (.I0(n5634), .I1(n5642), .I2(n5643), .O(n5644));
  LUT3 #(.INIT(8'h96)) lut_n5645 (.I0(x216), .I1(x217), .I2(x218), .O(n5645));
  LUT5 #(.INIT(32'h96696996)) lut_n5646 (.I0(x207), .I1(x208), .I2(x209), .I3(n5638), .I4(n5639), .O(n5646));
  LUT5 #(.INIT(32'hFF969600)) lut_n5647 (.I0(x213), .I1(x214), .I2(x215), .I3(n5645), .I4(n5646), .O(n5647));
  LUT3 #(.INIT(8'h96)) lut_n5648 (.I0(x222), .I1(x223), .I2(x224), .O(n5648));
  LUT5 #(.INIT(32'h96696996)) lut_n5649 (.I0(x213), .I1(x214), .I2(x215), .I3(n5645), .I4(n5646), .O(n5649));
  LUT5 #(.INIT(32'hFF969600)) lut_n5650 (.I0(x219), .I1(x220), .I2(x221), .I3(n5648), .I4(n5649), .O(n5650));
  LUT3 #(.INIT(8'h96)) lut_n5651 (.I0(n5637), .I1(n5640), .I2(n5641), .O(n5651));
  LUT3 #(.INIT(8'hE8)) lut_n5652 (.I0(n5647), .I1(n5650), .I2(n5651), .O(n5652));
  LUT3 #(.INIT(8'h96)) lut_n5653 (.I0(x228), .I1(x229), .I2(x230), .O(n5653));
  LUT5 #(.INIT(32'h96696996)) lut_n5654 (.I0(x219), .I1(x220), .I2(x221), .I3(n5648), .I4(n5649), .O(n5654));
  LUT5 #(.INIT(32'hFF969600)) lut_n5655 (.I0(x225), .I1(x226), .I2(x227), .I3(n5653), .I4(n5654), .O(n5655));
  LUT3 #(.INIT(8'h96)) lut_n5656 (.I0(x234), .I1(x235), .I2(x236), .O(n5656));
  LUT5 #(.INIT(32'h96696996)) lut_n5657 (.I0(x225), .I1(x226), .I2(x227), .I3(n5653), .I4(n5654), .O(n5657));
  LUT5 #(.INIT(32'hFF969600)) lut_n5658 (.I0(x231), .I1(x232), .I2(x233), .I3(n5656), .I4(n5657), .O(n5658));
  LUT3 #(.INIT(8'h96)) lut_n5659 (.I0(n5647), .I1(n5650), .I2(n5651), .O(n5659));
  LUT3 #(.INIT(8'hE8)) lut_n5660 (.I0(n5655), .I1(n5658), .I2(n5659), .O(n5660));
  LUT3 #(.INIT(8'h96)) lut_n5661 (.I0(n5634), .I1(n5642), .I2(n5643), .O(n5661));
  LUT3 #(.INIT(8'hE8)) lut_n5662 (.I0(n5652), .I1(n5660), .I2(n5661), .O(n5662));
  LUT3 #(.INIT(8'h96)) lut_n5663 (.I0(n5606), .I1(n5624), .I2(n5625), .O(n5663));
  LUT3 #(.INIT(8'hE8)) lut_n5664 (.I0(n5644), .I1(n5662), .I2(n5663), .O(n5664));
  LUT3 #(.INIT(8'h96)) lut_n5665 (.I0(n5539), .I1(n5577), .I2(n5578), .O(n5665));
  LUT3 #(.INIT(8'hE8)) lut_n5666 (.I0(n5626), .I1(n5664), .I2(n5665), .O(n5666));
  LUT3 #(.INIT(8'h96)) lut_n5667 (.I0(x240), .I1(x241), .I2(x242), .O(n5667));
  LUT5 #(.INIT(32'h96696996)) lut_n5668 (.I0(x231), .I1(x232), .I2(x233), .I3(n5656), .I4(n5657), .O(n5668));
  LUT5 #(.INIT(32'hFF969600)) lut_n5669 (.I0(x237), .I1(x238), .I2(x239), .I3(n5667), .I4(n5668), .O(n5669));
  LUT3 #(.INIT(8'h96)) lut_n5670 (.I0(x246), .I1(x247), .I2(x248), .O(n5670));
  LUT5 #(.INIT(32'h96696996)) lut_n5671 (.I0(x237), .I1(x238), .I2(x239), .I3(n5667), .I4(n5668), .O(n5671));
  LUT5 #(.INIT(32'hFF969600)) lut_n5672 (.I0(x243), .I1(x244), .I2(x245), .I3(n5670), .I4(n5671), .O(n5672));
  LUT3 #(.INIT(8'h96)) lut_n5673 (.I0(n5655), .I1(n5658), .I2(n5659), .O(n5673));
  LUT3 #(.INIT(8'hE8)) lut_n5674 (.I0(n5669), .I1(n5672), .I2(n5673), .O(n5674));
  LUT3 #(.INIT(8'h96)) lut_n5675 (.I0(x252), .I1(x253), .I2(x254), .O(n5675));
  LUT5 #(.INIT(32'h96696996)) lut_n5676 (.I0(x243), .I1(x244), .I2(x245), .I3(n5670), .I4(n5671), .O(n5676));
  LUT5 #(.INIT(32'hFF969600)) lut_n5677 (.I0(x249), .I1(x250), .I2(x251), .I3(n5675), .I4(n5676), .O(n5677));
  LUT3 #(.INIT(8'h96)) lut_n5678 (.I0(x258), .I1(x259), .I2(x260), .O(n5678));
  LUT5 #(.INIT(32'h96696996)) lut_n5679 (.I0(x249), .I1(x250), .I2(x251), .I3(n5675), .I4(n5676), .O(n5679));
  LUT5 #(.INIT(32'hFF969600)) lut_n5680 (.I0(x255), .I1(x256), .I2(x257), .I3(n5678), .I4(n5679), .O(n5680));
  LUT3 #(.INIT(8'h96)) lut_n5681 (.I0(n5669), .I1(n5672), .I2(n5673), .O(n5681));
  LUT3 #(.INIT(8'hE8)) lut_n5682 (.I0(n5677), .I1(n5680), .I2(n5681), .O(n5682));
  LUT3 #(.INIT(8'h96)) lut_n5683 (.I0(n5652), .I1(n5660), .I2(n5661), .O(n5683));
  LUT3 #(.INIT(8'hE8)) lut_n5684 (.I0(n5674), .I1(n5682), .I2(n5683), .O(n5684));
  LUT3 #(.INIT(8'h96)) lut_n5685 (.I0(x264), .I1(x265), .I2(x266), .O(n5685));
  LUT5 #(.INIT(32'h96696996)) lut_n5686 (.I0(x255), .I1(x256), .I2(x257), .I3(n5678), .I4(n5679), .O(n5686));
  LUT5 #(.INIT(32'hFF969600)) lut_n5687 (.I0(x261), .I1(x262), .I2(x263), .I3(n5685), .I4(n5686), .O(n5687));
  LUT3 #(.INIT(8'h96)) lut_n5688 (.I0(x270), .I1(x271), .I2(x272), .O(n5688));
  LUT5 #(.INIT(32'h96696996)) lut_n5689 (.I0(x261), .I1(x262), .I2(x263), .I3(n5685), .I4(n5686), .O(n5689));
  LUT5 #(.INIT(32'hFF969600)) lut_n5690 (.I0(x267), .I1(x268), .I2(x269), .I3(n5688), .I4(n5689), .O(n5690));
  LUT3 #(.INIT(8'h96)) lut_n5691 (.I0(n5677), .I1(n5680), .I2(n5681), .O(n5691));
  LUT3 #(.INIT(8'hE8)) lut_n5692 (.I0(n5687), .I1(n5690), .I2(n5691), .O(n5692));
  LUT3 #(.INIT(8'h96)) lut_n5693 (.I0(x276), .I1(x277), .I2(x278), .O(n5693));
  LUT5 #(.INIT(32'h96696996)) lut_n5694 (.I0(x267), .I1(x268), .I2(x269), .I3(n5688), .I4(n5689), .O(n5694));
  LUT5 #(.INIT(32'hFF969600)) lut_n5695 (.I0(x273), .I1(x274), .I2(x275), .I3(n5693), .I4(n5694), .O(n5695));
  LUT3 #(.INIT(8'h96)) lut_n5696 (.I0(x282), .I1(x283), .I2(x284), .O(n5696));
  LUT5 #(.INIT(32'h96696996)) lut_n5697 (.I0(x273), .I1(x274), .I2(x275), .I3(n5693), .I4(n5694), .O(n5697));
  LUT5 #(.INIT(32'hFF969600)) lut_n5698 (.I0(x279), .I1(x280), .I2(x281), .I3(n5696), .I4(n5697), .O(n5698));
  LUT3 #(.INIT(8'h96)) lut_n5699 (.I0(n5687), .I1(n5690), .I2(n5691), .O(n5699));
  LUT3 #(.INIT(8'hE8)) lut_n5700 (.I0(n5695), .I1(n5698), .I2(n5699), .O(n5700));
  LUT3 #(.INIT(8'h96)) lut_n5701 (.I0(n5674), .I1(n5682), .I2(n5683), .O(n5701));
  LUT3 #(.INIT(8'hE8)) lut_n5702 (.I0(n5692), .I1(n5700), .I2(n5701), .O(n5702));
  LUT3 #(.INIT(8'h96)) lut_n5703 (.I0(n5644), .I1(n5662), .I2(n5663), .O(n5703));
  LUT3 #(.INIT(8'hE8)) lut_n5704 (.I0(n5684), .I1(n5702), .I2(n5703), .O(n5704));
  LUT3 #(.INIT(8'h96)) lut_n5705 (.I0(x288), .I1(x289), .I2(x290), .O(n5705));
  LUT5 #(.INIT(32'h96696996)) lut_n5706 (.I0(x279), .I1(x280), .I2(x281), .I3(n5696), .I4(n5697), .O(n5706));
  LUT5 #(.INIT(32'hFF969600)) lut_n5707 (.I0(x285), .I1(x286), .I2(x287), .I3(n5705), .I4(n5706), .O(n5707));
  LUT3 #(.INIT(8'h96)) lut_n5708 (.I0(x294), .I1(x295), .I2(x296), .O(n5708));
  LUT5 #(.INIT(32'h96696996)) lut_n5709 (.I0(x285), .I1(x286), .I2(x287), .I3(n5705), .I4(n5706), .O(n5709));
  LUT5 #(.INIT(32'hFF969600)) lut_n5710 (.I0(x291), .I1(x292), .I2(x293), .I3(n5708), .I4(n5709), .O(n5710));
  LUT3 #(.INIT(8'h96)) lut_n5711 (.I0(n5695), .I1(n5698), .I2(n5699), .O(n5711));
  LUT3 #(.INIT(8'hE8)) lut_n5712 (.I0(n5707), .I1(n5710), .I2(n5711), .O(n5712));
  LUT3 #(.INIT(8'h96)) lut_n5713 (.I0(x297), .I1(x298), .I2(x299), .O(n5713));
  LUT5 #(.INIT(32'h96696996)) lut_n5714 (.I0(x291), .I1(x292), .I2(x293), .I3(n5708), .I4(n5709), .O(n5714));
  LUT5 #(.INIT(32'hFF969600)) lut_n5715 (.I0(x300), .I1(x301), .I2(x302), .I3(n5713), .I4(n5714), .O(n5715));
  LUT3 #(.INIT(8'h96)) lut_n5716 (.I0(x306), .I1(x307), .I2(x308), .O(n5716));
  LUT5 #(.INIT(32'h96696996)) lut_n5717 (.I0(x300), .I1(x301), .I2(x302), .I3(n5713), .I4(n5714), .O(n5717));
  LUT5 #(.INIT(32'hFF969600)) lut_n5718 (.I0(x303), .I1(x304), .I2(x305), .I3(n5716), .I4(n5717), .O(n5718));
  LUT3 #(.INIT(8'h96)) lut_n5719 (.I0(n5707), .I1(n5710), .I2(n5711), .O(n5719));
  LUT3 #(.INIT(8'hE8)) lut_n5720 (.I0(n5715), .I1(n5718), .I2(n5719), .O(n5720));
  LUT3 #(.INIT(8'h96)) lut_n5721 (.I0(n5692), .I1(n5700), .I2(n5701), .O(n5721));
  LUT3 #(.INIT(8'hE8)) lut_n5722 (.I0(n5712), .I1(n5720), .I2(n5721), .O(n5722));
  LUT3 #(.INIT(8'h96)) lut_n5723 (.I0(x312), .I1(x313), .I2(x314), .O(n5723));
  LUT5 #(.INIT(32'h96696996)) lut_n5724 (.I0(x303), .I1(x304), .I2(x305), .I3(n5716), .I4(n5717), .O(n5724));
  LUT5 #(.INIT(32'hFF969600)) lut_n5725 (.I0(x309), .I1(x310), .I2(x311), .I3(n5723), .I4(n5724), .O(n5725));
  LUT3 #(.INIT(8'h96)) lut_n5726 (.I0(x318), .I1(x319), .I2(x320), .O(n5726));
  LUT5 #(.INIT(32'h96696996)) lut_n5727 (.I0(x309), .I1(x310), .I2(x311), .I3(n5723), .I4(n5724), .O(n5727));
  LUT5 #(.INIT(32'hFF969600)) lut_n5728 (.I0(x315), .I1(x316), .I2(x317), .I3(n5726), .I4(n5727), .O(n5728));
  LUT3 #(.INIT(8'h96)) lut_n5729 (.I0(n5715), .I1(n5718), .I2(n5719), .O(n5729));
  LUT3 #(.INIT(8'hE8)) lut_n5730 (.I0(n5725), .I1(n5728), .I2(n5729), .O(n5730));
  LUT3 #(.INIT(8'h96)) lut_n5731 (.I0(x324), .I1(x325), .I2(x326), .O(n5731));
  LUT5 #(.INIT(32'h96696996)) lut_n5732 (.I0(x315), .I1(x316), .I2(x317), .I3(n5726), .I4(n5727), .O(n5732));
  LUT5 #(.INIT(32'hFF969600)) lut_n5733 (.I0(x321), .I1(x322), .I2(x323), .I3(n5731), .I4(n5732), .O(n5733));
  LUT3 #(.INIT(8'h96)) lut_n5734 (.I0(x330), .I1(x331), .I2(x332), .O(n5734));
  LUT5 #(.INIT(32'h96696996)) lut_n5735 (.I0(x321), .I1(x322), .I2(x323), .I3(n5731), .I4(n5732), .O(n5735));
  LUT5 #(.INIT(32'hFF969600)) lut_n5736 (.I0(x327), .I1(x328), .I2(x329), .I3(n5734), .I4(n5735), .O(n5736));
  LUT3 #(.INIT(8'h96)) lut_n5737 (.I0(n5725), .I1(n5728), .I2(n5729), .O(n5737));
  LUT3 #(.INIT(8'hE8)) lut_n5738 (.I0(n5733), .I1(n5736), .I2(n5737), .O(n5738));
  LUT3 #(.INIT(8'h96)) lut_n5739 (.I0(n5712), .I1(n5720), .I2(n5721), .O(n5739));
  LUT3 #(.INIT(8'hE8)) lut_n5740 (.I0(n5730), .I1(n5738), .I2(n5739), .O(n5740));
  LUT3 #(.INIT(8'h96)) lut_n5741 (.I0(n5684), .I1(n5702), .I2(n5703), .O(n5741));
  LUT3 #(.INIT(8'hE8)) lut_n5742 (.I0(n5722), .I1(n5740), .I2(n5741), .O(n5742));
  LUT3 #(.INIT(8'h96)) lut_n5743 (.I0(n5626), .I1(n5664), .I2(n5665), .O(n5743));
  LUT3 #(.INIT(8'hE8)) lut_n5744 (.I0(n5704), .I1(n5742), .I2(n5743), .O(n5744));
  LUT3 #(.INIT(8'h96)) lut_n5745 (.I0(n5501), .I1(n5579), .I2(n5580), .O(n5745));
  LUT3 #(.INIT(8'hE8)) lut_n5746 (.I0(n5666), .I1(n5744), .I2(n5745), .O(n5746));
  LUT3 #(.INIT(8'h96)) lut_n5747 (.I0(x336), .I1(x337), .I2(x338), .O(n5747));
  LUT5 #(.INIT(32'h96696996)) lut_n5748 (.I0(x327), .I1(x328), .I2(x329), .I3(n5734), .I4(n5735), .O(n5748));
  LUT5 #(.INIT(32'hFF969600)) lut_n5749 (.I0(x333), .I1(x334), .I2(x335), .I3(n5747), .I4(n5748), .O(n5749));
  LUT3 #(.INIT(8'h96)) lut_n5750 (.I0(x342), .I1(x343), .I2(x344), .O(n5750));
  LUT5 #(.INIT(32'h96696996)) lut_n5751 (.I0(x333), .I1(x334), .I2(x335), .I3(n5747), .I4(n5748), .O(n5751));
  LUT5 #(.INIT(32'hFF969600)) lut_n5752 (.I0(x339), .I1(x340), .I2(x341), .I3(n5750), .I4(n5751), .O(n5752));
  LUT3 #(.INIT(8'h96)) lut_n5753 (.I0(n5733), .I1(n5736), .I2(n5737), .O(n5753));
  LUT3 #(.INIT(8'hE8)) lut_n5754 (.I0(n5749), .I1(n5752), .I2(n5753), .O(n5754));
  LUT3 #(.INIT(8'h96)) lut_n5755 (.I0(x348), .I1(x349), .I2(x350), .O(n5755));
  LUT5 #(.INIT(32'h96696996)) lut_n5756 (.I0(x339), .I1(x340), .I2(x341), .I3(n5750), .I4(n5751), .O(n5756));
  LUT5 #(.INIT(32'hFF969600)) lut_n5757 (.I0(x345), .I1(x346), .I2(x347), .I3(n5755), .I4(n5756), .O(n5757));
  LUT3 #(.INIT(8'h96)) lut_n5758 (.I0(x354), .I1(x355), .I2(x356), .O(n5758));
  LUT5 #(.INIT(32'h96696996)) lut_n5759 (.I0(x345), .I1(x346), .I2(x347), .I3(n5755), .I4(n5756), .O(n5759));
  LUT5 #(.INIT(32'hFF969600)) lut_n5760 (.I0(x351), .I1(x352), .I2(x353), .I3(n5758), .I4(n5759), .O(n5760));
  LUT3 #(.INIT(8'h96)) lut_n5761 (.I0(n5749), .I1(n5752), .I2(n5753), .O(n5761));
  LUT3 #(.INIT(8'hE8)) lut_n5762 (.I0(n5757), .I1(n5760), .I2(n5761), .O(n5762));
  LUT3 #(.INIT(8'h96)) lut_n5763 (.I0(n5730), .I1(n5738), .I2(n5739), .O(n5763));
  LUT3 #(.INIT(8'hE8)) lut_n5764 (.I0(n5754), .I1(n5762), .I2(n5763), .O(n5764));
  LUT3 #(.INIT(8'h96)) lut_n5765 (.I0(x360), .I1(x361), .I2(x362), .O(n5765));
  LUT5 #(.INIT(32'h96696996)) lut_n5766 (.I0(x351), .I1(x352), .I2(x353), .I3(n5758), .I4(n5759), .O(n5766));
  LUT5 #(.INIT(32'hFF969600)) lut_n5767 (.I0(x357), .I1(x358), .I2(x359), .I3(n5765), .I4(n5766), .O(n5767));
  LUT3 #(.INIT(8'h96)) lut_n5768 (.I0(x366), .I1(x367), .I2(x368), .O(n5768));
  LUT5 #(.INIT(32'h96696996)) lut_n5769 (.I0(x357), .I1(x358), .I2(x359), .I3(n5765), .I4(n5766), .O(n5769));
  LUT5 #(.INIT(32'hFF969600)) lut_n5770 (.I0(x363), .I1(x364), .I2(x365), .I3(n5768), .I4(n5769), .O(n5770));
  LUT3 #(.INIT(8'h96)) lut_n5771 (.I0(n5757), .I1(n5760), .I2(n5761), .O(n5771));
  LUT3 #(.INIT(8'hE8)) lut_n5772 (.I0(n5767), .I1(n5770), .I2(n5771), .O(n5772));
  LUT3 #(.INIT(8'h96)) lut_n5773 (.I0(x372), .I1(x373), .I2(x374), .O(n5773));
  LUT5 #(.INIT(32'h96696996)) lut_n5774 (.I0(x363), .I1(x364), .I2(x365), .I3(n5768), .I4(n5769), .O(n5774));
  LUT5 #(.INIT(32'hFF969600)) lut_n5775 (.I0(x369), .I1(x370), .I2(x371), .I3(n5773), .I4(n5774), .O(n5775));
  LUT3 #(.INIT(8'h96)) lut_n5776 (.I0(x378), .I1(x379), .I2(x380), .O(n5776));
  LUT5 #(.INIT(32'h96696996)) lut_n5777 (.I0(x369), .I1(x370), .I2(x371), .I3(n5773), .I4(n5774), .O(n5777));
  LUT5 #(.INIT(32'hFF969600)) lut_n5778 (.I0(x375), .I1(x376), .I2(x377), .I3(n5776), .I4(n5777), .O(n5778));
  LUT3 #(.INIT(8'h96)) lut_n5779 (.I0(n5767), .I1(n5770), .I2(n5771), .O(n5779));
  LUT3 #(.INIT(8'hE8)) lut_n5780 (.I0(n5775), .I1(n5778), .I2(n5779), .O(n5780));
  LUT3 #(.INIT(8'h96)) lut_n5781 (.I0(n5754), .I1(n5762), .I2(n5763), .O(n5781));
  LUT3 #(.INIT(8'hE8)) lut_n5782 (.I0(n5772), .I1(n5780), .I2(n5781), .O(n5782));
  LUT3 #(.INIT(8'h96)) lut_n5783 (.I0(n5722), .I1(n5740), .I2(n5741), .O(n5783));
  LUT3 #(.INIT(8'hE8)) lut_n5784 (.I0(n5764), .I1(n5782), .I2(n5783), .O(n5784));
  LUT3 #(.INIT(8'h96)) lut_n5785 (.I0(x384), .I1(x385), .I2(x386), .O(n5785));
  LUT5 #(.INIT(32'h96696996)) lut_n5786 (.I0(x375), .I1(x376), .I2(x377), .I3(n5776), .I4(n5777), .O(n5786));
  LUT5 #(.INIT(32'hFF969600)) lut_n5787 (.I0(x381), .I1(x382), .I2(x383), .I3(n5785), .I4(n5786), .O(n5787));
  LUT3 #(.INIT(8'h96)) lut_n5788 (.I0(x390), .I1(x391), .I2(x392), .O(n5788));
  LUT5 #(.INIT(32'h96696996)) lut_n5789 (.I0(x381), .I1(x382), .I2(x383), .I3(n5785), .I4(n5786), .O(n5789));
  LUT5 #(.INIT(32'hFF969600)) lut_n5790 (.I0(x387), .I1(x388), .I2(x389), .I3(n5788), .I4(n5789), .O(n5790));
  LUT3 #(.INIT(8'h96)) lut_n5791 (.I0(n5775), .I1(n5778), .I2(n5779), .O(n5791));
  LUT3 #(.INIT(8'hE8)) lut_n5792 (.I0(n5787), .I1(n5790), .I2(n5791), .O(n5792));
  LUT3 #(.INIT(8'h96)) lut_n5793 (.I0(x396), .I1(x397), .I2(x398), .O(n5793));
  LUT5 #(.INIT(32'h96696996)) lut_n5794 (.I0(x387), .I1(x388), .I2(x389), .I3(n5788), .I4(n5789), .O(n5794));
  LUT5 #(.INIT(32'hFF969600)) lut_n5795 (.I0(x393), .I1(x394), .I2(x395), .I3(n5793), .I4(n5794), .O(n5795));
  LUT3 #(.INIT(8'h96)) lut_n5796 (.I0(x402), .I1(x403), .I2(x404), .O(n5796));
  LUT5 #(.INIT(32'h96696996)) lut_n5797 (.I0(x393), .I1(x394), .I2(x395), .I3(n5793), .I4(n5794), .O(n5797));
  LUT5 #(.INIT(32'hFF969600)) lut_n5798 (.I0(x399), .I1(x400), .I2(x401), .I3(n5796), .I4(n5797), .O(n5798));
  LUT3 #(.INIT(8'h96)) lut_n5799 (.I0(n5787), .I1(n5790), .I2(n5791), .O(n5799));
  LUT3 #(.INIT(8'hE8)) lut_n5800 (.I0(n5795), .I1(n5798), .I2(n5799), .O(n5800));
  LUT3 #(.INIT(8'h96)) lut_n5801 (.I0(n5772), .I1(n5780), .I2(n5781), .O(n5801));
  LUT3 #(.INIT(8'hE8)) lut_n5802 (.I0(n5792), .I1(n5800), .I2(n5801), .O(n5802));
  LUT3 #(.INIT(8'h96)) lut_n5803 (.I0(x408), .I1(x409), .I2(x410), .O(n5803));
  LUT5 #(.INIT(32'h96696996)) lut_n5804 (.I0(x399), .I1(x400), .I2(x401), .I3(n5796), .I4(n5797), .O(n5804));
  LUT5 #(.INIT(32'hFF969600)) lut_n5805 (.I0(x405), .I1(x406), .I2(x407), .I3(n5803), .I4(n5804), .O(n5805));
  LUT3 #(.INIT(8'h96)) lut_n5806 (.I0(x414), .I1(x415), .I2(x416), .O(n5806));
  LUT5 #(.INIT(32'h96696996)) lut_n5807 (.I0(x405), .I1(x406), .I2(x407), .I3(n5803), .I4(n5804), .O(n5807));
  LUT5 #(.INIT(32'hFF969600)) lut_n5808 (.I0(x411), .I1(x412), .I2(x413), .I3(n5806), .I4(n5807), .O(n5808));
  LUT3 #(.INIT(8'h96)) lut_n5809 (.I0(n5795), .I1(n5798), .I2(n5799), .O(n5809));
  LUT3 #(.INIT(8'hE8)) lut_n5810 (.I0(n5805), .I1(n5808), .I2(n5809), .O(n5810));
  LUT3 #(.INIT(8'h96)) lut_n5811 (.I0(x420), .I1(x421), .I2(x422), .O(n5811));
  LUT5 #(.INIT(32'h96696996)) lut_n5812 (.I0(x411), .I1(x412), .I2(x413), .I3(n5806), .I4(n5807), .O(n5812));
  LUT5 #(.INIT(32'hFF969600)) lut_n5813 (.I0(x417), .I1(x418), .I2(x419), .I3(n5811), .I4(n5812), .O(n5813));
  LUT3 #(.INIT(8'h96)) lut_n5814 (.I0(x426), .I1(x427), .I2(x428), .O(n5814));
  LUT5 #(.INIT(32'h96696996)) lut_n5815 (.I0(x417), .I1(x418), .I2(x419), .I3(n5811), .I4(n5812), .O(n5815));
  LUT5 #(.INIT(32'hFF969600)) lut_n5816 (.I0(x423), .I1(x424), .I2(x425), .I3(n5814), .I4(n5815), .O(n5816));
  LUT3 #(.INIT(8'h96)) lut_n5817 (.I0(n5805), .I1(n5808), .I2(n5809), .O(n5817));
  LUT3 #(.INIT(8'hE8)) lut_n5818 (.I0(n5813), .I1(n5816), .I2(n5817), .O(n5818));
  LUT3 #(.INIT(8'h96)) lut_n5819 (.I0(n5792), .I1(n5800), .I2(n5801), .O(n5819));
  LUT3 #(.INIT(8'hE8)) lut_n5820 (.I0(n5810), .I1(n5818), .I2(n5819), .O(n5820));
  LUT3 #(.INIT(8'h96)) lut_n5821 (.I0(n5764), .I1(n5782), .I2(n5783), .O(n5821));
  LUT3 #(.INIT(8'hE8)) lut_n5822 (.I0(n5802), .I1(n5820), .I2(n5821), .O(n5822));
  LUT3 #(.INIT(8'h96)) lut_n5823 (.I0(n5704), .I1(n5742), .I2(n5743), .O(n5823));
  LUT3 #(.INIT(8'hE8)) lut_n5824 (.I0(n5784), .I1(n5822), .I2(n5823), .O(n5824));
  LUT3 #(.INIT(8'h96)) lut_n5825 (.I0(x432), .I1(x433), .I2(x434), .O(n5825));
  LUT5 #(.INIT(32'h96696996)) lut_n5826 (.I0(x423), .I1(x424), .I2(x425), .I3(n5814), .I4(n5815), .O(n5826));
  LUT5 #(.INIT(32'hFF969600)) lut_n5827 (.I0(x429), .I1(x430), .I2(x431), .I3(n5825), .I4(n5826), .O(n5827));
  LUT3 #(.INIT(8'h96)) lut_n5828 (.I0(x438), .I1(x439), .I2(x440), .O(n5828));
  LUT5 #(.INIT(32'h96696996)) lut_n5829 (.I0(x429), .I1(x430), .I2(x431), .I3(n5825), .I4(n5826), .O(n5829));
  LUT5 #(.INIT(32'hFF969600)) lut_n5830 (.I0(x435), .I1(x436), .I2(x437), .I3(n5828), .I4(n5829), .O(n5830));
  LUT3 #(.INIT(8'h96)) lut_n5831 (.I0(n5813), .I1(n5816), .I2(n5817), .O(n5831));
  LUT3 #(.INIT(8'hE8)) lut_n5832 (.I0(n5827), .I1(n5830), .I2(n5831), .O(n5832));
  LUT3 #(.INIT(8'h96)) lut_n5833 (.I0(x444), .I1(x445), .I2(x446), .O(n5833));
  LUT5 #(.INIT(32'h96696996)) lut_n5834 (.I0(x435), .I1(x436), .I2(x437), .I3(n5828), .I4(n5829), .O(n5834));
  LUT5 #(.INIT(32'hFF969600)) lut_n5835 (.I0(x441), .I1(x442), .I2(x443), .I3(n5833), .I4(n5834), .O(n5835));
  LUT3 #(.INIT(8'h96)) lut_n5836 (.I0(x450), .I1(x451), .I2(x452), .O(n5836));
  LUT5 #(.INIT(32'h96696996)) lut_n5837 (.I0(x441), .I1(x442), .I2(x443), .I3(n5833), .I4(n5834), .O(n5837));
  LUT5 #(.INIT(32'hFF969600)) lut_n5838 (.I0(x447), .I1(x448), .I2(x449), .I3(n5836), .I4(n5837), .O(n5838));
  LUT3 #(.INIT(8'h96)) lut_n5839 (.I0(n5827), .I1(n5830), .I2(n5831), .O(n5839));
  LUT3 #(.INIT(8'hE8)) lut_n5840 (.I0(n5835), .I1(n5838), .I2(n5839), .O(n5840));
  LUT3 #(.INIT(8'h96)) lut_n5841 (.I0(n5810), .I1(n5818), .I2(n5819), .O(n5841));
  LUT3 #(.INIT(8'hE8)) lut_n5842 (.I0(n5832), .I1(n5840), .I2(n5841), .O(n5842));
  LUT3 #(.INIT(8'h96)) lut_n5843 (.I0(x456), .I1(x457), .I2(x458), .O(n5843));
  LUT5 #(.INIT(32'h96696996)) lut_n5844 (.I0(x447), .I1(x448), .I2(x449), .I3(n5836), .I4(n5837), .O(n5844));
  LUT5 #(.INIT(32'hFF969600)) lut_n5845 (.I0(x453), .I1(x454), .I2(x455), .I3(n5843), .I4(n5844), .O(n5845));
  LUT3 #(.INIT(8'h96)) lut_n5846 (.I0(x462), .I1(x463), .I2(x464), .O(n5846));
  LUT5 #(.INIT(32'h96696996)) lut_n5847 (.I0(x453), .I1(x454), .I2(x455), .I3(n5843), .I4(n5844), .O(n5847));
  LUT5 #(.INIT(32'hFF969600)) lut_n5848 (.I0(x459), .I1(x460), .I2(x461), .I3(n5846), .I4(n5847), .O(n5848));
  LUT3 #(.INIT(8'h96)) lut_n5849 (.I0(n5835), .I1(n5838), .I2(n5839), .O(n5849));
  LUT3 #(.INIT(8'hE8)) lut_n5850 (.I0(n5845), .I1(n5848), .I2(n5849), .O(n5850));
  LUT3 #(.INIT(8'h96)) lut_n5851 (.I0(x468), .I1(x469), .I2(x470), .O(n5851));
  LUT5 #(.INIT(32'h96696996)) lut_n5852 (.I0(x459), .I1(x460), .I2(x461), .I3(n5846), .I4(n5847), .O(n5852));
  LUT5 #(.INIT(32'hFF969600)) lut_n5853 (.I0(x465), .I1(x466), .I2(x467), .I3(n5851), .I4(n5852), .O(n5853));
  LUT3 #(.INIT(8'h96)) lut_n5854 (.I0(x474), .I1(x475), .I2(x476), .O(n5854));
  LUT5 #(.INIT(32'h96696996)) lut_n5855 (.I0(x465), .I1(x466), .I2(x467), .I3(n5851), .I4(n5852), .O(n5855));
  LUT5 #(.INIT(32'hFF969600)) lut_n5856 (.I0(x471), .I1(x472), .I2(x473), .I3(n5854), .I4(n5855), .O(n5856));
  LUT3 #(.INIT(8'h96)) lut_n5857 (.I0(n5845), .I1(n5848), .I2(n5849), .O(n5857));
  LUT3 #(.INIT(8'hE8)) lut_n5858 (.I0(n5853), .I1(n5856), .I2(n5857), .O(n5858));
  LUT3 #(.INIT(8'h96)) lut_n5859 (.I0(n5832), .I1(n5840), .I2(n5841), .O(n5859));
  LUT3 #(.INIT(8'hE8)) lut_n5860 (.I0(n5850), .I1(n5858), .I2(n5859), .O(n5860));
  LUT3 #(.INIT(8'h96)) lut_n5861 (.I0(n5802), .I1(n5820), .I2(n5821), .O(n5861));
  LUT3 #(.INIT(8'hE8)) lut_n5862 (.I0(n5842), .I1(n5860), .I2(n5861), .O(n5862));
  LUT3 #(.INIT(8'h96)) lut_n5863 (.I0(x480), .I1(x481), .I2(x482), .O(n5863));
  LUT5 #(.INIT(32'h96696996)) lut_n5864 (.I0(x471), .I1(x472), .I2(x473), .I3(n5854), .I4(n5855), .O(n5864));
  LUT5 #(.INIT(32'hFF969600)) lut_n5865 (.I0(x477), .I1(x478), .I2(x479), .I3(n5863), .I4(n5864), .O(n5865));
  LUT3 #(.INIT(8'h96)) lut_n5866 (.I0(x486), .I1(x487), .I2(x488), .O(n5866));
  LUT5 #(.INIT(32'h96696996)) lut_n5867 (.I0(x477), .I1(x478), .I2(x479), .I3(n5863), .I4(n5864), .O(n5867));
  LUT5 #(.INIT(32'hFF969600)) lut_n5868 (.I0(x483), .I1(x484), .I2(x485), .I3(n5866), .I4(n5867), .O(n5868));
  LUT3 #(.INIT(8'h96)) lut_n5869 (.I0(n5853), .I1(n5856), .I2(n5857), .O(n5869));
  LUT3 #(.INIT(8'hE8)) lut_n5870 (.I0(n5865), .I1(n5868), .I2(n5869), .O(n5870));
  LUT3 #(.INIT(8'h96)) lut_n5871 (.I0(x492), .I1(x493), .I2(x494), .O(n5871));
  LUT5 #(.INIT(32'h96696996)) lut_n5872 (.I0(x483), .I1(x484), .I2(x485), .I3(n5866), .I4(n5867), .O(n5872));
  LUT5 #(.INIT(32'hFF969600)) lut_n5873 (.I0(x489), .I1(x490), .I2(x491), .I3(n5871), .I4(n5872), .O(n5873));
  LUT3 #(.INIT(8'h96)) lut_n5874 (.I0(x498), .I1(x499), .I2(x500), .O(n5874));
  LUT5 #(.INIT(32'h96696996)) lut_n5875 (.I0(x489), .I1(x490), .I2(x491), .I3(n5871), .I4(n5872), .O(n5875));
  LUT5 #(.INIT(32'hFF969600)) lut_n5876 (.I0(x495), .I1(x496), .I2(x497), .I3(n5874), .I4(n5875), .O(n5876));
  LUT3 #(.INIT(8'h96)) lut_n5877 (.I0(n5865), .I1(n5868), .I2(n5869), .O(n5877));
  LUT3 #(.INIT(8'hE8)) lut_n5878 (.I0(n5873), .I1(n5876), .I2(n5877), .O(n5878));
  LUT3 #(.INIT(8'h96)) lut_n5879 (.I0(n5850), .I1(n5858), .I2(n5859), .O(n5879));
  LUT3 #(.INIT(8'hE8)) lut_n5880 (.I0(n5870), .I1(n5878), .I2(n5879), .O(n5880));
  LUT3 #(.INIT(8'h96)) lut_n5881 (.I0(x504), .I1(x505), .I2(x506), .O(n5881));
  LUT5 #(.INIT(32'h96696996)) lut_n5882 (.I0(x495), .I1(x496), .I2(x497), .I3(n5874), .I4(n5875), .O(n5882));
  LUT5 #(.INIT(32'hFF969600)) lut_n5883 (.I0(x501), .I1(x502), .I2(x503), .I3(n5881), .I4(n5882), .O(n5883));
  LUT3 #(.INIT(8'h96)) lut_n5884 (.I0(x510), .I1(x511), .I2(x512), .O(n5884));
  LUT5 #(.INIT(32'h96696996)) lut_n5885 (.I0(x501), .I1(x502), .I2(x503), .I3(n5881), .I4(n5882), .O(n5885));
  LUT5 #(.INIT(32'hFF969600)) lut_n5886 (.I0(x507), .I1(x508), .I2(x509), .I3(n5884), .I4(n5885), .O(n5886));
  LUT3 #(.INIT(8'h96)) lut_n5887 (.I0(n5873), .I1(n5876), .I2(n5877), .O(n5887));
  LUT3 #(.INIT(8'hE8)) lut_n5888 (.I0(n5883), .I1(n5886), .I2(n5887), .O(n5888));
  LUT3 #(.INIT(8'h96)) lut_n5889 (.I0(x516), .I1(x517), .I2(x518), .O(n5889));
  LUT5 #(.INIT(32'h96696996)) lut_n5890 (.I0(x507), .I1(x508), .I2(x509), .I3(n5884), .I4(n5885), .O(n5890));
  LUT5 #(.INIT(32'hFF969600)) lut_n5891 (.I0(x513), .I1(x514), .I2(x515), .I3(n5889), .I4(n5890), .O(n5891));
  LUT3 #(.INIT(8'h96)) lut_n5892 (.I0(x522), .I1(x523), .I2(x524), .O(n5892));
  LUT5 #(.INIT(32'h96696996)) lut_n5893 (.I0(x513), .I1(x514), .I2(x515), .I3(n5889), .I4(n5890), .O(n5893));
  LUT5 #(.INIT(32'hFF969600)) lut_n5894 (.I0(x519), .I1(x520), .I2(x521), .I3(n5892), .I4(n5893), .O(n5894));
  LUT3 #(.INIT(8'h96)) lut_n5895 (.I0(n5883), .I1(n5886), .I2(n5887), .O(n5895));
  LUT3 #(.INIT(8'hE8)) lut_n5896 (.I0(n5891), .I1(n5894), .I2(n5895), .O(n5896));
  LUT3 #(.INIT(8'h96)) lut_n5897 (.I0(n5870), .I1(n5878), .I2(n5879), .O(n5897));
  LUT3 #(.INIT(8'hE8)) lut_n5898 (.I0(n5888), .I1(n5896), .I2(n5897), .O(n5898));
  LUT3 #(.INIT(8'h96)) lut_n5899 (.I0(n5842), .I1(n5860), .I2(n5861), .O(n5899));
  LUT3 #(.INIT(8'hE8)) lut_n5900 (.I0(n5880), .I1(n5898), .I2(n5899), .O(n5900));
  LUT3 #(.INIT(8'h96)) lut_n5901 (.I0(n5784), .I1(n5822), .I2(n5823), .O(n5901));
  LUT3 #(.INIT(8'hE8)) lut_n5902 (.I0(n5862), .I1(n5900), .I2(n5901), .O(n5902));
  LUT3 #(.INIT(8'h96)) lut_n5903 (.I0(n5666), .I1(n5744), .I2(n5745), .O(n5903));
  LUT3 #(.INIT(8'hE8)) lut_n5904 (.I0(n5824), .I1(n5902), .I2(n5903), .O(n5904));
  LUT3 #(.INIT(8'h96)) lut_n5905 (.I0(n5446), .I1(n5581), .I2(n5582), .O(n5905));
  LUT3 #(.INIT(8'hE8)) lut_n5906 (.I0(n5746), .I1(n5904), .I2(n5905), .O(n5906));
  LUT3 #(.INIT(8'h96)) lut_n5907 (.I0(x528), .I1(x529), .I2(x530), .O(n5907));
  LUT5 #(.INIT(32'h96696996)) lut_n5908 (.I0(x519), .I1(x520), .I2(x521), .I3(n5892), .I4(n5893), .O(n5908));
  LUT5 #(.INIT(32'hFF969600)) lut_n5909 (.I0(x525), .I1(x526), .I2(x527), .I3(n5907), .I4(n5908), .O(n5909));
  LUT3 #(.INIT(8'h96)) lut_n5910 (.I0(x534), .I1(x535), .I2(x536), .O(n5910));
  LUT5 #(.INIT(32'h96696996)) lut_n5911 (.I0(x525), .I1(x526), .I2(x527), .I3(n5907), .I4(n5908), .O(n5911));
  LUT5 #(.INIT(32'hFF969600)) lut_n5912 (.I0(x531), .I1(x532), .I2(x533), .I3(n5910), .I4(n5911), .O(n5912));
  LUT3 #(.INIT(8'h96)) lut_n5913 (.I0(n5891), .I1(n5894), .I2(n5895), .O(n5913));
  LUT3 #(.INIT(8'hE8)) lut_n5914 (.I0(n5909), .I1(n5912), .I2(n5913), .O(n5914));
  LUT3 #(.INIT(8'h96)) lut_n5915 (.I0(x540), .I1(x541), .I2(x542), .O(n5915));
  LUT5 #(.INIT(32'h96696996)) lut_n5916 (.I0(x531), .I1(x532), .I2(x533), .I3(n5910), .I4(n5911), .O(n5916));
  LUT5 #(.INIT(32'hFF969600)) lut_n5917 (.I0(x537), .I1(x538), .I2(x539), .I3(n5915), .I4(n5916), .O(n5917));
  LUT3 #(.INIT(8'h96)) lut_n5918 (.I0(x546), .I1(x547), .I2(x548), .O(n5918));
  LUT5 #(.INIT(32'h96696996)) lut_n5919 (.I0(x537), .I1(x538), .I2(x539), .I3(n5915), .I4(n5916), .O(n5919));
  LUT5 #(.INIT(32'hFF969600)) lut_n5920 (.I0(x543), .I1(x544), .I2(x545), .I3(n5918), .I4(n5919), .O(n5920));
  LUT3 #(.INIT(8'h96)) lut_n5921 (.I0(n5909), .I1(n5912), .I2(n5913), .O(n5921));
  LUT3 #(.INIT(8'hE8)) lut_n5922 (.I0(n5917), .I1(n5920), .I2(n5921), .O(n5922));
  LUT3 #(.INIT(8'h96)) lut_n5923 (.I0(n5888), .I1(n5896), .I2(n5897), .O(n5923));
  LUT3 #(.INIT(8'hE8)) lut_n5924 (.I0(n5914), .I1(n5922), .I2(n5923), .O(n5924));
  LUT3 #(.INIT(8'h96)) lut_n5925 (.I0(x552), .I1(x553), .I2(x554), .O(n5925));
  LUT5 #(.INIT(32'h96696996)) lut_n5926 (.I0(x543), .I1(x544), .I2(x545), .I3(n5918), .I4(n5919), .O(n5926));
  LUT5 #(.INIT(32'hFF969600)) lut_n5927 (.I0(x549), .I1(x550), .I2(x551), .I3(n5925), .I4(n5926), .O(n5927));
  LUT3 #(.INIT(8'h96)) lut_n5928 (.I0(x558), .I1(x559), .I2(x560), .O(n5928));
  LUT5 #(.INIT(32'h96696996)) lut_n5929 (.I0(x549), .I1(x550), .I2(x551), .I3(n5925), .I4(n5926), .O(n5929));
  LUT5 #(.INIT(32'hFF969600)) lut_n5930 (.I0(x555), .I1(x556), .I2(x557), .I3(n5928), .I4(n5929), .O(n5930));
  LUT3 #(.INIT(8'h96)) lut_n5931 (.I0(n5917), .I1(n5920), .I2(n5921), .O(n5931));
  LUT3 #(.INIT(8'hE8)) lut_n5932 (.I0(n5927), .I1(n5930), .I2(n5931), .O(n5932));
  LUT3 #(.INIT(8'h96)) lut_n5933 (.I0(x564), .I1(x565), .I2(x566), .O(n5933));
  LUT5 #(.INIT(32'h96696996)) lut_n5934 (.I0(x555), .I1(x556), .I2(x557), .I3(n5928), .I4(n5929), .O(n5934));
  LUT5 #(.INIT(32'hFF969600)) lut_n5935 (.I0(x561), .I1(x562), .I2(x563), .I3(n5933), .I4(n5934), .O(n5935));
  LUT3 #(.INIT(8'h96)) lut_n5936 (.I0(x570), .I1(x571), .I2(x572), .O(n5936));
  LUT5 #(.INIT(32'h96696996)) lut_n5937 (.I0(x561), .I1(x562), .I2(x563), .I3(n5933), .I4(n5934), .O(n5937));
  LUT5 #(.INIT(32'hFF969600)) lut_n5938 (.I0(x567), .I1(x568), .I2(x569), .I3(n5936), .I4(n5937), .O(n5938));
  LUT3 #(.INIT(8'h96)) lut_n5939 (.I0(n5927), .I1(n5930), .I2(n5931), .O(n5939));
  LUT3 #(.INIT(8'hE8)) lut_n5940 (.I0(n5935), .I1(n5938), .I2(n5939), .O(n5940));
  LUT3 #(.INIT(8'h96)) lut_n5941 (.I0(n5914), .I1(n5922), .I2(n5923), .O(n5941));
  LUT3 #(.INIT(8'hE8)) lut_n5942 (.I0(n5932), .I1(n5940), .I2(n5941), .O(n5942));
  LUT3 #(.INIT(8'h96)) lut_n5943 (.I0(n5880), .I1(n5898), .I2(n5899), .O(n5943));
  LUT3 #(.INIT(8'hE8)) lut_n5944 (.I0(n5924), .I1(n5942), .I2(n5943), .O(n5944));
  LUT3 #(.INIT(8'h96)) lut_n5945 (.I0(x576), .I1(x577), .I2(x578), .O(n5945));
  LUT5 #(.INIT(32'h96696996)) lut_n5946 (.I0(x567), .I1(x568), .I2(x569), .I3(n5936), .I4(n5937), .O(n5946));
  LUT5 #(.INIT(32'hFF969600)) lut_n5947 (.I0(x573), .I1(x574), .I2(x575), .I3(n5945), .I4(n5946), .O(n5947));
  LUT3 #(.INIT(8'h96)) lut_n5948 (.I0(x582), .I1(x583), .I2(x584), .O(n5948));
  LUT5 #(.INIT(32'h96696996)) lut_n5949 (.I0(x573), .I1(x574), .I2(x575), .I3(n5945), .I4(n5946), .O(n5949));
  LUT5 #(.INIT(32'hFF969600)) lut_n5950 (.I0(x579), .I1(x580), .I2(x581), .I3(n5948), .I4(n5949), .O(n5950));
  LUT3 #(.INIT(8'h96)) lut_n5951 (.I0(n5935), .I1(n5938), .I2(n5939), .O(n5951));
  LUT3 #(.INIT(8'hE8)) lut_n5952 (.I0(n5947), .I1(n5950), .I2(n5951), .O(n5952));
  LUT3 #(.INIT(8'h96)) lut_n5953 (.I0(x588), .I1(x589), .I2(x590), .O(n5953));
  LUT5 #(.INIT(32'h96696996)) lut_n5954 (.I0(x579), .I1(x580), .I2(x581), .I3(n5948), .I4(n5949), .O(n5954));
  LUT5 #(.INIT(32'hFF969600)) lut_n5955 (.I0(x585), .I1(x586), .I2(x587), .I3(n5953), .I4(n5954), .O(n5955));
  LUT3 #(.INIT(8'h96)) lut_n5956 (.I0(x594), .I1(x595), .I2(x596), .O(n5956));
  LUT5 #(.INIT(32'h96696996)) lut_n5957 (.I0(x585), .I1(x586), .I2(x587), .I3(n5953), .I4(n5954), .O(n5957));
  LUT5 #(.INIT(32'hFF969600)) lut_n5958 (.I0(x591), .I1(x592), .I2(x593), .I3(n5956), .I4(n5957), .O(n5958));
  LUT3 #(.INIT(8'h96)) lut_n5959 (.I0(n5947), .I1(n5950), .I2(n5951), .O(n5959));
  LUT3 #(.INIT(8'hE8)) lut_n5960 (.I0(n5955), .I1(n5958), .I2(n5959), .O(n5960));
  LUT3 #(.INIT(8'h96)) lut_n5961 (.I0(n5932), .I1(n5940), .I2(n5941), .O(n5961));
  LUT3 #(.INIT(8'hE8)) lut_n5962 (.I0(n5952), .I1(n5960), .I2(n5961), .O(n5962));
  LUT3 #(.INIT(8'h96)) lut_n5963 (.I0(x600), .I1(x601), .I2(x602), .O(n5963));
  LUT5 #(.INIT(32'h96696996)) lut_n5964 (.I0(x591), .I1(x592), .I2(x593), .I3(n5956), .I4(n5957), .O(n5964));
  LUT5 #(.INIT(32'hFF969600)) lut_n5965 (.I0(x597), .I1(x598), .I2(x599), .I3(n5963), .I4(n5964), .O(n5965));
  LUT3 #(.INIT(8'h96)) lut_n5966 (.I0(x606), .I1(x607), .I2(x608), .O(n5966));
  LUT5 #(.INIT(32'h96696996)) lut_n5967 (.I0(x597), .I1(x598), .I2(x599), .I3(n5963), .I4(n5964), .O(n5967));
  LUT5 #(.INIT(32'hFF969600)) lut_n5968 (.I0(x603), .I1(x604), .I2(x605), .I3(n5966), .I4(n5967), .O(n5968));
  LUT3 #(.INIT(8'h96)) lut_n5969 (.I0(n5955), .I1(n5958), .I2(n5959), .O(n5969));
  LUT3 #(.INIT(8'hE8)) lut_n5970 (.I0(n5965), .I1(n5968), .I2(n5969), .O(n5970));
  LUT3 #(.INIT(8'h96)) lut_n5971 (.I0(x612), .I1(x613), .I2(x614), .O(n5971));
  LUT5 #(.INIT(32'h96696996)) lut_n5972 (.I0(x603), .I1(x604), .I2(x605), .I3(n5966), .I4(n5967), .O(n5972));
  LUT5 #(.INIT(32'hFF969600)) lut_n5973 (.I0(x609), .I1(x610), .I2(x611), .I3(n5971), .I4(n5972), .O(n5973));
  LUT3 #(.INIT(8'h96)) lut_n5974 (.I0(x618), .I1(x619), .I2(x620), .O(n5974));
  LUT5 #(.INIT(32'h96696996)) lut_n5975 (.I0(x609), .I1(x610), .I2(x611), .I3(n5971), .I4(n5972), .O(n5975));
  LUT5 #(.INIT(32'hFF969600)) lut_n5976 (.I0(x615), .I1(x616), .I2(x617), .I3(n5974), .I4(n5975), .O(n5976));
  LUT3 #(.INIT(8'h96)) lut_n5977 (.I0(n5965), .I1(n5968), .I2(n5969), .O(n5977));
  LUT3 #(.INIT(8'hE8)) lut_n5978 (.I0(n5973), .I1(n5976), .I2(n5977), .O(n5978));
  LUT3 #(.INIT(8'h96)) lut_n5979 (.I0(n5952), .I1(n5960), .I2(n5961), .O(n5979));
  LUT3 #(.INIT(8'hE8)) lut_n5980 (.I0(n5970), .I1(n5978), .I2(n5979), .O(n5980));
  LUT3 #(.INIT(8'h96)) lut_n5981 (.I0(n5924), .I1(n5942), .I2(n5943), .O(n5981));
  LUT3 #(.INIT(8'hE8)) lut_n5982 (.I0(n5962), .I1(n5980), .I2(n5981), .O(n5982));
  LUT3 #(.INIT(8'h96)) lut_n5983 (.I0(n5862), .I1(n5900), .I2(n5901), .O(n5983));
  LUT3 #(.INIT(8'hE8)) lut_n5984 (.I0(n5944), .I1(n5982), .I2(n5983), .O(n5984));
  LUT3 #(.INIT(8'h96)) lut_n5985 (.I0(x624), .I1(x625), .I2(x626), .O(n5985));
  LUT5 #(.INIT(32'h96696996)) lut_n5986 (.I0(x615), .I1(x616), .I2(x617), .I3(n5974), .I4(n5975), .O(n5986));
  LUT5 #(.INIT(32'hFF969600)) lut_n5987 (.I0(x621), .I1(x622), .I2(x623), .I3(n5985), .I4(n5986), .O(n5987));
  LUT3 #(.INIT(8'h96)) lut_n5988 (.I0(x630), .I1(x631), .I2(x632), .O(n5988));
  LUT5 #(.INIT(32'h96696996)) lut_n5989 (.I0(x621), .I1(x622), .I2(x623), .I3(n5985), .I4(n5986), .O(n5989));
  LUT5 #(.INIT(32'hFF969600)) lut_n5990 (.I0(x627), .I1(x628), .I2(x629), .I3(n5988), .I4(n5989), .O(n5990));
  LUT3 #(.INIT(8'h96)) lut_n5991 (.I0(n5973), .I1(n5976), .I2(n5977), .O(n5991));
  LUT3 #(.INIT(8'hE8)) lut_n5992 (.I0(n5987), .I1(n5990), .I2(n5991), .O(n5992));
  LUT3 #(.INIT(8'h96)) lut_n5993 (.I0(x636), .I1(x637), .I2(x638), .O(n5993));
  LUT5 #(.INIT(32'h96696996)) lut_n5994 (.I0(x627), .I1(x628), .I2(x629), .I3(n5988), .I4(n5989), .O(n5994));
  LUT5 #(.INIT(32'hFF969600)) lut_n5995 (.I0(x633), .I1(x634), .I2(x635), .I3(n5993), .I4(n5994), .O(n5995));
  LUT3 #(.INIT(8'h96)) lut_n5996 (.I0(x642), .I1(x643), .I2(x644), .O(n5996));
  LUT5 #(.INIT(32'h96696996)) lut_n5997 (.I0(x633), .I1(x634), .I2(x635), .I3(n5993), .I4(n5994), .O(n5997));
  LUT5 #(.INIT(32'hFF969600)) lut_n5998 (.I0(x639), .I1(x640), .I2(x641), .I3(n5996), .I4(n5997), .O(n5998));
  LUT3 #(.INIT(8'h96)) lut_n5999 (.I0(n5987), .I1(n5990), .I2(n5991), .O(n5999));
  LUT3 #(.INIT(8'hE8)) lut_n6000 (.I0(n5995), .I1(n5998), .I2(n5999), .O(n6000));
  LUT3 #(.INIT(8'h96)) lut_n6001 (.I0(n5970), .I1(n5978), .I2(n5979), .O(n6001));
  LUT3 #(.INIT(8'hE8)) lut_n6002 (.I0(n5992), .I1(n6000), .I2(n6001), .O(n6002));
  LUT3 #(.INIT(8'h96)) lut_n6003 (.I0(x648), .I1(x649), .I2(x650), .O(n6003));
  LUT5 #(.INIT(32'h96696996)) lut_n6004 (.I0(x639), .I1(x640), .I2(x641), .I3(n5996), .I4(n5997), .O(n6004));
  LUT5 #(.INIT(32'hFF969600)) lut_n6005 (.I0(x645), .I1(x646), .I2(x647), .I3(n6003), .I4(n6004), .O(n6005));
  LUT3 #(.INIT(8'h96)) lut_n6006 (.I0(x654), .I1(x655), .I2(x656), .O(n6006));
  LUT5 #(.INIT(32'h96696996)) lut_n6007 (.I0(x645), .I1(x646), .I2(x647), .I3(n6003), .I4(n6004), .O(n6007));
  LUT5 #(.INIT(32'hFF969600)) lut_n6008 (.I0(x651), .I1(x652), .I2(x653), .I3(n6006), .I4(n6007), .O(n6008));
  LUT3 #(.INIT(8'h96)) lut_n6009 (.I0(n5995), .I1(n5998), .I2(n5999), .O(n6009));
  LUT3 #(.INIT(8'hE8)) lut_n6010 (.I0(n6005), .I1(n6008), .I2(n6009), .O(n6010));
  LUT3 #(.INIT(8'h96)) lut_n6011 (.I0(x660), .I1(x661), .I2(x662), .O(n6011));
  LUT5 #(.INIT(32'h96696996)) lut_n6012 (.I0(x651), .I1(x652), .I2(x653), .I3(n6006), .I4(n6007), .O(n6012));
  LUT5 #(.INIT(32'hFF969600)) lut_n6013 (.I0(x657), .I1(x658), .I2(x659), .I3(n6011), .I4(n6012), .O(n6013));
  LUT3 #(.INIT(8'h96)) lut_n6014 (.I0(x666), .I1(x667), .I2(x668), .O(n6014));
  LUT5 #(.INIT(32'h96696996)) lut_n6015 (.I0(x657), .I1(x658), .I2(x659), .I3(n6011), .I4(n6012), .O(n6015));
  LUT5 #(.INIT(32'hFF969600)) lut_n6016 (.I0(x663), .I1(x664), .I2(x665), .I3(n6014), .I4(n6015), .O(n6016));
  LUT3 #(.INIT(8'h96)) lut_n6017 (.I0(n6005), .I1(n6008), .I2(n6009), .O(n6017));
  LUT3 #(.INIT(8'hE8)) lut_n6018 (.I0(n6013), .I1(n6016), .I2(n6017), .O(n6018));
  LUT3 #(.INIT(8'h96)) lut_n6019 (.I0(n5992), .I1(n6000), .I2(n6001), .O(n6019));
  LUT3 #(.INIT(8'hE8)) lut_n6020 (.I0(n6010), .I1(n6018), .I2(n6019), .O(n6020));
  LUT3 #(.INIT(8'h96)) lut_n6021 (.I0(n5962), .I1(n5980), .I2(n5981), .O(n6021));
  LUT3 #(.INIT(8'hE8)) lut_n6022 (.I0(n6002), .I1(n6020), .I2(n6021), .O(n6022));
  LUT3 #(.INIT(8'h96)) lut_n6023 (.I0(x672), .I1(x673), .I2(x674), .O(n6023));
  LUT5 #(.INIT(32'h96696996)) lut_n6024 (.I0(x663), .I1(x664), .I2(x665), .I3(n6014), .I4(n6015), .O(n6024));
  LUT5 #(.INIT(32'hFF969600)) lut_n6025 (.I0(x669), .I1(x670), .I2(x671), .I3(n6023), .I4(n6024), .O(n6025));
  LUT3 #(.INIT(8'h96)) lut_n6026 (.I0(x678), .I1(x679), .I2(x680), .O(n6026));
  LUT5 #(.INIT(32'h96696996)) lut_n6027 (.I0(x669), .I1(x670), .I2(x671), .I3(n6023), .I4(n6024), .O(n6027));
  LUT5 #(.INIT(32'hFF969600)) lut_n6028 (.I0(x675), .I1(x676), .I2(x677), .I3(n6026), .I4(n6027), .O(n6028));
  LUT3 #(.INIT(8'h96)) lut_n6029 (.I0(n6013), .I1(n6016), .I2(n6017), .O(n6029));
  LUT3 #(.INIT(8'hE8)) lut_n6030 (.I0(n6025), .I1(n6028), .I2(n6029), .O(n6030));
  LUT3 #(.INIT(8'h96)) lut_n6031 (.I0(x684), .I1(x685), .I2(x686), .O(n6031));
  LUT5 #(.INIT(32'h96696996)) lut_n6032 (.I0(x675), .I1(x676), .I2(x677), .I3(n6026), .I4(n6027), .O(n6032));
  LUT5 #(.INIT(32'hFF969600)) lut_n6033 (.I0(x681), .I1(x682), .I2(x683), .I3(n6031), .I4(n6032), .O(n6033));
  LUT3 #(.INIT(8'h96)) lut_n6034 (.I0(x690), .I1(x691), .I2(x692), .O(n6034));
  LUT5 #(.INIT(32'h96696996)) lut_n6035 (.I0(x681), .I1(x682), .I2(x683), .I3(n6031), .I4(n6032), .O(n6035));
  LUT5 #(.INIT(32'hFF969600)) lut_n6036 (.I0(x687), .I1(x688), .I2(x689), .I3(n6034), .I4(n6035), .O(n6036));
  LUT3 #(.INIT(8'h96)) lut_n6037 (.I0(n6025), .I1(n6028), .I2(n6029), .O(n6037));
  LUT3 #(.INIT(8'hE8)) lut_n6038 (.I0(n6033), .I1(n6036), .I2(n6037), .O(n6038));
  LUT3 #(.INIT(8'h96)) lut_n6039 (.I0(n6010), .I1(n6018), .I2(n6019), .O(n6039));
  LUT3 #(.INIT(8'hE8)) lut_n6040 (.I0(n6030), .I1(n6038), .I2(n6039), .O(n6040));
  LUT3 #(.INIT(8'h96)) lut_n6041 (.I0(x696), .I1(x697), .I2(x698), .O(n6041));
  LUT5 #(.INIT(32'h96696996)) lut_n6042 (.I0(x687), .I1(x688), .I2(x689), .I3(n6034), .I4(n6035), .O(n6042));
  LUT5 #(.INIT(32'hFF969600)) lut_n6043 (.I0(x693), .I1(x694), .I2(x695), .I3(n6041), .I4(n6042), .O(n6043));
  LUT3 #(.INIT(8'h96)) lut_n6044 (.I0(x702), .I1(x703), .I2(x704), .O(n6044));
  LUT5 #(.INIT(32'h96696996)) lut_n6045 (.I0(x693), .I1(x694), .I2(x695), .I3(n6041), .I4(n6042), .O(n6045));
  LUT5 #(.INIT(32'hFF969600)) lut_n6046 (.I0(x699), .I1(x700), .I2(x701), .I3(n6044), .I4(n6045), .O(n6046));
  LUT3 #(.INIT(8'h96)) lut_n6047 (.I0(n6033), .I1(n6036), .I2(n6037), .O(n6047));
  LUT3 #(.INIT(8'hE8)) lut_n6048 (.I0(n6043), .I1(n6046), .I2(n6047), .O(n6048));
  LUT3 #(.INIT(8'h96)) lut_n6049 (.I0(x708), .I1(x709), .I2(x710), .O(n6049));
  LUT5 #(.INIT(32'h96696996)) lut_n6050 (.I0(x699), .I1(x700), .I2(x701), .I3(n6044), .I4(n6045), .O(n6050));
  LUT5 #(.INIT(32'hFF969600)) lut_n6051 (.I0(x705), .I1(x706), .I2(x707), .I3(n6049), .I4(n6050), .O(n6051));
  LUT3 #(.INIT(8'h96)) lut_n6052 (.I0(x714), .I1(x715), .I2(x716), .O(n6052));
  LUT5 #(.INIT(32'h96696996)) lut_n6053 (.I0(x705), .I1(x706), .I2(x707), .I3(n6049), .I4(n6050), .O(n6053));
  LUT5 #(.INIT(32'hFF969600)) lut_n6054 (.I0(x711), .I1(x712), .I2(x713), .I3(n6052), .I4(n6053), .O(n6054));
  LUT3 #(.INIT(8'h96)) lut_n6055 (.I0(n6043), .I1(n6046), .I2(n6047), .O(n6055));
  LUT3 #(.INIT(8'hE8)) lut_n6056 (.I0(n6051), .I1(n6054), .I2(n6055), .O(n6056));
  LUT3 #(.INIT(8'h96)) lut_n6057 (.I0(n6030), .I1(n6038), .I2(n6039), .O(n6057));
  LUT3 #(.INIT(8'hE8)) lut_n6058 (.I0(n6048), .I1(n6056), .I2(n6057), .O(n6058));
  LUT3 #(.INIT(8'h96)) lut_n6059 (.I0(n6002), .I1(n6020), .I2(n6021), .O(n6059));
  LUT3 #(.INIT(8'hE8)) lut_n6060 (.I0(n6040), .I1(n6058), .I2(n6059), .O(n6060));
  LUT3 #(.INIT(8'h96)) lut_n6061 (.I0(n5944), .I1(n5982), .I2(n5983), .O(n6061));
  LUT3 #(.INIT(8'hE8)) lut_n6062 (.I0(n6022), .I1(n6060), .I2(n6061), .O(n6062));
  LUT3 #(.INIT(8'h96)) lut_n6063 (.I0(n5824), .I1(n5902), .I2(n5903), .O(n6063));
  LUT3 #(.INIT(8'hE8)) lut_n6064 (.I0(n5984), .I1(n6062), .I2(n6063), .O(n6064));
  LUT3 #(.INIT(8'h96)) lut_n6065 (.I0(x720), .I1(x721), .I2(x722), .O(n6065));
  LUT5 #(.INIT(32'h96696996)) lut_n6066 (.I0(x711), .I1(x712), .I2(x713), .I3(n6052), .I4(n6053), .O(n6066));
  LUT5 #(.INIT(32'hFF969600)) lut_n6067 (.I0(x717), .I1(x718), .I2(x719), .I3(n6065), .I4(n6066), .O(n6067));
  LUT3 #(.INIT(8'h96)) lut_n6068 (.I0(x726), .I1(x727), .I2(x728), .O(n6068));
  LUT5 #(.INIT(32'h96696996)) lut_n6069 (.I0(x717), .I1(x718), .I2(x719), .I3(n6065), .I4(n6066), .O(n6069));
  LUT5 #(.INIT(32'hFF969600)) lut_n6070 (.I0(x723), .I1(x724), .I2(x725), .I3(n6068), .I4(n6069), .O(n6070));
  LUT3 #(.INIT(8'h96)) lut_n6071 (.I0(n6051), .I1(n6054), .I2(n6055), .O(n6071));
  LUT3 #(.INIT(8'hE8)) lut_n6072 (.I0(n6067), .I1(n6070), .I2(n6071), .O(n6072));
  LUT3 #(.INIT(8'h96)) lut_n6073 (.I0(x732), .I1(x733), .I2(x734), .O(n6073));
  LUT5 #(.INIT(32'h96696996)) lut_n6074 (.I0(x723), .I1(x724), .I2(x725), .I3(n6068), .I4(n6069), .O(n6074));
  LUT5 #(.INIT(32'hFF969600)) lut_n6075 (.I0(x729), .I1(x730), .I2(x731), .I3(n6073), .I4(n6074), .O(n6075));
  LUT3 #(.INIT(8'h96)) lut_n6076 (.I0(x738), .I1(x739), .I2(x740), .O(n6076));
  LUT5 #(.INIT(32'h96696996)) lut_n6077 (.I0(x729), .I1(x730), .I2(x731), .I3(n6073), .I4(n6074), .O(n6077));
  LUT5 #(.INIT(32'hFF969600)) lut_n6078 (.I0(x735), .I1(x736), .I2(x737), .I3(n6076), .I4(n6077), .O(n6078));
  LUT3 #(.INIT(8'h96)) lut_n6079 (.I0(n6067), .I1(n6070), .I2(n6071), .O(n6079));
  LUT3 #(.INIT(8'hE8)) lut_n6080 (.I0(n6075), .I1(n6078), .I2(n6079), .O(n6080));
  LUT3 #(.INIT(8'h96)) lut_n6081 (.I0(n6048), .I1(n6056), .I2(n6057), .O(n6081));
  LUT3 #(.INIT(8'hE8)) lut_n6082 (.I0(n6072), .I1(n6080), .I2(n6081), .O(n6082));
  LUT3 #(.INIT(8'h96)) lut_n6083 (.I0(x744), .I1(x745), .I2(x746), .O(n6083));
  LUT5 #(.INIT(32'h96696996)) lut_n6084 (.I0(x735), .I1(x736), .I2(x737), .I3(n6076), .I4(n6077), .O(n6084));
  LUT5 #(.INIT(32'hFF969600)) lut_n6085 (.I0(x741), .I1(x742), .I2(x743), .I3(n6083), .I4(n6084), .O(n6085));
  LUT3 #(.INIT(8'h96)) lut_n6086 (.I0(x750), .I1(x751), .I2(x752), .O(n6086));
  LUT5 #(.INIT(32'h96696996)) lut_n6087 (.I0(x741), .I1(x742), .I2(x743), .I3(n6083), .I4(n6084), .O(n6087));
  LUT5 #(.INIT(32'hFF969600)) lut_n6088 (.I0(x747), .I1(x748), .I2(x749), .I3(n6086), .I4(n6087), .O(n6088));
  LUT3 #(.INIT(8'h96)) lut_n6089 (.I0(n6075), .I1(n6078), .I2(n6079), .O(n6089));
  LUT3 #(.INIT(8'hE8)) lut_n6090 (.I0(n6085), .I1(n6088), .I2(n6089), .O(n6090));
  LUT3 #(.INIT(8'h96)) lut_n6091 (.I0(x756), .I1(x757), .I2(x758), .O(n6091));
  LUT5 #(.INIT(32'h96696996)) lut_n6092 (.I0(x747), .I1(x748), .I2(x749), .I3(n6086), .I4(n6087), .O(n6092));
  LUT5 #(.INIT(32'hFF969600)) lut_n6093 (.I0(x753), .I1(x754), .I2(x755), .I3(n6091), .I4(n6092), .O(n6093));
  LUT3 #(.INIT(8'h96)) lut_n6094 (.I0(x762), .I1(x763), .I2(x764), .O(n6094));
  LUT5 #(.INIT(32'h96696996)) lut_n6095 (.I0(x753), .I1(x754), .I2(x755), .I3(n6091), .I4(n6092), .O(n6095));
  LUT5 #(.INIT(32'hFF969600)) lut_n6096 (.I0(x759), .I1(x760), .I2(x761), .I3(n6094), .I4(n6095), .O(n6096));
  LUT3 #(.INIT(8'h96)) lut_n6097 (.I0(n6085), .I1(n6088), .I2(n6089), .O(n6097));
  LUT3 #(.INIT(8'hE8)) lut_n6098 (.I0(n6093), .I1(n6096), .I2(n6097), .O(n6098));
  LUT3 #(.INIT(8'h96)) lut_n6099 (.I0(n6072), .I1(n6080), .I2(n6081), .O(n6099));
  LUT3 #(.INIT(8'hE8)) lut_n6100 (.I0(n6090), .I1(n6098), .I2(n6099), .O(n6100));
  LUT3 #(.INIT(8'h96)) lut_n6101 (.I0(n6040), .I1(n6058), .I2(n6059), .O(n6101));
  LUT3 #(.INIT(8'hE8)) lut_n6102 (.I0(n6082), .I1(n6100), .I2(n6101), .O(n6102));
  LUT3 #(.INIT(8'h96)) lut_n6103 (.I0(x768), .I1(x769), .I2(x770), .O(n6103));
  LUT5 #(.INIT(32'h96696996)) lut_n6104 (.I0(x759), .I1(x760), .I2(x761), .I3(n6094), .I4(n6095), .O(n6104));
  LUT5 #(.INIT(32'hFF969600)) lut_n6105 (.I0(x765), .I1(x766), .I2(x767), .I3(n6103), .I4(n6104), .O(n6105));
  LUT3 #(.INIT(8'h96)) lut_n6106 (.I0(x774), .I1(x775), .I2(x776), .O(n6106));
  LUT5 #(.INIT(32'h96696996)) lut_n6107 (.I0(x765), .I1(x766), .I2(x767), .I3(n6103), .I4(n6104), .O(n6107));
  LUT5 #(.INIT(32'hFF969600)) lut_n6108 (.I0(x771), .I1(x772), .I2(x773), .I3(n6106), .I4(n6107), .O(n6108));
  LUT3 #(.INIT(8'h96)) lut_n6109 (.I0(n6093), .I1(n6096), .I2(n6097), .O(n6109));
  LUT3 #(.INIT(8'hE8)) lut_n6110 (.I0(n6105), .I1(n6108), .I2(n6109), .O(n6110));
  LUT3 #(.INIT(8'h96)) lut_n6111 (.I0(x780), .I1(x781), .I2(x782), .O(n6111));
  LUT5 #(.INIT(32'h96696996)) lut_n6112 (.I0(x771), .I1(x772), .I2(x773), .I3(n6106), .I4(n6107), .O(n6112));
  LUT5 #(.INIT(32'hFF969600)) lut_n6113 (.I0(x777), .I1(x778), .I2(x779), .I3(n6111), .I4(n6112), .O(n6113));
  LUT3 #(.INIT(8'h96)) lut_n6114 (.I0(x786), .I1(x787), .I2(x788), .O(n6114));
  LUT5 #(.INIT(32'h96696996)) lut_n6115 (.I0(x777), .I1(x778), .I2(x779), .I3(n6111), .I4(n6112), .O(n6115));
  LUT5 #(.INIT(32'hFF969600)) lut_n6116 (.I0(x783), .I1(x784), .I2(x785), .I3(n6114), .I4(n6115), .O(n6116));
  LUT3 #(.INIT(8'h96)) lut_n6117 (.I0(n6105), .I1(n6108), .I2(n6109), .O(n6117));
  LUT3 #(.INIT(8'hE8)) lut_n6118 (.I0(n6113), .I1(n6116), .I2(n6117), .O(n6118));
  LUT3 #(.INIT(8'h96)) lut_n6119 (.I0(n6090), .I1(n6098), .I2(n6099), .O(n6119));
  LUT3 #(.INIT(8'hE8)) lut_n6120 (.I0(n6110), .I1(n6118), .I2(n6119), .O(n6120));
  LUT3 #(.INIT(8'h96)) lut_n6121 (.I0(x792), .I1(x793), .I2(x794), .O(n6121));
  LUT5 #(.INIT(32'h96696996)) lut_n6122 (.I0(x783), .I1(x784), .I2(x785), .I3(n6114), .I4(n6115), .O(n6122));
  LUT5 #(.INIT(32'hFF969600)) lut_n6123 (.I0(x789), .I1(x790), .I2(x791), .I3(n6121), .I4(n6122), .O(n6123));
  LUT3 #(.INIT(8'h96)) lut_n6124 (.I0(x798), .I1(x799), .I2(x800), .O(n6124));
  LUT5 #(.INIT(32'h96696996)) lut_n6125 (.I0(x789), .I1(x790), .I2(x791), .I3(n6121), .I4(n6122), .O(n6125));
  LUT5 #(.INIT(32'hFF969600)) lut_n6126 (.I0(x795), .I1(x796), .I2(x797), .I3(n6124), .I4(n6125), .O(n6126));
  LUT3 #(.INIT(8'h96)) lut_n6127 (.I0(n6113), .I1(n6116), .I2(n6117), .O(n6127));
  LUT3 #(.INIT(8'hE8)) lut_n6128 (.I0(n6123), .I1(n6126), .I2(n6127), .O(n6128));
  LUT3 #(.INIT(8'h96)) lut_n6129 (.I0(x804), .I1(x805), .I2(x806), .O(n6129));
  LUT5 #(.INIT(32'h96696996)) lut_n6130 (.I0(x795), .I1(x796), .I2(x797), .I3(n6124), .I4(n6125), .O(n6130));
  LUT5 #(.INIT(32'hFF969600)) lut_n6131 (.I0(x801), .I1(x802), .I2(x803), .I3(n6129), .I4(n6130), .O(n6131));
  LUT3 #(.INIT(8'h96)) lut_n6132 (.I0(x810), .I1(x811), .I2(x812), .O(n6132));
  LUT5 #(.INIT(32'h96696996)) lut_n6133 (.I0(x801), .I1(x802), .I2(x803), .I3(n6129), .I4(n6130), .O(n6133));
  LUT5 #(.INIT(32'hFF969600)) lut_n6134 (.I0(x807), .I1(x808), .I2(x809), .I3(n6132), .I4(n6133), .O(n6134));
  LUT3 #(.INIT(8'h96)) lut_n6135 (.I0(n6123), .I1(n6126), .I2(n6127), .O(n6135));
  LUT3 #(.INIT(8'hE8)) lut_n6136 (.I0(n6131), .I1(n6134), .I2(n6135), .O(n6136));
  LUT3 #(.INIT(8'h96)) lut_n6137 (.I0(n6110), .I1(n6118), .I2(n6119), .O(n6137));
  LUT3 #(.INIT(8'hE8)) lut_n6138 (.I0(n6128), .I1(n6136), .I2(n6137), .O(n6138));
  LUT3 #(.INIT(8'h96)) lut_n6139 (.I0(n6082), .I1(n6100), .I2(n6101), .O(n6139));
  LUT3 #(.INIT(8'hE8)) lut_n6140 (.I0(n6120), .I1(n6138), .I2(n6139), .O(n6140));
  LUT3 #(.INIT(8'h96)) lut_n6141 (.I0(n6022), .I1(n6060), .I2(n6061), .O(n6141));
  LUT3 #(.INIT(8'hE8)) lut_n6142 (.I0(n6102), .I1(n6140), .I2(n6141), .O(n6142));
  LUT3 #(.INIT(8'h96)) lut_n6143 (.I0(x816), .I1(x817), .I2(x818), .O(n6143));
  LUT5 #(.INIT(32'h96696996)) lut_n6144 (.I0(x807), .I1(x808), .I2(x809), .I3(n6132), .I4(n6133), .O(n6144));
  LUT5 #(.INIT(32'hFF969600)) lut_n6145 (.I0(x813), .I1(x814), .I2(x815), .I3(n6143), .I4(n6144), .O(n6145));
  LUT3 #(.INIT(8'h96)) lut_n6146 (.I0(x822), .I1(x823), .I2(x824), .O(n6146));
  LUT5 #(.INIT(32'h96696996)) lut_n6147 (.I0(x813), .I1(x814), .I2(x815), .I3(n6143), .I4(n6144), .O(n6147));
  LUT5 #(.INIT(32'hFF969600)) lut_n6148 (.I0(x819), .I1(x820), .I2(x821), .I3(n6146), .I4(n6147), .O(n6148));
  LUT3 #(.INIT(8'h96)) lut_n6149 (.I0(n6131), .I1(n6134), .I2(n6135), .O(n6149));
  LUT3 #(.INIT(8'hE8)) lut_n6150 (.I0(n6145), .I1(n6148), .I2(n6149), .O(n6150));
  LUT3 #(.INIT(8'h96)) lut_n6151 (.I0(x828), .I1(x829), .I2(x830), .O(n6151));
  LUT5 #(.INIT(32'h96696996)) lut_n6152 (.I0(x819), .I1(x820), .I2(x821), .I3(n6146), .I4(n6147), .O(n6152));
  LUT5 #(.INIT(32'hFF969600)) lut_n6153 (.I0(x825), .I1(x826), .I2(x827), .I3(n6151), .I4(n6152), .O(n6153));
  LUT3 #(.INIT(8'h96)) lut_n6154 (.I0(x834), .I1(x835), .I2(x836), .O(n6154));
  LUT5 #(.INIT(32'h96696996)) lut_n6155 (.I0(x825), .I1(x826), .I2(x827), .I3(n6151), .I4(n6152), .O(n6155));
  LUT5 #(.INIT(32'hFF969600)) lut_n6156 (.I0(x831), .I1(x832), .I2(x833), .I3(n6154), .I4(n6155), .O(n6156));
  LUT3 #(.INIT(8'h96)) lut_n6157 (.I0(n6145), .I1(n6148), .I2(n6149), .O(n6157));
  LUT3 #(.INIT(8'hE8)) lut_n6158 (.I0(n6153), .I1(n6156), .I2(n6157), .O(n6158));
  LUT3 #(.INIT(8'h96)) lut_n6159 (.I0(n6128), .I1(n6136), .I2(n6137), .O(n6159));
  LUT3 #(.INIT(8'hE8)) lut_n6160 (.I0(n6150), .I1(n6158), .I2(n6159), .O(n6160));
  LUT3 #(.INIT(8'h96)) lut_n6161 (.I0(x840), .I1(x841), .I2(x842), .O(n6161));
  LUT5 #(.INIT(32'h96696996)) lut_n6162 (.I0(x831), .I1(x832), .I2(x833), .I3(n6154), .I4(n6155), .O(n6162));
  LUT5 #(.INIT(32'hFF969600)) lut_n6163 (.I0(x837), .I1(x838), .I2(x839), .I3(n6161), .I4(n6162), .O(n6163));
  LUT3 #(.INIT(8'h96)) lut_n6164 (.I0(x846), .I1(x847), .I2(x848), .O(n6164));
  LUT5 #(.INIT(32'h96696996)) lut_n6165 (.I0(x837), .I1(x838), .I2(x839), .I3(n6161), .I4(n6162), .O(n6165));
  LUT5 #(.INIT(32'hFF969600)) lut_n6166 (.I0(x843), .I1(x844), .I2(x845), .I3(n6164), .I4(n6165), .O(n6166));
  LUT3 #(.INIT(8'h96)) lut_n6167 (.I0(n6153), .I1(n6156), .I2(n6157), .O(n6167));
  LUT3 #(.INIT(8'hE8)) lut_n6168 (.I0(n6163), .I1(n6166), .I2(n6167), .O(n6168));
  LUT3 #(.INIT(8'h96)) lut_n6169 (.I0(x852), .I1(x853), .I2(x854), .O(n6169));
  LUT5 #(.INIT(32'h96696996)) lut_n6170 (.I0(x843), .I1(x844), .I2(x845), .I3(n6164), .I4(n6165), .O(n6170));
  LUT5 #(.INIT(32'hFF969600)) lut_n6171 (.I0(x849), .I1(x850), .I2(x851), .I3(n6169), .I4(n6170), .O(n6171));
  LUT3 #(.INIT(8'h96)) lut_n6172 (.I0(x858), .I1(x859), .I2(x860), .O(n6172));
  LUT5 #(.INIT(32'h96696996)) lut_n6173 (.I0(x849), .I1(x850), .I2(x851), .I3(n6169), .I4(n6170), .O(n6173));
  LUT5 #(.INIT(32'hFF969600)) lut_n6174 (.I0(x855), .I1(x856), .I2(x857), .I3(n6172), .I4(n6173), .O(n6174));
  LUT3 #(.INIT(8'h96)) lut_n6175 (.I0(n6163), .I1(n6166), .I2(n6167), .O(n6175));
  LUT3 #(.INIT(8'hE8)) lut_n6176 (.I0(n6171), .I1(n6174), .I2(n6175), .O(n6176));
  LUT3 #(.INIT(8'h96)) lut_n6177 (.I0(n6150), .I1(n6158), .I2(n6159), .O(n6177));
  LUT3 #(.INIT(8'hE8)) lut_n6178 (.I0(n6168), .I1(n6176), .I2(n6177), .O(n6178));
  LUT3 #(.INIT(8'h96)) lut_n6179 (.I0(n6120), .I1(n6138), .I2(n6139), .O(n6179));
  LUT3 #(.INIT(8'hE8)) lut_n6180 (.I0(n6160), .I1(n6178), .I2(n6179), .O(n6180));
  LUT3 #(.INIT(8'h96)) lut_n6181 (.I0(x864), .I1(x865), .I2(x866), .O(n6181));
  LUT5 #(.INIT(32'h96696996)) lut_n6182 (.I0(x855), .I1(x856), .I2(x857), .I3(n6172), .I4(n6173), .O(n6182));
  LUT5 #(.INIT(32'hFF969600)) lut_n6183 (.I0(x861), .I1(x862), .I2(x863), .I3(n6181), .I4(n6182), .O(n6183));
  LUT3 #(.INIT(8'h96)) lut_n6184 (.I0(x870), .I1(x871), .I2(x872), .O(n6184));
  LUT5 #(.INIT(32'h96696996)) lut_n6185 (.I0(x861), .I1(x862), .I2(x863), .I3(n6181), .I4(n6182), .O(n6185));
  LUT5 #(.INIT(32'hFF969600)) lut_n6186 (.I0(x867), .I1(x868), .I2(x869), .I3(n6184), .I4(n6185), .O(n6186));
  LUT3 #(.INIT(8'h96)) lut_n6187 (.I0(n6171), .I1(n6174), .I2(n6175), .O(n6187));
  LUT3 #(.INIT(8'hE8)) lut_n6188 (.I0(n6183), .I1(n6186), .I2(n6187), .O(n6188));
  LUT3 #(.INIT(8'h96)) lut_n6189 (.I0(x876), .I1(x877), .I2(x878), .O(n6189));
  LUT5 #(.INIT(32'h96696996)) lut_n6190 (.I0(x867), .I1(x868), .I2(x869), .I3(n6184), .I4(n6185), .O(n6190));
  LUT5 #(.INIT(32'hFF969600)) lut_n6191 (.I0(x873), .I1(x874), .I2(x875), .I3(n6189), .I4(n6190), .O(n6191));
  LUT3 #(.INIT(8'h96)) lut_n6192 (.I0(x882), .I1(x883), .I2(x884), .O(n6192));
  LUT5 #(.INIT(32'h96696996)) lut_n6193 (.I0(x873), .I1(x874), .I2(x875), .I3(n6189), .I4(n6190), .O(n6193));
  LUT5 #(.INIT(32'hFF969600)) lut_n6194 (.I0(x879), .I1(x880), .I2(x881), .I3(n6192), .I4(n6193), .O(n6194));
  LUT3 #(.INIT(8'h96)) lut_n6195 (.I0(n6183), .I1(n6186), .I2(n6187), .O(n6195));
  LUT3 #(.INIT(8'hE8)) lut_n6196 (.I0(n6191), .I1(n6194), .I2(n6195), .O(n6196));
  LUT3 #(.INIT(8'h96)) lut_n6197 (.I0(n6168), .I1(n6176), .I2(n6177), .O(n6197));
  LUT3 #(.INIT(8'hE8)) lut_n6198 (.I0(n6188), .I1(n6196), .I2(n6197), .O(n6198));
  LUT3 #(.INIT(8'h96)) lut_n6199 (.I0(x888), .I1(x889), .I2(x890), .O(n6199));
  LUT5 #(.INIT(32'h96696996)) lut_n6200 (.I0(x879), .I1(x880), .I2(x881), .I3(n6192), .I4(n6193), .O(n6200));
  LUT5 #(.INIT(32'hFF969600)) lut_n6201 (.I0(x885), .I1(x886), .I2(x887), .I3(n6199), .I4(n6200), .O(n6201));
  LUT3 #(.INIT(8'h96)) lut_n6202 (.I0(x894), .I1(x895), .I2(x896), .O(n6202));
  LUT5 #(.INIT(32'h96696996)) lut_n6203 (.I0(x885), .I1(x886), .I2(x887), .I3(n6199), .I4(n6200), .O(n6203));
  LUT5 #(.INIT(32'hFF969600)) lut_n6204 (.I0(x891), .I1(x892), .I2(x893), .I3(n6202), .I4(n6203), .O(n6204));
  LUT3 #(.INIT(8'h96)) lut_n6205 (.I0(n6191), .I1(n6194), .I2(n6195), .O(n6205));
  LUT3 #(.INIT(8'hE8)) lut_n6206 (.I0(n6201), .I1(n6204), .I2(n6205), .O(n6206));
  LUT3 #(.INIT(8'h96)) lut_n6207 (.I0(x900), .I1(x901), .I2(x902), .O(n6207));
  LUT5 #(.INIT(32'h96696996)) lut_n6208 (.I0(x891), .I1(x892), .I2(x893), .I3(n6202), .I4(n6203), .O(n6208));
  LUT5 #(.INIT(32'hFF969600)) lut_n6209 (.I0(x897), .I1(x898), .I2(x899), .I3(n6207), .I4(n6208), .O(n6209));
  LUT3 #(.INIT(8'h96)) lut_n6210 (.I0(x906), .I1(x907), .I2(x908), .O(n6210));
  LUT5 #(.INIT(32'h96696996)) lut_n6211 (.I0(x897), .I1(x898), .I2(x899), .I3(n6207), .I4(n6208), .O(n6211));
  LUT5 #(.INIT(32'hFF969600)) lut_n6212 (.I0(x903), .I1(x904), .I2(x905), .I3(n6210), .I4(n6211), .O(n6212));
  LUT3 #(.INIT(8'h96)) lut_n6213 (.I0(n6201), .I1(n6204), .I2(n6205), .O(n6213));
  LUT3 #(.INIT(8'hE8)) lut_n6214 (.I0(n6209), .I1(n6212), .I2(n6213), .O(n6214));
  LUT3 #(.INIT(8'h96)) lut_n6215 (.I0(n6188), .I1(n6196), .I2(n6197), .O(n6215));
  LUT3 #(.INIT(8'hE8)) lut_n6216 (.I0(n6206), .I1(n6214), .I2(n6215), .O(n6216));
  LUT3 #(.INIT(8'h96)) lut_n6217 (.I0(n6160), .I1(n6178), .I2(n6179), .O(n6217));
  LUT3 #(.INIT(8'hE8)) lut_n6218 (.I0(n6198), .I1(n6216), .I2(n6217), .O(n6218));
  LUT3 #(.INIT(8'h96)) lut_n6219 (.I0(n6102), .I1(n6140), .I2(n6141), .O(n6219));
  LUT3 #(.INIT(8'hE8)) lut_n6220 (.I0(n6180), .I1(n6218), .I2(n6219), .O(n6220));
  LUT3 #(.INIT(8'h96)) lut_n6221 (.I0(n5984), .I1(n6062), .I2(n6063), .O(n6221));
  LUT3 #(.INIT(8'hE8)) lut_n6222 (.I0(n6142), .I1(n6220), .I2(n6221), .O(n6222));
  LUT3 #(.INIT(8'h96)) lut_n6223 (.I0(n5746), .I1(n5904), .I2(n5905), .O(n6223));
  LUT3 #(.INIT(8'hE8)) lut_n6224 (.I0(n6064), .I1(n6222), .I2(n6223), .O(n6224));
  LUT3 #(.INIT(8'h96)) lut_n6225 (.I0(n5368), .I1(n5583), .I2(n5584), .O(n6225));
  LUT3 #(.INIT(8'hE8)) lut_n6226 (.I0(n5906), .I1(n6224), .I2(n6225), .O(n6226));
  LUT3 #(.INIT(8'h96)) lut_n6227 (.I0(x912), .I1(x913), .I2(x914), .O(n6227));
  LUT5 #(.INIT(32'h96696996)) lut_n6228 (.I0(x903), .I1(x904), .I2(x905), .I3(n6210), .I4(n6211), .O(n6228));
  LUT5 #(.INIT(32'hFF969600)) lut_n6229 (.I0(x909), .I1(x910), .I2(x911), .I3(n6227), .I4(n6228), .O(n6229));
  LUT3 #(.INIT(8'h96)) lut_n6230 (.I0(x918), .I1(x919), .I2(x920), .O(n6230));
  LUT5 #(.INIT(32'h96696996)) lut_n6231 (.I0(x909), .I1(x910), .I2(x911), .I3(n6227), .I4(n6228), .O(n6231));
  LUT5 #(.INIT(32'hFF969600)) lut_n6232 (.I0(x915), .I1(x916), .I2(x917), .I3(n6230), .I4(n6231), .O(n6232));
  LUT3 #(.INIT(8'h96)) lut_n6233 (.I0(n6209), .I1(n6212), .I2(n6213), .O(n6233));
  LUT3 #(.INIT(8'hE8)) lut_n6234 (.I0(n6229), .I1(n6232), .I2(n6233), .O(n6234));
  LUT3 #(.INIT(8'h96)) lut_n6235 (.I0(x924), .I1(x925), .I2(x926), .O(n6235));
  LUT5 #(.INIT(32'h96696996)) lut_n6236 (.I0(x915), .I1(x916), .I2(x917), .I3(n6230), .I4(n6231), .O(n6236));
  LUT5 #(.INIT(32'hFF969600)) lut_n6237 (.I0(x921), .I1(x922), .I2(x923), .I3(n6235), .I4(n6236), .O(n6237));
  LUT3 #(.INIT(8'h96)) lut_n6238 (.I0(x930), .I1(x931), .I2(x932), .O(n6238));
  LUT5 #(.INIT(32'h96696996)) lut_n6239 (.I0(x921), .I1(x922), .I2(x923), .I3(n6235), .I4(n6236), .O(n6239));
  LUT5 #(.INIT(32'hFF969600)) lut_n6240 (.I0(x927), .I1(x928), .I2(x929), .I3(n6238), .I4(n6239), .O(n6240));
  LUT3 #(.INIT(8'h96)) lut_n6241 (.I0(n6229), .I1(n6232), .I2(n6233), .O(n6241));
  LUT3 #(.INIT(8'hE8)) lut_n6242 (.I0(n6237), .I1(n6240), .I2(n6241), .O(n6242));
  LUT3 #(.INIT(8'h96)) lut_n6243 (.I0(n6206), .I1(n6214), .I2(n6215), .O(n6243));
  LUT3 #(.INIT(8'hE8)) lut_n6244 (.I0(n6234), .I1(n6242), .I2(n6243), .O(n6244));
  LUT3 #(.INIT(8'h96)) lut_n6245 (.I0(x936), .I1(x937), .I2(x938), .O(n6245));
  LUT5 #(.INIT(32'h96696996)) lut_n6246 (.I0(x927), .I1(x928), .I2(x929), .I3(n6238), .I4(n6239), .O(n6246));
  LUT5 #(.INIT(32'hFF969600)) lut_n6247 (.I0(x933), .I1(x934), .I2(x935), .I3(n6245), .I4(n6246), .O(n6247));
  LUT3 #(.INIT(8'h96)) lut_n6248 (.I0(x942), .I1(x943), .I2(x944), .O(n6248));
  LUT5 #(.INIT(32'h96696996)) lut_n6249 (.I0(x933), .I1(x934), .I2(x935), .I3(n6245), .I4(n6246), .O(n6249));
  LUT5 #(.INIT(32'hFF969600)) lut_n6250 (.I0(x939), .I1(x940), .I2(x941), .I3(n6248), .I4(n6249), .O(n6250));
  LUT3 #(.INIT(8'h96)) lut_n6251 (.I0(n6237), .I1(n6240), .I2(n6241), .O(n6251));
  LUT3 #(.INIT(8'hE8)) lut_n6252 (.I0(n6247), .I1(n6250), .I2(n6251), .O(n6252));
  LUT3 #(.INIT(8'h96)) lut_n6253 (.I0(x948), .I1(x949), .I2(x950), .O(n6253));
  LUT5 #(.INIT(32'h96696996)) lut_n6254 (.I0(x939), .I1(x940), .I2(x941), .I3(n6248), .I4(n6249), .O(n6254));
  LUT5 #(.INIT(32'hFF969600)) lut_n6255 (.I0(x945), .I1(x946), .I2(x947), .I3(n6253), .I4(n6254), .O(n6255));
  LUT3 #(.INIT(8'h96)) lut_n6256 (.I0(x954), .I1(x955), .I2(x956), .O(n6256));
  LUT5 #(.INIT(32'h96696996)) lut_n6257 (.I0(x945), .I1(x946), .I2(x947), .I3(n6253), .I4(n6254), .O(n6257));
  LUT5 #(.INIT(32'hFF969600)) lut_n6258 (.I0(x951), .I1(x952), .I2(x953), .I3(n6256), .I4(n6257), .O(n6258));
  LUT3 #(.INIT(8'h96)) lut_n6259 (.I0(n6247), .I1(n6250), .I2(n6251), .O(n6259));
  LUT3 #(.INIT(8'hE8)) lut_n6260 (.I0(n6255), .I1(n6258), .I2(n6259), .O(n6260));
  LUT3 #(.INIT(8'h96)) lut_n6261 (.I0(n6234), .I1(n6242), .I2(n6243), .O(n6261));
  LUT3 #(.INIT(8'hE8)) lut_n6262 (.I0(n6252), .I1(n6260), .I2(n6261), .O(n6262));
  LUT3 #(.INIT(8'h96)) lut_n6263 (.I0(n6198), .I1(n6216), .I2(n6217), .O(n6263));
  LUT3 #(.INIT(8'hE8)) lut_n6264 (.I0(n6244), .I1(n6262), .I2(n6263), .O(n6264));
  LUT3 #(.INIT(8'h96)) lut_n6265 (.I0(x960), .I1(x961), .I2(x962), .O(n6265));
  LUT5 #(.INIT(32'h96696996)) lut_n6266 (.I0(x951), .I1(x952), .I2(x953), .I3(n6256), .I4(n6257), .O(n6266));
  LUT5 #(.INIT(32'hFF969600)) lut_n6267 (.I0(x957), .I1(x958), .I2(x959), .I3(n6265), .I4(n6266), .O(n6267));
  LUT3 #(.INIT(8'h96)) lut_n6268 (.I0(x966), .I1(x967), .I2(x968), .O(n6268));
  LUT5 #(.INIT(32'h96696996)) lut_n6269 (.I0(x957), .I1(x958), .I2(x959), .I3(n6265), .I4(n6266), .O(n6269));
  LUT5 #(.INIT(32'hFF969600)) lut_n6270 (.I0(x963), .I1(x964), .I2(x965), .I3(n6268), .I4(n6269), .O(n6270));
  LUT3 #(.INIT(8'h96)) lut_n6271 (.I0(n6255), .I1(n6258), .I2(n6259), .O(n6271));
  LUT3 #(.INIT(8'hE8)) lut_n6272 (.I0(n6267), .I1(n6270), .I2(n6271), .O(n6272));
  LUT3 #(.INIT(8'h96)) lut_n6273 (.I0(x972), .I1(x973), .I2(x974), .O(n6273));
  LUT5 #(.INIT(32'h96696996)) lut_n6274 (.I0(x963), .I1(x964), .I2(x965), .I3(n6268), .I4(n6269), .O(n6274));
  LUT5 #(.INIT(32'hFF969600)) lut_n6275 (.I0(x969), .I1(x970), .I2(x971), .I3(n6273), .I4(n6274), .O(n6275));
  LUT3 #(.INIT(8'h96)) lut_n6276 (.I0(x978), .I1(x979), .I2(x980), .O(n6276));
  LUT5 #(.INIT(32'h96696996)) lut_n6277 (.I0(x969), .I1(x970), .I2(x971), .I3(n6273), .I4(n6274), .O(n6277));
  LUT5 #(.INIT(32'hFF969600)) lut_n6278 (.I0(x975), .I1(x976), .I2(x977), .I3(n6276), .I4(n6277), .O(n6278));
  LUT3 #(.INIT(8'h96)) lut_n6279 (.I0(n6267), .I1(n6270), .I2(n6271), .O(n6279));
  LUT3 #(.INIT(8'hE8)) lut_n6280 (.I0(n6275), .I1(n6278), .I2(n6279), .O(n6280));
  LUT3 #(.INIT(8'h96)) lut_n6281 (.I0(n6252), .I1(n6260), .I2(n6261), .O(n6281));
  LUT3 #(.INIT(8'hE8)) lut_n6282 (.I0(n6272), .I1(n6280), .I2(n6281), .O(n6282));
  LUT3 #(.INIT(8'h96)) lut_n6283 (.I0(x984), .I1(x985), .I2(x986), .O(n6283));
  LUT5 #(.INIT(32'h96696996)) lut_n6284 (.I0(x975), .I1(x976), .I2(x977), .I3(n6276), .I4(n6277), .O(n6284));
  LUT5 #(.INIT(32'hFF969600)) lut_n6285 (.I0(x981), .I1(x982), .I2(x983), .I3(n6283), .I4(n6284), .O(n6285));
  LUT3 #(.INIT(8'h96)) lut_n6286 (.I0(x990), .I1(x991), .I2(x992), .O(n6286));
  LUT5 #(.INIT(32'h96696996)) lut_n6287 (.I0(x981), .I1(x982), .I2(x983), .I3(n6283), .I4(n6284), .O(n6287));
  LUT5 #(.INIT(32'hFF969600)) lut_n6288 (.I0(x987), .I1(x988), .I2(x989), .I3(n6286), .I4(n6287), .O(n6288));
  LUT3 #(.INIT(8'h96)) lut_n6289 (.I0(n6275), .I1(n6278), .I2(n6279), .O(n6289));
  LUT3 #(.INIT(8'hE8)) lut_n6290 (.I0(n6285), .I1(n6288), .I2(n6289), .O(n6290));
  LUT3 #(.INIT(8'h96)) lut_n6291 (.I0(x996), .I1(x997), .I2(x998), .O(n6291));
  LUT5 #(.INIT(32'h96696996)) lut_n6292 (.I0(x987), .I1(x988), .I2(x989), .I3(n6286), .I4(n6287), .O(n6292));
  LUT5 #(.INIT(32'hFF969600)) lut_n6293 (.I0(x993), .I1(x994), .I2(x995), .I3(n6291), .I4(n6292), .O(n6293));
  LUT3 #(.INIT(8'h96)) lut_n6294 (.I0(x1002), .I1(x1003), .I2(x1004), .O(n6294));
  LUT5 #(.INIT(32'h96696996)) lut_n6295 (.I0(x993), .I1(x994), .I2(x995), .I3(n6291), .I4(n6292), .O(n6295));
  LUT5 #(.INIT(32'hFF969600)) lut_n6296 (.I0(x999), .I1(x1000), .I2(x1001), .I3(n6294), .I4(n6295), .O(n6296));
  LUT3 #(.INIT(8'h96)) lut_n6297 (.I0(n6285), .I1(n6288), .I2(n6289), .O(n6297));
  LUT3 #(.INIT(8'hE8)) lut_n6298 (.I0(n6293), .I1(n6296), .I2(n6297), .O(n6298));
  LUT3 #(.INIT(8'h96)) lut_n6299 (.I0(n6272), .I1(n6280), .I2(n6281), .O(n6299));
  LUT3 #(.INIT(8'hE8)) lut_n6300 (.I0(n6290), .I1(n6298), .I2(n6299), .O(n6300));
  LUT3 #(.INIT(8'h96)) lut_n6301 (.I0(n6244), .I1(n6262), .I2(n6263), .O(n6301));
  LUT3 #(.INIT(8'hE8)) lut_n6302 (.I0(n6282), .I1(n6300), .I2(n6301), .O(n6302));
  LUT3 #(.INIT(8'h96)) lut_n6303 (.I0(n6180), .I1(n6218), .I2(n6219), .O(n6303));
  LUT3 #(.INIT(8'hE8)) lut_n6304 (.I0(n6264), .I1(n6302), .I2(n6303), .O(n6304));
  LUT3 #(.INIT(8'h96)) lut_n6305 (.I0(x1008), .I1(x1009), .I2(x1010), .O(n6305));
  LUT5 #(.INIT(32'h96696996)) lut_n6306 (.I0(x999), .I1(x1000), .I2(x1001), .I3(n6294), .I4(n6295), .O(n6306));
  LUT5 #(.INIT(32'hFF969600)) lut_n6307 (.I0(x1005), .I1(x1006), .I2(x1007), .I3(n6305), .I4(n6306), .O(n6307));
  LUT3 #(.INIT(8'h96)) lut_n6308 (.I0(x1014), .I1(x1015), .I2(x1016), .O(n6308));
  LUT5 #(.INIT(32'h96696996)) lut_n6309 (.I0(x1005), .I1(x1006), .I2(x1007), .I3(n6305), .I4(n6306), .O(n6309));
  LUT5 #(.INIT(32'hFF969600)) lut_n6310 (.I0(x1011), .I1(x1012), .I2(x1013), .I3(n6308), .I4(n6309), .O(n6310));
  LUT3 #(.INIT(8'h96)) lut_n6311 (.I0(n6293), .I1(n6296), .I2(n6297), .O(n6311));
  LUT3 #(.INIT(8'hE8)) lut_n6312 (.I0(n6307), .I1(n6310), .I2(n6311), .O(n6312));
  LUT3 #(.INIT(8'h96)) lut_n6313 (.I0(x1020), .I1(x1021), .I2(x1022), .O(n6313));
  LUT5 #(.INIT(32'h96696996)) lut_n6314 (.I0(x1011), .I1(x1012), .I2(x1013), .I3(n6308), .I4(n6309), .O(n6314));
  LUT5 #(.INIT(32'hFF969600)) lut_n6315 (.I0(x1017), .I1(x1018), .I2(x1019), .I3(n6313), .I4(n6314), .O(n6315));
  LUT3 #(.INIT(8'h96)) lut_n6316 (.I0(x1026), .I1(x1027), .I2(x1028), .O(n6316));
  LUT5 #(.INIT(32'h96696996)) lut_n6317 (.I0(x1017), .I1(x1018), .I2(x1019), .I3(n6313), .I4(n6314), .O(n6317));
  LUT5 #(.INIT(32'hFF969600)) lut_n6318 (.I0(x1023), .I1(x1024), .I2(x1025), .I3(n6316), .I4(n6317), .O(n6318));
  LUT3 #(.INIT(8'h96)) lut_n6319 (.I0(n6307), .I1(n6310), .I2(n6311), .O(n6319));
  LUT3 #(.INIT(8'hE8)) lut_n6320 (.I0(n6315), .I1(n6318), .I2(n6319), .O(n6320));
  LUT3 #(.INIT(8'h96)) lut_n6321 (.I0(n6290), .I1(n6298), .I2(n6299), .O(n6321));
  LUT3 #(.INIT(8'hE8)) lut_n6322 (.I0(n6312), .I1(n6320), .I2(n6321), .O(n6322));
  LUT3 #(.INIT(8'h96)) lut_n6323 (.I0(x1032), .I1(x1033), .I2(x1034), .O(n6323));
  LUT5 #(.INIT(32'h96696996)) lut_n6324 (.I0(x1023), .I1(x1024), .I2(x1025), .I3(n6316), .I4(n6317), .O(n6324));
  LUT5 #(.INIT(32'hFF969600)) lut_n6325 (.I0(x1029), .I1(x1030), .I2(x1031), .I3(n6323), .I4(n6324), .O(n6325));
  LUT3 #(.INIT(8'h96)) lut_n6326 (.I0(x1038), .I1(x1039), .I2(x1040), .O(n6326));
  LUT5 #(.INIT(32'h96696996)) lut_n6327 (.I0(x1029), .I1(x1030), .I2(x1031), .I3(n6323), .I4(n6324), .O(n6327));
  LUT5 #(.INIT(32'hFF969600)) lut_n6328 (.I0(x1035), .I1(x1036), .I2(x1037), .I3(n6326), .I4(n6327), .O(n6328));
  LUT3 #(.INIT(8'h96)) lut_n6329 (.I0(n6315), .I1(n6318), .I2(n6319), .O(n6329));
  LUT3 #(.INIT(8'hE8)) lut_n6330 (.I0(n6325), .I1(n6328), .I2(n6329), .O(n6330));
  LUT3 #(.INIT(8'h96)) lut_n6331 (.I0(x1044), .I1(x1045), .I2(x1046), .O(n6331));
  LUT5 #(.INIT(32'h96696996)) lut_n6332 (.I0(x1035), .I1(x1036), .I2(x1037), .I3(n6326), .I4(n6327), .O(n6332));
  LUT5 #(.INIT(32'hFF969600)) lut_n6333 (.I0(x1041), .I1(x1042), .I2(x1043), .I3(n6331), .I4(n6332), .O(n6333));
  LUT3 #(.INIT(8'h96)) lut_n6334 (.I0(x1050), .I1(x1051), .I2(x1052), .O(n6334));
  LUT5 #(.INIT(32'h96696996)) lut_n6335 (.I0(x1041), .I1(x1042), .I2(x1043), .I3(n6331), .I4(n6332), .O(n6335));
  LUT5 #(.INIT(32'hFF969600)) lut_n6336 (.I0(x1047), .I1(x1048), .I2(x1049), .I3(n6334), .I4(n6335), .O(n6336));
  LUT3 #(.INIT(8'h96)) lut_n6337 (.I0(n6325), .I1(n6328), .I2(n6329), .O(n6337));
  LUT3 #(.INIT(8'hE8)) lut_n6338 (.I0(n6333), .I1(n6336), .I2(n6337), .O(n6338));
  LUT3 #(.INIT(8'h96)) lut_n6339 (.I0(n6312), .I1(n6320), .I2(n6321), .O(n6339));
  LUT3 #(.INIT(8'hE8)) lut_n6340 (.I0(n6330), .I1(n6338), .I2(n6339), .O(n6340));
  LUT3 #(.INIT(8'h96)) lut_n6341 (.I0(n6282), .I1(n6300), .I2(n6301), .O(n6341));
  LUT3 #(.INIT(8'hE8)) lut_n6342 (.I0(n6322), .I1(n6340), .I2(n6341), .O(n6342));
  LUT3 #(.INIT(8'h96)) lut_n6343 (.I0(x1056), .I1(x1057), .I2(x1058), .O(n6343));
  LUT5 #(.INIT(32'h96696996)) lut_n6344 (.I0(x1047), .I1(x1048), .I2(x1049), .I3(n6334), .I4(n6335), .O(n6344));
  LUT5 #(.INIT(32'hFF969600)) lut_n6345 (.I0(x1053), .I1(x1054), .I2(x1055), .I3(n6343), .I4(n6344), .O(n6345));
  LUT3 #(.INIT(8'h96)) lut_n6346 (.I0(x1062), .I1(x1063), .I2(x1064), .O(n6346));
  LUT5 #(.INIT(32'h96696996)) lut_n6347 (.I0(x1053), .I1(x1054), .I2(x1055), .I3(n6343), .I4(n6344), .O(n6347));
  LUT5 #(.INIT(32'hFF969600)) lut_n6348 (.I0(x1059), .I1(x1060), .I2(x1061), .I3(n6346), .I4(n6347), .O(n6348));
  LUT3 #(.INIT(8'h96)) lut_n6349 (.I0(n6333), .I1(n6336), .I2(n6337), .O(n6349));
  LUT3 #(.INIT(8'hE8)) lut_n6350 (.I0(n6345), .I1(n6348), .I2(n6349), .O(n6350));
  LUT3 #(.INIT(8'h96)) lut_n6351 (.I0(x1068), .I1(x1069), .I2(x1070), .O(n6351));
  LUT5 #(.INIT(32'h96696996)) lut_n6352 (.I0(x1059), .I1(x1060), .I2(x1061), .I3(n6346), .I4(n6347), .O(n6352));
  LUT5 #(.INIT(32'hFF969600)) lut_n6353 (.I0(x1065), .I1(x1066), .I2(x1067), .I3(n6351), .I4(n6352), .O(n6353));
  LUT3 #(.INIT(8'h96)) lut_n6354 (.I0(x1074), .I1(x1075), .I2(x1076), .O(n6354));
  LUT5 #(.INIT(32'h96696996)) lut_n6355 (.I0(x1065), .I1(x1066), .I2(x1067), .I3(n6351), .I4(n6352), .O(n6355));
  LUT5 #(.INIT(32'hFF969600)) lut_n6356 (.I0(x1071), .I1(x1072), .I2(x1073), .I3(n6354), .I4(n6355), .O(n6356));
  LUT3 #(.INIT(8'h96)) lut_n6357 (.I0(n6345), .I1(n6348), .I2(n6349), .O(n6357));
  LUT3 #(.INIT(8'hE8)) lut_n6358 (.I0(n6353), .I1(n6356), .I2(n6357), .O(n6358));
  LUT3 #(.INIT(8'h96)) lut_n6359 (.I0(n6330), .I1(n6338), .I2(n6339), .O(n6359));
  LUT3 #(.INIT(8'hE8)) lut_n6360 (.I0(n6350), .I1(n6358), .I2(n6359), .O(n6360));
  LUT3 #(.INIT(8'h96)) lut_n6361 (.I0(x1080), .I1(x1081), .I2(x1082), .O(n6361));
  LUT5 #(.INIT(32'h96696996)) lut_n6362 (.I0(x1071), .I1(x1072), .I2(x1073), .I3(n6354), .I4(n6355), .O(n6362));
  LUT5 #(.INIT(32'hFF969600)) lut_n6363 (.I0(x1077), .I1(x1078), .I2(x1079), .I3(n6361), .I4(n6362), .O(n6363));
  LUT3 #(.INIT(8'h96)) lut_n6364 (.I0(x1086), .I1(x1087), .I2(x1088), .O(n6364));
  LUT5 #(.INIT(32'h96696996)) lut_n6365 (.I0(x1077), .I1(x1078), .I2(x1079), .I3(n6361), .I4(n6362), .O(n6365));
  LUT5 #(.INIT(32'hFF969600)) lut_n6366 (.I0(x1083), .I1(x1084), .I2(x1085), .I3(n6364), .I4(n6365), .O(n6366));
  LUT3 #(.INIT(8'h96)) lut_n6367 (.I0(n6353), .I1(n6356), .I2(n6357), .O(n6367));
  LUT3 #(.INIT(8'hE8)) lut_n6368 (.I0(n6363), .I1(n6366), .I2(n6367), .O(n6368));
  LUT3 #(.INIT(8'h96)) lut_n6369 (.I0(x1092), .I1(x1093), .I2(x1094), .O(n6369));
  LUT5 #(.INIT(32'h96696996)) lut_n6370 (.I0(x1083), .I1(x1084), .I2(x1085), .I3(n6364), .I4(n6365), .O(n6370));
  LUT5 #(.INIT(32'hFF969600)) lut_n6371 (.I0(x1089), .I1(x1090), .I2(x1091), .I3(n6369), .I4(n6370), .O(n6371));
  LUT3 #(.INIT(8'h96)) lut_n6372 (.I0(x1098), .I1(x1099), .I2(x1100), .O(n6372));
  LUT5 #(.INIT(32'h96696996)) lut_n6373 (.I0(x1089), .I1(x1090), .I2(x1091), .I3(n6369), .I4(n6370), .O(n6373));
  LUT5 #(.INIT(32'hFF969600)) lut_n6374 (.I0(x1095), .I1(x1096), .I2(x1097), .I3(n6372), .I4(n6373), .O(n6374));
  LUT3 #(.INIT(8'h96)) lut_n6375 (.I0(n6363), .I1(n6366), .I2(n6367), .O(n6375));
  LUT3 #(.INIT(8'hE8)) lut_n6376 (.I0(n6371), .I1(n6374), .I2(n6375), .O(n6376));
  LUT3 #(.INIT(8'h96)) lut_n6377 (.I0(n6350), .I1(n6358), .I2(n6359), .O(n6377));
  LUT3 #(.INIT(8'hE8)) lut_n6378 (.I0(n6368), .I1(n6376), .I2(n6377), .O(n6378));
  LUT3 #(.INIT(8'h96)) lut_n6379 (.I0(n6322), .I1(n6340), .I2(n6341), .O(n6379));
  LUT3 #(.INIT(8'hE8)) lut_n6380 (.I0(n6360), .I1(n6378), .I2(n6379), .O(n6380));
  LUT3 #(.INIT(8'h96)) lut_n6381 (.I0(n6264), .I1(n6302), .I2(n6303), .O(n6381));
  LUT3 #(.INIT(8'hE8)) lut_n6382 (.I0(n6342), .I1(n6380), .I2(n6381), .O(n6382));
  LUT3 #(.INIT(8'h96)) lut_n6383 (.I0(n6142), .I1(n6220), .I2(n6221), .O(n6383));
  LUT3 #(.INIT(8'hE8)) lut_n6384 (.I0(n6304), .I1(n6382), .I2(n6383), .O(n6384));
  LUT3 #(.INIT(8'h96)) lut_n6385 (.I0(x1104), .I1(x1105), .I2(x1106), .O(n6385));
  LUT5 #(.INIT(32'h96696996)) lut_n6386 (.I0(x1095), .I1(x1096), .I2(x1097), .I3(n6372), .I4(n6373), .O(n6386));
  LUT5 #(.INIT(32'hFF969600)) lut_n6387 (.I0(x1101), .I1(x1102), .I2(x1103), .I3(n6385), .I4(n6386), .O(n6387));
  LUT3 #(.INIT(8'h96)) lut_n6388 (.I0(x1110), .I1(x1111), .I2(x1112), .O(n6388));
  LUT5 #(.INIT(32'h96696996)) lut_n6389 (.I0(x1101), .I1(x1102), .I2(x1103), .I3(n6385), .I4(n6386), .O(n6389));
  LUT5 #(.INIT(32'hFF969600)) lut_n6390 (.I0(x1107), .I1(x1108), .I2(x1109), .I3(n6388), .I4(n6389), .O(n6390));
  LUT3 #(.INIT(8'h96)) lut_n6391 (.I0(n6371), .I1(n6374), .I2(n6375), .O(n6391));
  LUT3 #(.INIT(8'hE8)) lut_n6392 (.I0(n6387), .I1(n6390), .I2(n6391), .O(n6392));
  LUT3 #(.INIT(8'h96)) lut_n6393 (.I0(x1116), .I1(x1117), .I2(x1118), .O(n6393));
  LUT5 #(.INIT(32'h96696996)) lut_n6394 (.I0(x1107), .I1(x1108), .I2(x1109), .I3(n6388), .I4(n6389), .O(n6394));
  LUT5 #(.INIT(32'hFF969600)) lut_n6395 (.I0(x1113), .I1(x1114), .I2(x1115), .I3(n6393), .I4(n6394), .O(n6395));
  LUT3 #(.INIT(8'h96)) lut_n6396 (.I0(x1122), .I1(x1123), .I2(x1124), .O(n6396));
  LUT5 #(.INIT(32'h96696996)) lut_n6397 (.I0(x1113), .I1(x1114), .I2(x1115), .I3(n6393), .I4(n6394), .O(n6397));
  LUT5 #(.INIT(32'hFF969600)) lut_n6398 (.I0(x1119), .I1(x1120), .I2(x1121), .I3(n6396), .I4(n6397), .O(n6398));
  LUT3 #(.INIT(8'h96)) lut_n6399 (.I0(n6387), .I1(n6390), .I2(n6391), .O(n6399));
  LUT3 #(.INIT(8'hE8)) lut_n6400 (.I0(n6395), .I1(n6398), .I2(n6399), .O(n6400));
  LUT3 #(.INIT(8'h96)) lut_n6401 (.I0(n6368), .I1(n6376), .I2(n6377), .O(n6401));
  LUT3 #(.INIT(8'hE8)) lut_n6402 (.I0(n6392), .I1(n6400), .I2(n6401), .O(n6402));
  LUT3 #(.INIT(8'h96)) lut_n6403 (.I0(x1128), .I1(x1129), .I2(x1130), .O(n6403));
  LUT5 #(.INIT(32'h96696996)) lut_n6404 (.I0(x1119), .I1(x1120), .I2(x1121), .I3(n6396), .I4(n6397), .O(n6404));
  LUT5 #(.INIT(32'hFF969600)) lut_n6405 (.I0(x1125), .I1(x1126), .I2(x1127), .I3(n6403), .I4(n6404), .O(n6405));
  LUT3 #(.INIT(8'h96)) lut_n6406 (.I0(x1134), .I1(x1135), .I2(x1136), .O(n6406));
  LUT5 #(.INIT(32'h96696996)) lut_n6407 (.I0(x1125), .I1(x1126), .I2(x1127), .I3(n6403), .I4(n6404), .O(n6407));
  LUT5 #(.INIT(32'hFF969600)) lut_n6408 (.I0(x1131), .I1(x1132), .I2(x1133), .I3(n6406), .I4(n6407), .O(n6408));
  LUT3 #(.INIT(8'h96)) lut_n6409 (.I0(n6395), .I1(n6398), .I2(n6399), .O(n6409));
  LUT3 #(.INIT(8'hE8)) lut_n6410 (.I0(n6405), .I1(n6408), .I2(n6409), .O(n6410));
  LUT3 #(.INIT(8'h96)) lut_n6411 (.I0(x1140), .I1(x1141), .I2(x1142), .O(n6411));
  LUT5 #(.INIT(32'h96696996)) lut_n6412 (.I0(x1131), .I1(x1132), .I2(x1133), .I3(n6406), .I4(n6407), .O(n6412));
  LUT5 #(.INIT(32'hFF969600)) lut_n6413 (.I0(x1137), .I1(x1138), .I2(x1139), .I3(n6411), .I4(n6412), .O(n6413));
  LUT3 #(.INIT(8'h96)) lut_n6414 (.I0(x1146), .I1(x1147), .I2(x1148), .O(n6414));
  LUT5 #(.INIT(32'h96696996)) lut_n6415 (.I0(x1137), .I1(x1138), .I2(x1139), .I3(n6411), .I4(n6412), .O(n6415));
  LUT5 #(.INIT(32'hFF969600)) lut_n6416 (.I0(x1143), .I1(x1144), .I2(x1145), .I3(n6414), .I4(n6415), .O(n6416));
  LUT3 #(.INIT(8'h96)) lut_n6417 (.I0(n6405), .I1(n6408), .I2(n6409), .O(n6417));
  LUT3 #(.INIT(8'hE8)) lut_n6418 (.I0(n6413), .I1(n6416), .I2(n6417), .O(n6418));
  LUT3 #(.INIT(8'h96)) lut_n6419 (.I0(n6392), .I1(n6400), .I2(n6401), .O(n6419));
  LUT3 #(.INIT(8'hE8)) lut_n6420 (.I0(n6410), .I1(n6418), .I2(n6419), .O(n6420));
  LUT3 #(.INIT(8'h96)) lut_n6421 (.I0(n6360), .I1(n6378), .I2(n6379), .O(n6421));
  LUT3 #(.INIT(8'hE8)) lut_n6422 (.I0(n6402), .I1(n6420), .I2(n6421), .O(n6422));
  LUT3 #(.INIT(8'h96)) lut_n6423 (.I0(x1152), .I1(x1153), .I2(x1154), .O(n6423));
  LUT5 #(.INIT(32'h96696996)) lut_n6424 (.I0(x1143), .I1(x1144), .I2(x1145), .I3(n6414), .I4(n6415), .O(n6424));
  LUT5 #(.INIT(32'hFF969600)) lut_n6425 (.I0(x1149), .I1(x1150), .I2(x1151), .I3(n6423), .I4(n6424), .O(n6425));
  LUT3 #(.INIT(8'h96)) lut_n6426 (.I0(x1158), .I1(x1159), .I2(x1160), .O(n6426));
  LUT5 #(.INIT(32'h96696996)) lut_n6427 (.I0(x1149), .I1(x1150), .I2(x1151), .I3(n6423), .I4(n6424), .O(n6427));
  LUT5 #(.INIT(32'hFF969600)) lut_n6428 (.I0(x1155), .I1(x1156), .I2(x1157), .I3(n6426), .I4(n6427), .O(n6428));
  LUT3 #(.INIT(8'h96)) lut_n6429 (.I0(n6413), .I1(n6416), .I2(n6417), .O(n6429));
  LUT3 #(.INIT(8'hE8)) lut_n6430 (.I0(n6425), .I1(n6428), .I2(n6429), .O(n6430));
  LUT3 #(.INIT(8'h96)) lut_n6431 (.I0(x1164), .I1(x1165), .I2(x1166), .O(n6431));
  LUT5 #(.INIT(32'h96696996)) lut_n6432 (.I0(x1155), .I1(x1156), .I2(x1157), .I3(n6426), .I4(n6427), .O(n6432));
  LUT5 #(.INIT(32'hFF969600)) lut_n6433 (.I0(x1161), .I1(x1162), .I2(x1163), .I3(n6431), .I4(n6432), .O(n6433));
  LUT3 #(.INIT(8'h96)) lut_n6434 (.I0(x1170), .I1(x1171), .I2(x1172), .O(n6434));
  LUT5 #(.INIT(32'h96696996)) lut_n6435 (.I0(x1161), .I1(x1162), .I2(x1163), .I3(n6431), .I4(n6432), .O(n6435));
  LUT5 #(.INIT(32'hFF969600)) lut_n6436 (.I0(x1167), .I1(x1168), .I2(x1169), .I3(n6434), .I4(n6435), .O(n6436));
  LUT3 #(.INIT(8'h96)) lut_n6437 (.I0(n6425), .I1(n6428), .I2(n6429), .O(n6437));
  LUT3 #(.INIT(8'hE8)) lut_n6438 (.I0(n6433), .I1(n6436), .I2(n6437), .O(n6438));
  LUT3 #(.INIT(8'h96)) lut_n6439 (.I0(n6410), .I1(n6418), .I2(n6419), .O(n6439));
  LUT3 #(.INIT(8'hE8)) lut_n6440 (.I0(n6430), .I1(n6438), .I2(n6439), .O(n6440));
  LUT3 #(.INIT(8'h96)) lut_n6441 (.I0(x1176), .I1(x1177), .I2(x1178), .O(n6441));
  LUT5 #(.INIT(32'h96696996)) lut_n6442 (.I0(x1167), .I1(x1168), .I2(x1169), .I3(n6434), .I4(n6435), .O(n6442));
  LUT5 #(.INIT(32'hFF969600)) lut_n6443 (.I0(x1173), .I1(x1174), .I2(x1175), .I3(n6441), .I4(n6442), .O(n6443));
  LUT3 #(.INIT(8'h96)) lut_n6444 (.I0(x1182), .I1(x1183), .I2(x1184), .O(n6444));
  LUT5 #(.INIT(32'h96696996)) lut_n6445 (.I0(x1173), .I1(x1174), .I2(x1175), .I3(n6441), .I4(n6442), .O(n6445));
  LUT5 #(.INIT(32'hFF969600)) lut_n6446 (.I0(x1179), .I1(x1180), .I2(x1181), .I3(n6444), .I4(n6445), .O(n6446));
  LUT3 #(.INIT(8'h96)) lut_n6447 (.I0(n6433), .I1(n6436), .I2(n6437), .O(n6447));
  LUT3 #(.INIT(8'hE8)) lut_n6448 (.I0(n6443), .I1(n6446), .I2(n6447), .O(n6448));
  LUT3 #(.INIT(8'h96)) lut_n6449 (.I0(x1188), .I1(x1189), .I2(x1190), .O(n6449));
  LUT5 #(.INIT(32'h96696996)) lut_n6450 (.I0(x1179), .I1(x1180), .I2(x1181), .I3(n6444), .I4(n6445), .O(n6450));
  LUT5 #(.INIT(32'hFF969600)) lut_n6451 (.I0(x1185), .I1(x1186), .I2(x1187), .I3(n6449), .I4(n6450), .O(n6451));
  LUT3 #(.INIT(8'h96)) lut_n6452 (.I0(x1194), .I1(x1195), .I2(x1196), .O(n6452));
  LUT5 #(.INIT(32'h96696996)) lut_n6453 (.I0(x1185), .I1(x1186), .I2(x1187), .I3(n6449), .I4(n6450), .O(n6453));
  LUT5 #(.INIT(32'hFF969600)) lut_n6454 (.I0(x1191), .I1(x1192), .I2(x1193), .I3(n6452), .I4(n6453), .O(n6454));
  LUT3 #(.INIT(8'h96)) lut_n6455 (.I0(n6443), .I1(n6446), .I2(n6447), .O(n6455));
  LUT3 #(.INIT(8'hE8)) lut_n6456 (.I0(n6451), .I1(n6454), .I2(n6455), .O(n6456));
  LUT3 #(.INIT(8'h96)) lut_n6457 (.I0(n6430), .I1(n6438), .I2(n6439), .O(n6457));
  LUT3 #(.INIT(8'hE8)) lut_n6458 (.I0(n6448), .I1(n6456), .I2(n6457), .O(n6458));
  LUT3 #(.INIT(8'h96)) lut_n6459 (.I0(n6402), .I1(n6420), .I2(n6421), .O(n6459));
  LUT3 #(.INIT(8'hE8)) lut_n6460 (.I0(n6440), .I1(n6458), .I2(n6459), .O(n6460));
  LUT3 #(.INIT(8'h96)) lut_n6461 (.I0(n6342), .I1(n6380), .I2(n6381), .O(n6461));
  LUT3 #(.INIT(8'hE8)) lut_n6462 (.I0(n6422), .I1(n6460), .I2(n6461), .O(n6462));
  LUT3 #(.INIT(8'h96)) lut_n6463 (.I0(x1200), .I1(x1201), .I2(x1202), .O(n6463));
  LUT5 #(.INIT(32'h96696996)) lut_n6464 (.I0(x1191), .I1(x1192), .I2(x1193), .I3(n6452), .I4(n6453), .O(n6464));
  LUT5 #(.INIT(32'hFF969600)) lut_n6465 (.I0(x1197), .I1(x1198), .I2(x1199), .I3(n6463), .I4(n6464), .O(n6465));
  LUT3 #(.INIT(8'h96)) lut_n6466 (.I0(x1206), .I1(x1207), .I2(x1208), .O(n6466));
  LUT5 #(.INIT(32'h96696996)) lut_n6467 (.I0(x1197), .I1(x1198), .I2(x1199), .I3(n6463), .I4(n6464), .O(n6467));
  LUT5 #(.INIT(32'hFF969600)) lut_n6468 (.I0(x1203), .I1(x1204), .I2(x1205), .I3(n6466), .I4(n6467), .O(n6468));
  LUT3 #(.INIT(8'h96)) lut_n6469 (.I0(n6451), .I1(n6454), .I2(n6455), .O(n6469));
  LUT3 #(.INIT(8'hE8)) lut_n6470 (.I0(n6465), .I1(n6468), .I2(n6469), .O(n6470));
  LUT3 #(.INIT(8'h96)) lut_n6471 (.I0(x1212), .I1(x1213), .I2(x1214), .O(n6471));
  LUT5 #(.INIT(32'h96696996)) lut_n6472 (.I0(x1203), .I1(x1204), .I2(x1205), .I3(n6466), .I4(n6467), .O(n6472));
  LUT5 #(.INIT(32'hFF969600)) lut_n6473 (.I0(x1209), .I1(x1210), .I2(x1211), .I3(n6471), .I4(n6472), .O(n6473));
  LUT3 #(.INIT(8'h96)) lut_n6474 (.I0(x1218), .I1(x1219), .I2(x1220), .O(n6474));
  LUT5 #(.INIT(32'h96696996)) lut_n6475 (.I0(x1209), .I1(x1210), .I2(x1211), .I3(n6471), .I4(n6472), .O(n6475));
  LUT5 #(.INIT(32'hFF969600)) lut_n6476 (.I0(x1215), .I1(x1216), .I2(x1217), .I3(n6474), .I4(n6475), .O(n6476));
  LUT3 #(.INIT(8'h96)) lut_n6477 (.I0(n6465), .I1(n6468), .I2(n6469), .O(n6477));
  LUT3 #(.INIT(8'hE8)) lut_n6478 (.I0(n6473), .I1(n6476), .I2(n6477), .O(n6478));
  LUT3 #(.INIT(8'h96)) lut_n6479 (.I0(n6448), .I1(n6456), .I2(n6457), .O(n6479));
  LUT3 #(.INIT(8'hE8)) lut_n6480 (.I0(n6470), .I1(n6478), .I2(n6479), .O(n6480));
  LUT3 #(.INIT(8'h96)) lut_n6481 (.I0(x1224), .I1(x1225), .I2(x1226), .O(n6481));
  LUT5 #(.INIT(32'h96696996)) lut_n6482 (.I0(x1215), .I1(x1216), .I2(x1217), .I3(n6474), .I4(n6475), .O(n6482));
  LUT5 #(.INIT(32'hFF969600)) lut_n6483 (.I0(x1221), .I1(x1222), .I2(x1223), .I3(n6481), .I4(n6482), .O(n6483));
  LUT3 #(.INIT(8'h96)) lut_n6484 (.I0(x1230), .I1(x1231), .I2(x1232), .O(n6484));
  LUT5 #(.INIT(32'h96696996)) lut_n6485 (.I0(x1221), .I1(x1222), .I2(x1223), .I3(n6481), .I4(n6482), .O(n6485));
  LUT5 #(.INIT(32'hFF969600)) lut_n6486 (.I0(x1227), .I1(x1228), .I2(x1229), .I3(n6484), .I4(n6485), .O(n6486));
  LUT3 #(.INIT(8'h96)) lut_n6487 (.I0(n6473), .I1(n6476), .I2(n6477), .O(n6487));
  LUT3 #(.INIT(8'hE8)) lut_n6488 (.I0(n6483), .I1(n6486), .I2(n6487), .O(n6488));
  LUT3 #(.INIT(8'h96)) lut_n6489 (.I0(x1236), .I1(x1237), .I2(x1238), .O(n6489));
  LUT5 #(.INIT(32'h96696996)) lut_n6490 (.I0(x1227), .I1(x1228), .I2(x1229), .I3(n6484), .I4(n6485), .O(n6490));
  LUT5 #(.INIT(32'hFF969600)) lut_n6491 (.I0(x1233), .I1(x1234), .I2(x1235), .I3(n6489), .I4(n6490), .O(n6491));
  LUT3 #(.INIT(8'h96)) lut_n6492 (.I0(x1242), .I1(x1243), .I2(x1244), .O(n6492));
  LUT5 #(.INIT(32'h96696996)) lut_n6493 (.I0(x1233), .I1(x1234), .I2(x1235), .I3(n6489), .I4(n6490), .O(n6493));
  LUT5 #(.INIT(32'hFF969600)) lut_n6494 (.I0(x1239), .I1(x1240), .I2(x1241), .I3(n6492), .I4(n6493), .O(n6494));
  LUT3 #(.INIT(8'h96)) lut_n6495 (.I0(n6483), .I1(n6486), .I2(n6487), .O(n6495));
  LUT3 #(.INIT(8'hE8)) lut_n6496 (.I0(n6491), .I1(n6494), .I2(n6495), .O(n6496));
  LUT3 #(.INIT(8'h96)) lut_n6497 (.I0(n6470), .I1(n6478), .I2(n6479), .O(n6497));
  LUT3 #(.INIT(8'hE8)) lut_n6498 (.I0(n6488), .I1(n6496), .I2(n6497), .O(n6498));
  LUT3 #(.INIT(8'h96)) lut_n6499 (.I0(n6440), .I1(n6458), .I2(n6459), .O(n6499));
  LUT3 #(.INIT(8'hE8)) lut_n6500 (.I0(n6480), .I1(n6498), .I2(n6499), .O(n6500));
  LUT3 #(.INIT(8'h96)) lut_n6501 (.I0(x1248), .I1(x1249), .I2(x1250), .O(n6501));
  LUT5 #(.INIT(32'h96696996)) lut_n6502 (.I0(x1239), .I1(x1240), .I2(x1241), .I3(n6492), .I4(n6493), .O(n6502));
  LUT5 #(.INIT(32'hFF969600)) lut_n6503 (.I0(x1245), .I1(x1246), .I2(x1247), .I3(n6501), .I4(n6502), .O(n6503));
  LUT3 #(.INIT(8'h96)) lut_n6504 (.I0(x1254), .I1(x1255), .I2(x1256), .O(n6504));
  LUT5 #(.INIT(32'h96696996)) lut_n6505 (.I0(x1245), .I1(x1246), .I2(x1247), .I3(n6501), .I4(n6502), .O(n6505));
  LUT5 #(.INIT(32'hFF969600)) lut_n6506 (.I0(x1251), .I1(x1252), .I2(x1253), .I3(n6504), .I4(n6505), .O(n6506));
  LUT3 #(.INIT(8'h96)) lut_n6507 (.I0(n6491), .I1(n6494), .I2(n6495), .O(n6507));
  LUT3 #(.INIT(8'hE8)) lut_n6508 (.I0(n6503), .I1(n6506), .I2(n6507), .O(n6508));
  LUT3 #(.INIT(8'h96)) lut_n6509 (.I0(x1260), .I1(x1261), .I2(x1262), .O(n6509));
  LUT5 #(.INIT(32'h96696996)) lut_n6510 (.I0(x1251), .I1(x1252), .I2(x1253), .I3(n6504), .I4(n6505), .O(n6510));
  LUT5 #(.INIT(32'hFF969600)) lut_n6511 (.I0(x1257), .I1(x1258), .I2(x1259), .I3(n6509), .I4(n6510), .O(n6511));
  LUT3 #(.INIT(8'h96)) lut_n6512 (.I0(x1266), .I1(x1267), .I2(x1268), .O(n6512));
  LUT5 #(.INIT(32'h96696996)) lut_n6513 (.I0(x1257), .I1(x1258), .I2(x1259), .I3(n6509), .I4(n6510), .O(n6513));
  LUT5 #(.INIT(32'hFF969600)) lut_n6514 (.I0(x1263), .I1(x1264), .I2(x1265), .I3(n6512), .I4(n6513), .O(n6514));
  LUT3 #(.INIT(8'h96)) lut_n6515 (.I0(n6503), .I1(n6506), .I2(n6507), .O(n6515));
  LUT3 #(.INIT(8'hE8)) lut_n6516 (.I0(n6511), .I1(n6514), .I2(n6515), .O(n6516));
  LUT3 #(.INIT(8'h96)) lut_n6517 (.I0(n6488), .I1(n6496), .I2(n6497), .O(n6517));
  LUT3 #(.INIT(8'hE8)) lut_n6518 (.I0(n6508), .I1(n6516), .I2(n6517), .O(n6518));
  LUT3 #(.INIT(8'h96)) lut_n6519 (.I0(x1272), .I1(x1273), .I2(x1274), .O(n6519));
  LUT5 #(.INIT(32'h96696996)) lut_n6520 (.I0(x1263), .I1(x1264), .I2(x1265), .I3(n6512), .I4(n6513), .O(n6520));
  LUT5 #(.INIT(32'hFF969600)) lut_n6521 (.I0(x1269), .I1(x1270), .I2(x1271), .I3(n6519), .I4(n6520), .O(n6521));
  LUT3 #(.INIT(8'h96)) lut_n6522 (.I0(x1278), .I1(x1279), .I2(x1280), .O(n6522));
  LUT5 #(.INIT(32'h96696996)) lut_n6523 (.I0(x1269), .I1(x1270), .I2(x1271), .I3(n6519), .I4(n6520), .O(n6523));
  LUT5 #(.INIT(32'hFF969600)) lut_n6524 (.I0(x1275), .I1(x1276), .I2(x1277), .I3(n6522), .I4(n6523), .O(n6524));
  LUT3 #(.INIT(8'h96)) lut_n6525 (.I0(n6511), .I1(n6514), .I2(n6515), .O(n6525));
  LUT3 #(.INIT(8'hE8)) lut_n6526 (.I0(n6521), .I1(n6524), .I2(n6525), .O(n6526));
  LUT3 #(.INIT(8'h96)) lut_n6527 (.I0(x1284), .I1(x1285), .I2(x1286), .O(n6527));
  LUT5 #(.INIT(32'h96696996)) lut_n6528 (.I0(x1275), .I1(x1276), .I2(x1277), .I3(n6522), .I4(n6523), .O(n6528));
  LUT5 #(.INIT(32'hFF969600)) lut_n6529 (.I0(x1281), .I1(x1282), .I2(x1283), .I3(n6527), .I4(n6528), .O(n6529));
  LUT3 #(.INIT(8'h96)) lut_n6530 (.I0(x1290), .I1(x1291), .I2(x1292), .O(n6530));
  LUT5 #(.INIT(32'h96696996)) lut_n6531 (.I0(x1281), .I1(x1282), .I2(x1283), .I3(n6527), .I4(n6528), .O(n6531));
  LUT5 #(.INIT(32'hFF969600)) lut_n6532 (.I0(x1287), .I1(x1288), .I2(x1289), .I3(n6530), .I4(n6531), .O(n6532));
  LUT3 #(.INIT(8'h96)) lut_n6533 (.I0(n6521), .I1(n6524), .I2(n6525), .O(n6533));
  LUT3 #(.INIT(8'hE8)) lut_n6534 (.I0(n6529), .I1(n6532), .I2(n6533), .O(n6534));
  LUT3 #(.INIT(8'h96)) lut_n6535 (.I0(n6508), .I1(n6516), .I2(n6517), .O(n6535));
  LUT3 #(.INIT(8'hE8)) lut_n6536 (.I0(n6526), .I1(n6534), .I2(n6535), .O(n6536));
  LUT3 #(.INIT(8'h96)) lut_n6537 (.I0(n6480), .I1(n6498), .I2(n6499), .O(n6537));
  LUT3 #(.INIT(8'hE8)) lut_n6538 (.I0(n6518), .I1(n6536), .I2(n6537), .O(n6538));
  LUT3 #(.INIT(8'h96)) lut_n6539 (.I0(n6422), .I1(n6460), .I2(n6461), .O(n6539));
  LUT3 #(.INIT(8'hE8)) lut_n6540 (.I0(n6500), .I1(n6538), .I2(n6539), .O(n6540));
  LUT3 #(.INIT(8'h96)) lut_n6541 (.I0(n6304), .I1(n6382), .I2(n6383), .O(n6541));
  LUT3 #(.INIT(8'hE8)) lut_n6542 (.I0(n6462), .I1(n6540), .I2(n6541), .O(n6542));
  LUT3 #(.INIT(8'h96)) lut_n6543 (.I0(n6064), .I1(n6222), .I2(n6223), .O(n6543));
  LUT3 #(.INIT(8'hE8)) lut_n6544 (.I0(n6384), .I1(n6542), .I2(n6543), .O(n6544));
  LUT3 #(.INIT(8'h96)) lut_n6545 (.I0(x1296), .I1(x1297), .I2(x1298), .O(n6545));
  LUT5 #(.INIT(32'h96696996)) lut_n6546 (.I0(x1287), .I1(x1288), .I2(x1289), .I3(n6530), .I4(n6531), .O(n6546));
  LUT5 #(.INIT(32'hFF969600)) lut_n6547 (.I0(x1293), .I1(x1294), .I2(x1295), .I3(n6545), .I4(n6546), .O(n6547));
  LUT3 #(.INIT(8'h96)) lut_n6548 (.I0(x1302), .I1(x1303), .I2(x1304), .O(n6548));
  LUT5 #(.INIT(32'h96696996)) lut_n6549 (.I0(x1293), .I1(x1294), .I2(x1295), .I3(n6545), .I4(n6546), .O(n6549));
  LUT5 #(.INIT(32'hFF969600)) lut_n6550 (.I0(x1299), .I1(x1300), .I2(x1301), .I3(n6548), .I4(n6549), .O(n6550));
  LUT3 #(.INIT(8'h96)) lut_n6551 (.I0(n6529), .I1(n6532), .I2(n6533), .O(n6551));
  LUT3 #(.INIT(8'hE8)) lut_n6552 (.I0(n6547), .I1(n6550), .I2(n6551), .O(n6552));
  LUT3 #(.INIT(8'h96)) lut_n6553 (.I0(x1308), .I1(x1309), .I2(x1310), .O(n6553));
  LUT5 #(.INIT(32'h96696996)) lut_n6554 (.I0(x1299), .I1(x1300), .I2(x1301), .I3(n6548), .I4(n6549), .O(n6554));
  LUT5 #(.INIT(32'hFF969600)) lut_n6555 (.I0(x1305), .I1(x1306), .I2(x1307), .I3(n6553), .I4(n6554), .O(n6555));
  LUT3 #(.INIT(8'h96)) lut_n6556 (.I0(x1314), .I1(x1315), .I2(x1316), .O(n6556));
  LUT5 #(.INIT(32'h96696996)) lut_n6557 (.I0(x1305), .I1(x1306), .I2(x1307), .I3(n6553), .I4(n6554), .O(n6557));
  LUT5 #(.INIT(32'hFF969600)) lut_n6558 (.I0(x1311), .I1(x1312), .I2(x1313), .I3(n6556), .I4(n6557), .O(n6558));
  LUT3 #(.INIT(8'h96)) lut_n6559 (.I0(n6547), .I1(n6550), .I2(n6551), .O(n6559));
  LUT3 #(.INIT(8'hE8)) lut_n6560 (.I0(n6555), .I1(n6558), .I2(n6559), .O(n6560));
  LUT3 #(.INIT(8'h96)) lut_n6561 (.I0(n6526), .I1(n6534), .I2(n6535), .O(n6561));
  LUT3 #(.INIT(8'hE8)) lut_n6562 (.I0(n6552), .I1(n6560), .I2(n6561), .O(n6562));
  LUT3 #(.INIT(8'h96)) lut_n6563 (.I0(x1320), .I1(x1321), .I2(x1322), .O(n6563));
  LUT5 #(.INIT(32'h96696996)) lut_n6564 (.I0(x1311), .I1(x1312), .I2(x1313), .I3(n6556), .I4(n6557), .O(n6564));
  LUT5 #(.INIT(32'hFF969600)) lut_n6565 (.I0(x1317), .I1(x1318), .I2(x1319), .I3(n6563), .I4(n6564), .O(n6565));
  LUT3 #(.INIT(8'h96)) lut_n6566 (.I0(x1326), .I1(x1327), .I2(x1328), .O(n6566));
  LUT5 #(.INIT(32'h96696996)) lut_n6567 (.I0(x1317), .I1(x1318), .I2(x1319), .I3(n6563), .I4(n6564), .O(n6567));
  LUT5 #(.INIT(32'hFF969600)) lut_n6568 (.I0(x1323), .I1(x1324), .I2(x1325), .I3(n6566), .I4(n6567), .O(n6568));
  LUT3 #(.INIT(8'h96)) lut_n6569 (.I0(n6555), .I1(n6558), .I2(n6559), .O(n6569));
  LUT3 #(.INIT(8'hE8)) lut_n6570 (.I0(n6565), .I1(n6568), .I2(n6569), .O(n6570));
  LUT3 #(.INIT(8'h96)) lut_n6571 (.I0(x1332), .I1(x1333), .I2(x1334), .O(n6571));
  LUT5 #(.INIT(32'h96696996)) lut_n6572 (.I0(x1323), .I1(x1324), .I2(x1325), .I3(n6566), .I4(n6567), .O(n6572));
  LUT5 #(.INIT(32'hFF969600)) lut_n6573 (.I0(x1329), .I1(x1330), .I2(x1331), .I3(n6571), .I4(n6572), .O(n6573));
  LUT3 #(.INIT(8'h96)) lut_n6574 (.I0(x1338), .I1(x1339), .I2(x1340), .O(n6574));
  LUT5 #(.INIT(32'h96696996)) lut_n6575 (.I0(x1329), .I1(x1330), .I2(x1331), .I3(n6571), .I4(n6572), .O(n6575));
  LUT5 #(.INIT(32'hFF969600)) lut_n6576 (.I0(x1335), .I1(x1336), .I2(x1337), .I3(n6574), .I4(n6575), .O(n6576));
  LUT3 #(.INIT(8'h96)) lut_n6577 (.I0(n6565), .I1(n6568), .I2(n6569), .O(n6577));
  LUT3 #(.INIT(8'hE8)) lut_n6578 (.I0(n6573), .I1(n6576), .I2(n6577), .O(n6578));
  LUT3 #(.INIT(8'h96)) lut_n6579 (.I0(n6552), .I1(n6560), .I2(n6561), .O(n6579));
  LUT3 #(.INIT(8'hE8)) lut_n6580 (.I0(n6570), .I1(n6578), .I2(n6579), .O(n6580));
  LUT3 #(.INIT(8'h96)) lut_n6581 (.I0(n6518), .I1(n6536), .I2(n6537), .O(n6581));
  LUT3 #(.INIT(8'hE8)) lut_n6582 (.I0(n6562), .I1(n6580), .I2(n6581), .O(n6582));
  LUT3 #(.INIT(8'h96)) lut_n6583 (.I0(x1344), .I1(x1345), .I2(x1346), .O(n6583));
  LUT5 #(.INIT(32'h96696996)) lut_n6584 (.I0(x1335), .I1(x1336), .I2(x1337), .I3(n6574), .I4(n6575), .O(n6584));
  LUT5 #(.INIT(32'hFF969600)) lut_n6585 (.I0(x1341), .I1(x1342), .I2(x1343), .I3(n6583), .I4(n6584), .O(n6585));
  LUT3 #(.INIT(8'h96)) lut_n6586 (.I0(x1350), .I1(x1351), .I2(x1352), .O(n6586));
  LUT5 #(.INIT(32'h96696996)) lut_n6587 (.I0(x1341), .I1(x1342), .I2(x1343), .I3(n6583), .I4(n6584), .O(n6587));
  LUT5 #(.INIT(32'hFF969600)) lut_n6588 (.I0(x1347), .I1(x1348), .I2(x1349), .I3(n6586), .I4(n6587), .O(n6588));
  LUT3 #(.INIT(8'h96)) lut_n6589 (.I0(n6573), .I1(n6576), .I2(n6577), .O(n6589));
  LUT3 #(.INIT(8'hE8)) lut_n6590 (.I0(n6585), .I1(n6588), .I2(n6589), .O(n6590));
  LUT3 #(.INIT(8'h96)) lut_n6591 (.I0(x1356), .I1(x1357), .I2(x1358), .O(n6591));
  LUT5 #(.INIT(32'h96696996)) lut_n6592 (.I0(x1347), .I1(x1348), .I2(x1349), .I3(n6586), .I4(n6587), .O(n6592));
  LUT5 #(.INIT(32'hFF969600)) lut_n6593 (.I0(x1353), .I1(x1354), .I2(x1355), .I3(n6591), .I4(n6592), .O(n6593));
  LUT3 #(.INIT(8'h96)) lut_n6594 (.I0(x1362), .I1(x1363), .I2(x1364), .O(n6594));
  LUT5 #(.INIT(32'h96696996)) lut_n6595 (.I0(x1353), .I1(x1354), .I2(x1355), .I3(n6591), .I4(n6592), .O(n6595));
  LUT5 #(.INIT(32'hFF969600)) lut_n6596 (.I0(x1359), .I1(x1360), .I2(x1361), .I3(n6594), .I4(n6595), .O(n6596));
  LUT3 #(.INIT(8'h96)) lut_n6597 (.I0(n6585), .I1(n6588), .I2(n6589), .O(n6597));
  LUT3 #(.INIT(8'hE8)) lut_n6598 (.I0(n6593), .I1(n6596), .I2(n6597), .O(n6598));
  LUT3 #(.INIT(8'h96)) lut_n6599 (.I0(n6570), .I1(n6578), .I2(n6579), .O(n6599));
  LUT3 #(.INIT(8'hE8)) lut_n6600 (.I0(n6590), .I1(n6598), .I2(n6599), .O(n6600));
  LUT3 #(.INIT(8'h96)) lut_n6601 (.I0(x1368), .I1(x1369), .I2(x1370), .O(n6601));
  LUT5 #(.INIT(32'h96696996)) lut_n6602 (.I0(x1359), .I1(x1360), .I2(x1361), .I3(n6594), .I4(n6595), .O(n6602));
  LUT5 #(.INIT(32'hFF969600)) lut_n6603 (.I0(x1365), .I1(x1366), .I2(x1367), .I3(n6601), .I4(n6602), .O(n6603));
  LUT3 #(.INIT(8'h96)) lut_n6604 (.I0(x1374), .I1(x1375), .I2(x1376), .O(n6604));
  LUT5 #(.INIT(32'h96696996)) lut_n6605 (.I0(x1365), .I1(x1366), .I2(x1367), .I3(n6601), .I4(n6602), .O(n6605));
  LUT5 #(.INIT(32'hFF969600)) lut_n6606 (.I0(x1371), .I1(x1372), .I2(x1373), .I3(n6604), .I4(n6605), .O(n6606));
  LUT3 #(.INIT(8'h96)) lut_n6607 (.I0(n6593), .I1(n6596), .I2(n6597), .O(n6607));
  LUT3 #(.INIT(8'hE8)) lut_n6608 (.I0(n6603), .I1(n6606), .I2(n6607), .O(n6608));
  LUT3 #(.INIT(8'h96)) lut_n6609 (.I0(x1380), .I1(x1381), .I2(x1382), .O(n6609));
  LUT5 #(.INIT(32'h96696996)) lut_n6610 (.I0(x1371), .I1(x1372), .I2(x1373), .I3(n6604), .I4(n6605), .O(n6610));
  LUT5 #(.INIT(32'hFF969600)) lut_n6611 (.I0(x1377), .I1(x1378), .I2(x1379), .I3(n6609), .I4(n6610), .O(n6611));
  LUT3 #(.INIT(8'h96)) lut_n6612 (.I0(x1386), .I1(x1387), .I2(x1388), .O(n6612));
  LUT5 #(.INIT(32'h96696996)) lut_n6613 (.I0(x1377), .I1(x1378), .I2(x1379), .I3(n6609), .I4(n6610), .O(n6613));
  LUT5 #(.INIT(32'hFF969600)) lut_n6614 (.I0(x1383), .I1(x1384), .I2(x1385), .I3(n6612), .I4(n6613), .O(n6614));
  LUT3 #(.INIT(8'h96)) lut_n6615 (.I0(n6603), .I1(n6606), .I2(n6607), .O(n6615));
  LUT3 #(.INIT(8'hE8)) lut_n6616 (.I0(n6611), .I1(n6614), .I2(n6615), .O(n6616));
  LUT3 #(.INIT(8'h96)) lut_n6617 (.I0(n6590), .I1(n6598), .I2(n6599), .O(n6617));
  LUT3 #(.INIT(8'hE8)) lut_n6618 (.I0(n6608), .I1(n6616), .I2(n6617), .O(n6618));
  LUT3 #(.INIT(8'h96)) lut_n6619 (.I0(n6562), .I1(n6580), .I2(n6581), .O(n6619));
  LUT3 #(.INIT(8'hE8)) lut_n6620 (.I0(n6600), .I1(n6618), .I2(n6619), .O(n6620));
  LUT3 #(.INIT(8'h96)) lut_n6621 (.I0(n6500), .I1(n6538), .I2(n6539), .O(n6621));
  LUT3 #(.INIT(8'hE8)) lut_n6622 (.I0(n6582), .I1(n6620), .I2(n6621), .O(n6622));
  LUT3 #(.INIT(8'h96)) lut_n6623 (.I0(x1392), .I1(x1393), .I2(x1394), .O(n6623));
  LUT5 #(.INIT(32'h96696996)) lut_n6624 (.I0(x1383), .I1(x1384), .I2(x1385), .I3(n6612), .I4(n6613), .O(n6624));
  LUT5 #(.INIT(32'hFF969600)) lut_n6625 (.I0(x1389), .I1(x1390), .I2(x1391), .I3(n6623), .I4(n6624), .O(n6625));
  LUT3 #(.INIT(8'h96)) lut_n6626 (.I0(x1398), .I1(x1399), .I2(x1400), .O(n6626));
  LUT5 #(.INIT(32'h96696996)) lut_n6627 (.I0(x1389), .I1(x1390), .I2(x1391), .I3(n6623), .I4(n6624), .O(n6627));
  LUT5 #(.INIT(32'hFF969600)) lut_n6628 (.I0(x1395), .I1(x1396), .I2(x1397), .I3(n6626), .I4(n6627), .O(n6628));
  LUT3 #(.INIT(8'h96)) lut_n6629 (.I0(n6611), .I1(n6614), .I2(n6615), .O(n6629));
  LUT3 #(.INIT(8'hE8)) lut_n6630 (.I0(n6625), .I1(n6628), .I2(n6629), .O(n6630));
  LUT3 #(.INIT(8'h96)) lut_n6631 (.I0(x1404), .I1(x1405), .I2(x1406), .O(n6631));
  LUT5 #(.INIT(32'h96696996)) lut_n6632 (.I0(x1395), .I1(x1396), .I2(x1397), .I3(n6626), .I4(n6627), .O(n6632));
  LUT5 #(.INIT(32'hFF969600)) lut_n6633 (.I0(x1401), .I1(x1402), .I2(x1403), .I3(n6631), .I4(n6632), .O(n6633));
  LUT3 #(.INIT(8'h96)) lut_n6634 (.I0(x1410), .I1(x1411), .I2(x1412), .O(n6634));
  LUT5 #(.INIT(32'h96696996)) lut_n6635 (.I0(x1401), .I1(x1402), .I2(x1403), .I3(n6631), .I4(n6632), .O(n6635));
  LUT5 #(.INIT(32'hFF969600)) lut_n6636 (.I0(x1407), .I1(x1408), .I2(x1409), .I3(n6634), .I4(n6635), .O(n6636));
  LUT3 #(.INIT(8'h96)) lut_n6637 (.I0(n6625), .I1(n6628), .I2(n6629), .O(n6637));
  LUT3 #(.INIT(8'hE8)) lut_n6638 (.I0(n6633), .I1(n6636), .I2(n6637), .O(n6638));
  LUT3 #(.INIT(8'h96)) lut_n6639 (.I0(n6608), .I1(n6616), .I2(n6617), .O(n6639));
  LUT3 #(.INIT(8'hE8)) lut_n6640 (.I0(n6630), .I1(n6638), .I2(n6639), .O(n6640));
  LUT3 #(.INIT(8'h96)) lut_n6641 (.I0(x1416), .I1(x1417), .I2(x1418), .O(n6641));
  LUT5 #(.INIT(32'h96696996)) lut_n6642 (.I0(x1407), .I1(x1408), .I2(x1409), .I3(n6634), .I4(n6635), .O(n6642));
  LUT5 #(.INIT(32'hFF969600)) lut_n6643 (.I0(x1413), .I1(x1414), .I2(x1415), .I3(n6641), .I4(n6642), .O(n6643));
  LUT3 #(.INIT(8'h96)) lut_n6644 (.I0(x1422), .I1(x1423), .I2(x1424), .O(n6644));
  LUT5 #(.INIT(32'h96696996)) lut_n6645 (.I0(x1413), .I1(x1414), .I2(x1415), .I3(n6641), .I4(n6642), .O(n6645));
  LUT5 #(.INIT(32'hFF969600)) lut_n6646 (.I0(x1419), .I1(x1420), .I2(x1421), .I3(n6644), .I4(n6645), .O(n6646));
  LUT3 #(.INIT(8'h96)) lut_n6647 (.I0(n6633), .I1(n6636), .I2(n6637), .O(n6647));
  LUT3 #(.INIT(8'hE8)) lut_n6648 (.I0(n6643), .I1(n6646), .I2(n6647), .O(n6648));
  LUT3 #(.INIT(8'h96)) lut_n6649 (.I0(x1428), .I1(x1429), .I2(x1430), .O(n6649));
  LUT5 #(.INIT(32'h96696996)) lut_n6650 (.I0(x1419), .I1(x1420), .I2(x1421), .I3(n6644), .I4(n6645), .O(n6650));
  LUT5 #(.INIT(32'hFF969600)) lut_n6651 (.I0(x1425), .I1(x1426), .I2(x1427), .I3(n6649), .I4(n6650), .O(n6651));
  LUT3 #(.INIT(8'h96)) lut_n6652 (.I0(x1434), .I1(x1435), .I2(x1436), .O(n6652));
  LUT5 #(.INIT(32'h96696996)) lut_n6653 (.I0(x1425), .I1(x1426), .I2(x1427), .I3(n6649), .I4(n6650), .O(n6653));
  LUT5 #(.INIT(32'hFF969600)) lut_n6654 (.I0(x1431), .I1(x1432), .I2(x1433), .I3(n6652), .I4(n6653), .O(n6654));
  LUT3 #(.INIT(8'h96)) lut_n6655 (.I0(n6643), .I1(n6646), .I2(n6647), .O(n6655));
  LUT3 #(.INIT(8'hE8)) lut_n6656 (.I0(n6651), .I1(n6654), .I2(n6655), .O(n6656));
  LUT3 #(.INIT(8'h96)) lut_n6657 (.I0(n6630), .I1(n6638), .I2(n6639), .O(n6657));
  LUT3 #(.INIT(8'hE8)) lut_n6658 (.I0(n6648), .I1(n6656), .I2(n6657), .O(n6658));
  LUT3 #(.INIT(8'h96)) lut_n6659 (.I0(n6600), .I1(n6618), .I2(n6619), .O(n6659));
  LUT3 #(.INIT(8'hE8)) lut_n6660 (.I0(n6640), .I1(n6658), .I2(n6659), .O(n6660));
  LUT3 #(.INIT(8'h96)) lut_n6661 (.I0(x1440), .I1(x1441), .I2(x1442), .O(n6661));
  LUT5 #(.INIT(32'h96696996)) lut_n6662 (.I0(x1431), .I1(x1432), .I2(x1433), .I3(n6652), .I4(n6653), .O(n6662));
  LUT5 #(.INIT(32'hFF969600)) lut_n6663 (.I0(x1437), .I1(x1438), .I2(x1439), .I3(n6661), .I4(n6662), .O(n6663));
  LUT3 #(.INIT(8'h96)) lut_n6664 (.I0(x1446), .I1(x1447), .I2(x1448), .O(n6664));
  LUT5 #(.INIT(32'h96696996)) lut_n6665 (.I0(x1437), .I1(x1438), .I2(x1439), .I3(n6661), .I4(n6662), .O(n6665));
  LUT5 #(.INIT(32'hFF969600)) lut_n6666 (.I0(x1443), .I1(x1444), .I2(x1445), .I3(n6664), .I4(n6665), .O(n6666));
  LUT3 #(.INIT(8'h96)) lut_n6667 (.I0(n6651), .I1(n6654), .I2(n6655), .O(n6667));
  LUT3 #(.INIT(8'hE8)) lut_n6668 (.I0(n6663), .I1(n6666), .I2(n6667), .O(n6668));
  LUT3 #(.INIT(8'h96)) lut_n6669 (.I0(x1452), .I1(x1453), .I2(x1454), .O(n6669));
  LUT5 #(.INIT(32'h96696996)) lut_n6670 (.I0(x1443), .I1(x1444), .I2(x1445), .I3(n6664), .I4(n6665), .O(n6670));
  LUT5 #(.INIT(32'hFF969600)) lut_n6671 (.I0(x1449), .I1(x1450), .I2(x1451), .I3(n6669), .I4(n6670), .O(n6671));
  LUT3 #(.INIT(8'h96)) lut_n6672 (.I0(x1458), .I1(x1459), .I2(x1460), .O(n6672));
  LUT5 #(.INIT(32'h96696996)) lut_n6673 (.I0(x1449), .I1(x1450), .I2(x1451), .I3(n6669), .I4(n6670), .O(n6673));
  LUT5 #(.INIT(32'hFF969600)) lut_n6674 (.I0(x1455), .I1(x1456), .I2(x1457), .I3(n6672), .I4(n6673), .O(n6674));
  LUT3 #(.INIT(8'h96)) lut_n6675 (.I0(n6663), .I1(n6666), .I2(n6667), .O(n6675));
  LUT3 #(.INIT(8'hE8)) lut_n6676 (.I0(n6671), .I1(n6674), .I2(n6675), .O(n6676));
  LUT3 #(.INIT(8'h96)) lut_n6677 (.I0(n6648), .I1(n6656), .I2(n6657), .O(n6677));
  LUT3 #(.INIT(8'hE8)) lut_n6678 (.I0(n6668), .I1(n6676), .I2(n6677), .O(n6678));
  LUT3 #(.INIT(8'h96)) lut_n6679 (.I0(x1464), .I1(x1465), .I2(x1466), .O(n6679));
  LUT5 #(.INIT(32'h96696996)) lut_n6680 (.I0(x1455), .I1(x1456), .I2(x1457), .I3(n6672), .I4(n6673), .O(n6680));
  LUT5 #(.INIT(32'hFF969600)) lut_n6681 (.I0(x1461), .I1(x1462), .I2(x1463), .I3(n6679), .I4(n6680), .O(n6681));
  LUT3 #(.INIT(8'h96)) lut_n6682 (.I0(x1470), .I1(x1471), .I2(x1472), .O(n6682));
  LUT5 #(.INIT(32'h96696996)) lut_n6683 (.I0(x1461), .I1(x1462), .I2(x1463), .I3(n6679), .I4(n6680), .O(n6683));
  LUT5 #(.INIT(32'hFF969600)) lut_n6684 (.I0(x1467), .I1(x1468), .I2(x1469), .I3(n6682), .I4(n6683), .O(n6684));
  LUT3 #(.INIT(8'h96)) lut_n6685 (.I0(n6671), .I1(n6674), .I2(n6675), .O(n6685));
  LUT3 #(.INIT(8'hE8)) lut_n6686 (.I0(n6681), .I1(n6684), .I2(n6685), .O(n6686));
  LUT3 #(.INIT(8'h96)) lut_n6687 (.I0(x1476), .I1(x1477), .I2(x1478), .O(n6687));
  LUT5 #(.INIT(32'h96696996)) lut_n6688 (.I0(x1467), .I1(x1468), .I2(x1469), .I3(n6682), .I4(n6683), .O(n6688));
  LUT5 #(.INIT(32'hFF969600)) lut_n6689 (.I0(x1473), .I1(x1474), .I2(x1475), .I3(n6687), .I4(n6688), .O(n6689));
  LUT3 #(.INIT(8'h96)) lut_n6690 (.I0(x1482), .I1(x1483), .I2(x1484), .O(n6690));
  LUT5 #(.INIT(32'h96696996)) lut_n6691 (.I0(x1473), .I1(x1474), .I2(x1475), .I3(n6687), .I4(n6688), .O(n6691));
  LUT5 #(.INIT(32'hFF969600)) lut_n6692 (.I0(x1479), .I1(x1480), .I2(x1481), .I3(n6690), .I4(n6691), .O(n6692));
  LUT3 #(.INIT(8'h96)) lut_n6693 (.I0(n6681), .I1(n6684), .I2(n6685), .O(n6693));
  LUT3 #(.INIT(8'hE8)) lut_n6694 (.I0(n6689), .I1(n6692), .I2(n6693), .O(n6694));
  LUT3 #(.INIT(8'h96)) lut_n6695 (.I0(n6668), .I1(n6676), .I2(n6677), .O(n6695));
  LUT3 #(.INIT(8'hE8)) lut_n6696 (.I0(n6686), .I1(n6694), .I2(n6695), .O(n6696));
  LUT3 #(.INIT(8'h96)) lut_n6697 (.I0(n6640), .I1(n6658), .I2(n6659), .O(n6697));
  LUT3 #(.INIT(8'hE8)) lut_n6698 (.I0(n6678), .I1(n6696), .I2(n6697), .O(n6698));
  LUT3 #(.INIT(8'h96)) lut_n6699 (.I0(n6582), .I1(n6620), .I2(n6621), .O(n6699));
  LUT3 #(.INIT(8'hE8)) lut_n6700 (.I0(n6660), .I1(n6698), .I2(n6699), .O(n6700));
  LUT3 #(.INIT(8'h96)) lut_n6701 (.I0(n6462), .I1(n6540), .I2(n6541), .O(n6701));
  LUT3 #(.INIT(8'hE8)) lut_n6702 (.I0(n6622), .I1(n6700), .I2(n6701), .O(n6702));
  LUT3 #(.INIT(8'h96)) lut_n6703 (.I0(x1488), .I1(x1489), .I2(x1490), .O(n6703));
  LUT5 #(.INIT(32'h96696996)) lut_n6704 (.I0(x1479), .I1(x1480), .I2(x1481), .I3(n6690), .I4(n6691), .O(n6704));
  LUT5 #(.INIT(32'hFF969600)) lut_n6705 (.I0(x1485), .I1(x1486), .I2(x1487), .I3(n6703), .I4(n6704), .O(n6705));
  LUT3 #(.INIT(8'h96)) lut_n6706 (.I0(x1494), .I1(x1495), .I2(x1496), .O(n6706));
  LUT5 #(.INIT(32'h96696996)) lut_n6707 (.I0(x1485), .I1(x1486), .I2(x1487), .I3(n6703), .I4(n6704), .O(n6707));
  LUT5 #(.INIT(32'hFF969600)) lut_n6708 (.I0(x1491), .I1(x1492), .I2(x1493), .I3(n6706), .I4(n6707), .O(n6708));
  LUT3 #(.INIT(8'h96)) lut_n6709 (.I0(n6689), .I1(n6692), .I2(n6693), .O(n6709));
  LUT3 #(.INIT(8'hE8)) lut_n6710 (.I0(n6705), .I1(n6708), .I2(n6709), .O(n6710));
  LUT3 #(.INIT(8'h96)) lut_n6711 (.I0(x1500), .I1(x1501), .I2(x1502), .O(n6711));
  LUT5 #(.INIT(32'h96696996)) lut_n6712 (.I0(x1491), .I1(x1492), .I2(x1493), .I3(n6706), .I4(n6707), .O(n6712));
  LUT5 #(.INIT(32'hFF969600)) lut_n6713 (.I0(x1497), .I1(x1498), .I2(x1499), .I3(n6711), .I4(n6712), .O(n6713));
  LUT3 #(.INIT(8'h96)) lut_n6714 (.I0(x1506), .I1(x1507), .I2(x1508), .O(n6714));
  LUT5 #(.INIT(32'h96696996)) lut_n6715 (.I0(x1497), .I1(x1498), .I2(x1499), .I3(n6711), .I4(n6712), .O(n6715));
  LUT5 #(.INIT(32'hFF969600)) lut_n6716 (.I0(x1503), .I1(x1504), .I2(x1505), .I3(n6714), .I4(n6715), .O(n6716));
  LUT3 #(.INIT(8'h96)) lut_n6717 (.I0(n6705), .I1(n6708), .I2(n6709), .O(n6717));
  LUT3 #(.INIT(8'hE8)) lut_n6718 (.I0(n6713), .I1(n6716), .I2(n6717), .O(n6718));
  LUT3 #(.INIT(8'h96)) lut_n6719 (.I0(n6686), .I1(n6694), .I2(n6695), .O(n6719));
  LUT3 #(.INIT(8'hE8)) lut_n6720 (.I0(n6710), .I1(n6718), .I2(n6719), .O(n6720));
  LUT3 #(.INIT(8'h96)) lut_n6721 (.I0(x1512), .I1(x1513), .I2(x1514), .O(n6721));
  LUT5 #(.INIT(32'h96696996)) lut_n6722 (.I0(x1503), .I1(x1504), .I2(x1505), .I3(n6714), .I4(n6715), .O(n6722));
  LUT5 #(.INIT(32'hFF969600)) lut_n6723 (.I0(x1509), .I1(x1510), .I2(x1511), .I3(n6721), .I4(n6722), .O(n6723));
  LUT3 #(.INIT(8'h96)) lut_n6724 (.I0(x1518), .I1(x1519), .I2(x1520), .O(n6724));
  LUT5 #(.INIT(32'h96696996)) lut_n6725 (.I0(x1509), .I1(x1510), .I2(x1511), .I3(n6721), .I4(n6722), .O(n6725));
  LUT5 #(.INIT(32'hFF969600)) lut_n6726 (.I0(x1515), .I1(x1516), .I2(x1517), .I3(n6724), .I4(n6725), .O(n6726));
  LUT3 #(.INIT(8'h96)) lut_n6727 (.I0(n6713), .I1(n6716), .I2(n6717), .O(n6727));
  LUT3 #(.INIT(8'hE8)) lut_n6728 (.I0(n6723), .I1(n6726), .I2(n6727), .O(n6728));
  LUT3 #(.INIT(8'h96)) lut_n6729 (.I0(x1524), .I1(x1525), .I2(x1526), .O(n6729));
  LUT5 #(.INIT(32'h96696996)) lut_n6730 (.I0(x1515), .I1(x1516), .I2(x1517), .I3(n6724), .I4(n6725), .O(n6730));
  LUT5 #(.INIT(32'hFF969600)) lut_n6731 (.I0(x1521), .I1(x1522), .I2(x1523), .I3(n6729), .I4(n6730), .O(n6731));
  LUT3 #(.INIT(8'h96)) lut_n6732 (.I0(x1530), .I1(x1531), .I2(x1532), .O(n6732));
  LUT5 #(.INIT(32'h96696996)) lut_n6733 (.I0(x1521), .I1(x1522), .I2(x1523), .I3(n6729), .I4(n6730), .O(n6733));
  LUT5 #(.INIT(32'hFF969600)) lut_n6734 (.I0(x1527), .I1(x1528), .I2(x1529), .I3(n6732), .I4(n6733), .O(n6734));
  LUT3 #(.INIT(8'h96)) lut_n6735 (.I0(n6723), .I1(n6726), .I2(n6727), .O(n6735));
  LUT3 #(.INIT(8'hE8)) lut_n6736 (.I0(n6731), .I1(n6734), .I2(n6735), .O(n6736));
  LUT3 #(.INIT(8'h96)) lut_n6737 (.I0(n6710), .I1(n6718), .I2(n6719), .O(n6737));
  LUT3 #(.INIT(8'hE8)) lut_n6738 (.I0(n6728), .I1(n6736), .I2(n6737), .O(n6738));
  LUT3 #(.INIT(8'h96)) lut_n6739 (.I0(n6678), .I1(n6696), .I2(n6697), .O(n6739));
  LUT3 #(.INIT(8'hE8)) lut_n6740 (.I0(n6720), .I1(n6738), .I2(n6739), .O(n6740));
  LUT3 #(.INIT(8'h96)) lut_n6741 (.I0(x1536), .I1(x1537), .I2(x1538), .O(n6741));
  LUT5 #(.INIT(32'h96696996)) lut_n6742 (.I0(x1527), .I1(x1528), .I2(x1529), .I3(n6732), .I4(n6733), .O(n6742));
  LUT5 #(.INIT(32'hFF969600)) lut_n6743 (.I0(x1533), .I1(x1534), .I2(x1535), .I3(n6741), .I4(n6742), .O(n6743));
  LUT3 #(.INIT(8'h96)) lut_n6744 (.I0(x1542), .I1(x1543), .I2(x1544), .O(n6744));
  LUT5 #(.INIT(32'h96696996)) lut_n6745 (.I0(x1533), .I1(x1534), .I2(x1535), .I3(n6741), .I4(n6742), .O(n6745));
  LUT5 #(.INIT(32'hFF969600)) lut_n6746 (.I0(x1539), .I1(x1540), .I2(x1541), .I3(n6744), .I4(n6745), .O(n6746));
  LUT3 #(.INIT(8'h96)) lut_n6747 (.I0(n6731), .I1(n6734), .I2(n6735), .O(n6747));
  LUT3 #(.INIT(8'hE8)) lut_n6748 (.I0(n6743), .I1(n6746), .I2(n6747), .O(n6748));
  LUT3 #(.INIT(8'h96)) lut_n6749 (.I0(x1548), .I1(x1549), .I2(x1550), .O(n6749));
  LUT5 #(.INIT(32'h96696996)) lut_n6750 (.I0(x1539), .I1(x1540), .I2(x1541), .I3(n6744), .I4(n6745), .O(n6750));
  LUT5 #(.INIT(32'hFF969600)) lut_n6751 (.I0(x1545), .I1(x1546), .I2(x1547), .I3(n6749), .I4(n6750), .O(n6751));
  LUT3 #(.INIT(8'h96)) lut_n6752 (.I0(x1554), .I1(x1555), .I2(x1556), .O(n6752));
  LUT5 #(.INIT(32'h96696996)) lut_n6753 (.I0(x1545), .I1(x1546), .I2(x1547), .I3(n6749), .I4(n6750), .O(n6753));
  LUT5 #(.INIT(32'hFF969600)) lut_n6754 (.I0(x1551), .I1(x1552), .I2(x1553), .I3(n6752), .I4(n6753), .O(n6754));
  LUT3 #(.INIT(8'h96)) lut_n6755 (.I0(n6743), .I1(n6746), .I2(n6747), .O(n6755));
  LUT3 #(.INIT(8'hE8)) lut_n6756 (.I0(n6751), .I1(n6754), .I2(n6755), .O(n6756));
  LUT3 #(.INIT(8'h96)) lut_n6757 (.I0(n6728), .I1(n6736), .I2(n6737), .O(n6757));
  LUT3 #(.INIT(8'hE8)) lut_n6758 (.I0(n6748), .I1(n6756), .I2(n6757), .O(n6758));
  LUT3 #(.INIT(8'h96)) lut_n6759 (.I0(x1560), .I1(x1561), .I2(x1562), .O(n6759));
  LUT5 #(.INIT(32'h96696996)) lut_n6760 (.I0(x1551), .I1(x1552), .I2(x1553), .I3(n6752), .I4(n6753), .O(n6760));
  LUT5 #(.INIT(32'hFF969600)) lut_n6761 (.I0(x1557), .I1(x1558), .I2(x1559), .I3(n6759), .I4(n6760), .O(n6761));
  LUT3 #(.INIT(8'h96)) lut_n6762 (.I0(x1566), .I1(x1567), .I2(x1568), .O(n6762));
  LUT5 #(.INIT(32'h96696996)) lut_n6763 (.I0(x1557), .I1(x1558), .I2(x1559), .I3(n6759), .I4(n6760), .O(n6763));
  LUT5 #(.INIT(32'hFF969600)) lut_n6764 (.I0(x1563), .I1(x1564), .I2(x1565), .I3(n6762), .I4(n6763), .O(n6764));
  LUT3 #(.INIT(8'h96)) lut_n6765 (.I0(n6751), .I1(n6754), .I2(n6755), .O(n6765));
  LUT3 #(.INIT(8'hE8)) lut_n6766 (.I0(n6761), .I1(n6764), .I2(n6765), .O(n6766));
  LUT3 #(.INIT(8'h96)) lut_n6767 (.I0(x1572), .I1(x1573), .I2(x1574), .O(n6767));
  LUT5 #(.INIT(32'h96696996)) lut_n6768 (.I0(x1563), .I1(x1564), .I2(x1565), .I3(n6762), .I4(n6763), .O(n6768));
  LUT5 #(.INIT(32'hFF969600)) lut_n6769 (.I0(x1569), .I1(x1570), .I2(x1571), .I3(n6767), .I4(n6768), .O(n6769));
  LUT3 #(.INIT(8'h96)) lut_n6770 (.I0(x1578), .I1(x1579), .I2(x1580), .O(n6770));
  LUT5 #(.INIT(32'h96696996)) lut_n6771 (.I0(x1569), .I1(x1570), .I2(x1571), .I3(n6767), .I4(n6768), .O(n6771));
  LUT5 #(.INIT(32'hFF969600)) lut_n6772 (.I0(x1575), .I1(x1576), .I2(x1577), .I3(n6770), .I4(n6771), .O(n6772));
  LUT3 #(.INIT(8'h96)) lut_n6773 (.I0(n6761), .I1(n6764), .I2(n6765), .O(n6773));
  LUT3 #(.INIT(8'hE8)) lut_n6774 (.I0(n6769), .I1(n6772), .I2(n6773), .O(n6774));
  LUT3 #(.INIT(8'h96)) lut_n6775 (.I0(n6748), .I1(n6756), .I2(n6757), .O(n6775));
  LUT3 #(.INIT(8'hE8)) lut_n6776 (.I0(n6766), .I1(n6774), .I2(n6775), .O(n6776));
  LUT3 #(.INIT(8'h96)) lut_n6777 (.I0(n6720), .I1(n6738), .I2(n6739), .O(n6777));
  LUT3 #(.INIT(8'hE8)) lut_n6778 (.I0(n6758), .I1(n6776), .I2(n6777), .O(n6778));
  LUT3 #(.INIT(8'h96)) lut_n6779 (.I0(n6660), .I1(n6698), .I2(n6699), .O(n6779));
  LUT3 #(.INIT(8'hE8)) lut_n6780 (.I0(n6740), .I1(n6778), .I2(n6779), .O(n6780));
  LUT3 #(.INIT(8'h96)) lut_n6781 (.I0(x1584), .I1(x1585), .I2(x1586), .O(n6781));
  LUT5 #(.INIT(32'h96696996)) lut_n6782 (.I0(x1575), .I1(x1576), .I2(x1577), .I3(n6770), .I4(n6771), .O(n6782));
  LUT5 #(.INIT(32'hFF969600)) lut_n6783 (.I0(x1581), .I1(x1582), .I2(x1583), .I3(n6781), .I4(n6782), .O(n6783));
  LUT3 #(.INIT(8'h96)) lut_n6784 (.I0(x1590), .I1(x1591), .I2(x1592), .O(n6784));
  LUT5 #(.INIT(32'h96696996)) lut_n6785 (.I0(x1581), .I1(x1582), .I2(x1583), .I3(n6781), .I4(n6782), .O(n6785));
  LUT5 #(.INIT(32'hFF969600)) lut_n6786 (.I0(x1587), .I1(x1588), .I2(x1589), .I3(n6784), .I4(n6785), .O(n6786));
  LUT3 #(.INIT(8'h96)) lut_n6787 (.I0(n6769), .I1(n6772), .I2(n6773), .O(n6787));
  LUT3 #(.INIT(8'hE8)) lut_n6788 (.I0(n6783), .I1(n6786), .I2(n6787), .O(n6788));
  LUT3 #(.INIT(8'h96)) lut_n6789 (.I0(x1596), .I1(x1597), .I2(x1598), .O(n6789));
  LUT5 #(.INIT(32'h96696996)) lut_n6790 (.I0(x1587), .I1(x1588), .I2(x1589), .I3(n6784), .I4(n6785), .O(n6790));
  LUT5 #(.INIT(32'hFF969600)) lut_n6791 (.I0(x1593), .I1(x1594), .I2(x1595), .I3(n6789), .I4(n6790), .O(n6791));
  LUT3 #(.INIT(8'h96)) lut_n6792 (.I0(x1602), .I1(x1603), .I2(x1604), .O(n6792));
  LUT5 #(.INIT(32'h96696996)) lut_n6793 (.I0(x1593), .I1(x1594), .I2(x1595), .I3(n6789), .I4(n6790), .O(n6793));
  LUT5 #(.INIT(32'hFF969600)) lut_n6794 (.I0(x1599), .I1(x1600), .I2(x1601), .I3(n6792), .I4(n6793), .O(n6794));
  LUT3 #(.INIT(8'h96)) lut_n6795 (.I0(n6783), .I1(n6786), .I2(n6787), .O(n6795));
  LUT3 #(.INIT(8'hE8)) lut_n6796 (.I0(n6791), .I1(n6794), .I2(n6795), .O(n6796));
  LUT3 #(.INIT(8'h96)) lut_n6797 (.I0(n6766), .I1(n6774), .I2(n6775), .O(n6797));
  LUT3 #(.INIT(8'hE8)) lut_n6798 (.I0(n6788), .I1(n6796), .I2(n6797), .O(n6798));
  LUT3 #(.INIT(8'h96)) lut_n6799 (.I0(x1608), .I1(x1609), .I2(x1610), .O(n6799));
  LUT5 #(.INIT(32'h96696996)) lut_n6800 (.I0(x1599), .I1(x1600), .I2(x1601), .I3(n6792), .I4(n6793), .O(n6800));
  LUT5 #(.INIT(32'hFF969600)) lut_n6801 (.I0(x1605), .I1(x1606), .I2(x1607), .I3(n6799), .I4(n6800), .O(n6801));
  LUT3 #(.INIT(8'h96)) lut_n6802 (.I0(x1614), .I1(x1615), .I2(x1616), .O(n6802));
  LUT5 #(.INIT(32'h96696996)) lut_n6803 (.I0(x1605), .I1(x1606), .I2(x1607), .I3(n6799), .I4(n6800), .O(n6803));
  LUT5 #(.INIT(32'hFF969600)) lut_n6804 (.I0(x1611), .I1(x1612), .I2(x1613), .I3(n6802), .I4(n6803), .O(n6804));
  LUT3 #(.INIT(8'h96)) lut_n6805 (.I0(n6791), .I1(n6794), .I2(n6795), .O(n6805));
  LUT3 #(.INIT(8'hE8)) lut_n6806 (.I0(n6801), .I1(n6804), .I2(n6805), .O(n6806));
  LUT3 #(.INIT(8'h96)) lut_n6807 (.I0(x1620), .I1(x1621), .I2(x1622), .O(n6807));
  LUT5 #(.INIT(32'h96696996)) lut_n6808 (.I0(x1611), .I1(x1612), .I2(x1613), .I3(n6802), .I4(n6803), .O(n6808));
  LUT5 #(.INIT(32'hFF969600)) lut_n6809 (.I0(x1617), .I1(x1618), .I2(x1619), .I3(n6807), .I4(n6808), .O(n6809));
  LUT3 #(.INIT(8'h96)) lut_n6810 (.I0(x1626), .I1(x1627), .I2(x1628), .O(n6810));
  LUT5 #(.INIT(32'h96696996)) lut_n6811 (.I0(x1617), .I1(x1618), .I2(x1619), .I3(n6807), .I4(n6808), .O(n6811));
  LUT5 #(.INIT(32'hFF969600)) lut_n6812 (.I0(x1623), .I1(x1624), .I2(x1625), .I3(n6810), .I4(n6811), .O(n6812));
  LUT3 #(.INIT(8'h96)) lut_n6813 (.I0(n6801), .I1(n6804), .I2(n6805), .O(n6813));
  LUT3 #(.INIT(8'hE8)) lut_n6814 (.I0(n6809), .I1(n6812), .I2(n6813), .O(n6814));
  LUT3 #(.INIT(8'h96)) lut_n6815 (.I0(n6788), .I1(n6796), .I2(n6797), .O(n6815));
  LUT3 #(.INIT(8'hE8)) lut_n6816 (.I0(n6806), .I1(n6814), .I2(n6815), .O(n6816));
  LUT3 #(.INIT(8'h96)) lut_n6817 (.I0(n6758), .I1(n6776), .I2(n6777), .O(n6817));
  LUT3 #(.INIT(8'hE8)) lut_n6818 (.I0(n6798), .I1(n6816), .I2(n6817), .O(n6818));
  LUT3 #(.INIT(8'h96)) lut_n6819 (.I0(x1632), .I1(x1633), .I2(x1634), .O(n6819));
  LUT5 #(.INIT(32'h96696996)) lut_n6820 (.I0(x1623), .I1(x1624), .I2(x1625), .I3(n6810), .I4(n6811), .O(n6820));
  LUT5 #(.INIT(32'hFF969600)) lut_n6821 (.I0(x1629), .I1(x1630), .I2(x1631), .I3(n6819), .I4(n6820), .O(n6821));
  LUT3 #(.INIT(8'h96)) lut_n6822 (.I0(x1638), .I1(x1639), .I2(x1640), .O(n6822));
  LUT5 #(.INIT(32'h96696996)) lut_n6823 (.I0(x1629), .I1(x1630), .I2(x1631), .I3(n6819), .I4(n6820), .O(n6823));
  LUT5 #(.INIT(32'hFF969600)) lut_n6824 (.I0(x1635), .I1(x1636), .I2(x1637), .I3(n6822), .I4(n6823), .O(n6824));
  LUT3 #(.INIT(8'h96)) lut_n6825 (.I0(n6809), .I1(n6812), .I2(n6813), .O(n6825));
  LUT3 #(.INIT(8'hE8)) lut_n6826 (.I0(n6821), .I1(n6824), .I2(n6825), .O(n6826));
  LUT3 #(.INIT(8'h96)) lut_n6827 (.I0(x1644), .I1(x1645), .I2(x1646), .O(n6827));
  LUT5 #(.INIT(32'h96696996)) lut_n6828 (.I0(x1635), .I1(x1636), .I2(x1637), .I3(n6822), .I4(n6823), .O(n6828));
  LUT5 #(.INIT(32'hFF969600)) lut_n6829 (.I0(x1641), .I1(x1642), .I2(x1643), .I3(n6827), .I4(n6828), .O(n6829));
  LUT3 #(.INIT(8'h96)) lut_n6830 (.I0(x1650), .I1(x1651), .I2(x1652), .O(n6830));
  LUT5 #(.INIT(32'h96696996)) lut_n6831 (.I0(x1641), .I1(x1642), .I2(x1643), .I3(n6827), .I4(n6828), .O(n6831));
  LUT5 #(.INIT(32'hFF969600)) lut_n6832 (.I0(x1647), .I1(x1648), .I2(x1649), .I3(n6830), .I4(n6831), .O(n6832));
  LUT3 #(.INIT(8'h96)) lut_n6833 (.I0(n6821), .I1(n6824), .I2(n6825), .O(n6833));
  LUT3 #(.INIT(8'hE8)) lut_n6834 (.I0(n6829), .I1(n6832), .I2(n6833), .O(n6834));
  LUT3 #(.INIT(8'h96)) lut_n6835 (.I0(n6806), .I1(n6814), .I2(n6815), .O(n6835));
  LUT3 #(.INIT(8'hE8)) lut_n6836 (.I0(n6826), .I1(n6834), .I2(n6835), .O(n6836));
  LUT3 #(.INIT(8'h96)) lut_n6837 (.I0(x1656), .I1(x1657), .I2(x1658), .O(n6837));
  LUT5 #(.INIT(32'h96696996)) lut_n6838 (.I0(x1647), .I1(x1648), .I2(x1649), .I3(n6830), .I4(n6831), .O(n6838));
  LUT5 #(.INIT(32'hFF969600)) lut_n6839 (.I0(x1653), .I1(x1654), .I2(x1655), .I3(n6837), .I4(n6838), .O(n6839));
  LUT3 #(.INIT(8'h96)) lut_n6840 (.I0(x1662), .I1(x1663), .I2(x1664), .O(n6840));
  LUT5 #(.INIT(32'h96696996)) lut_n6841 (.I0(x1653), .I1(x1654), .I2(x1655), .I3(n6837), .I4(n6838), .O(n6841));
  LUT5 #(.INIT(32'hFF969600)) lut_n6842 (.I0(x1659), .I1(x1660), .I2(x1661), .I3(n6840), .I4(n6841), .O(n6842));
  LUT3 #(.INIT(8'h96)) lut_n6843 (.I0(n6829), .I1(n6832), .I2(n6833), .O(n6843));
  LUT3 #(.INIT(8'hE8)) lut_n6844 (.I0(n6839), .I1(n6842), .I2(n6843), .O(n6844));
  LUT3 #(.INIT(8'h96)) lut_n6845 (.I0(x1668), .I1(x1669), .I2(x1670), .O(n6845));
  LUT5 #(.INIT(32'h96696996)) lut_n6846 (.I0(x1659), .I1(x1660), .I2(x1661), .I3(n6840), .I4(n6841), .O(n6846));
  LUT5 #(.INIT(32'hFF969600)) lut_n6847 (.I0(x1665), .I1(x1666), .I2(x1667), .I3(n6845), .I4(n6846), .O(n6847));
  LUT3 #(.INIT(8'h96)) lut_n6848 (.I0(x1674), .I1(x1675), .I2(x1676), .O(n6848));
  LUT5 #(.INIT(32'h96696996)) lut_n6849 (.I0(x1665), .I1(x1666), .I2(x1667), .I3(n6845), .I4(n6846), .O(n6849));
  LUT5 #(.INIT(32'hFF969600)) lut_n6850 (.I0(x1671), .I1(x1672), .I2(x1673), .I3(n6848), .I4(n6849), .O(n6850));
  LUT3 #(.INIT(8'h96)) lut_n6851 (.I0(n6839), .I1(n6842), .I2(n6843), .O(n6851));
  LUT3 #(.INIT(8'hE8)) lut_n6852 (.I0(n6847), .I1(n6850), .I2(n6851), .O(n6852));
  LUT3 #(.INIT(8'h96)) lut_n6853 (.I0(n6826), .I1(n6834), .I2(n6835), .O(n6853));
  LUT3 #(.INIT(8'hE8)) lut_n6854 (.I0(n6844), .I1(n6852), .I2(n6853), .O(n6854));
  LUT3 #(.INIT(8'h96)) lut_n6855 (.I0(n6798), .I1(n6816), .I2(n6817), .O(n6855));
  LUT3 #(.INIT(8'hE8)) lut_n6856 (.I0(n6836), .I1(n6854), .I2(n6855), .O(n6856));
  LUT3 #(.INIT(8'h96)) lut_n6857 (.I0(n6740), .I1(n6778), .I2(n6779), .O(n6857));
  LUT3 #(.INIT(8'hE8)) lut_n6858 (.I0(n6818), .I1(n6856), .I2(n6857), .O(n6858));
  LUT3 #(.INIT(8'h96)) lut_n6859 (.I0(n6622), .I1(n6700), .I2(n6701), .O(n6859));
  LUT3 #(.INIT(8'hE8)) lut_n6860 (.I0(n6780), .I1(n6858), .I2(n6859), .O(n6860));
  LUT3 #(.INIT(8'h96)) lut_n6861 (.I0(n6384), .I1(n6542), .I2(n6543), .O(n6861));
  LUT3 #(.INIT(8'hE8)) lut_n6862 (.I0(n6702), .I1(n6860), .I2(n6861), .O(n6862));
  LUT3 #(.INIT(8'h96)) lut_n6863 (.I0(n5906), .I1(n6224), .I2(n6225), .O(n6863));
  LUT3 #(.INIT(8'hE8)) lut_n6864 (.I0(n6544), .I1(n6862), .I2(n6863), .O(n6864));
  LUT3 #(.INIT(8'h96)) lut_n6865 (.I0(n5210), .I1(n5585), .I2(n5586), .O(n6865));
  LUT3 #(.INIT(8'hE8)) lut_n6866 (.I0(n6226), .I1(n6864), .I2(n6865), .O(n6866));
  LUT3 #(.INIT(8'h96)) lut_n6867 (.I0(x1680), .I1(x1681), .I2(x1682), .O(n6867));
  LUT5 #(.INIT(32'h96696996)) lut_n6868 (.I0(x1671), .I1(x1672), .I2(x1673), .I3(n6848), .I4(n6849), .O(n6868));
  LUT5 #(.INIT(32'hFF969600)) lut_n6869 (.I0(x1677), .I1(x1678), .I2(x1679), .I3(n6867), .I4(n6868), .O(n6869));
  LUT3 #(.INIT(8'h96)) lut_n6870 (.I0(x1686), .I1(x1687), .I2(x1688), .O(n6870));
  LUT5 #(.INIT(32'h96696996)) lut_n6871 (.I0(x1677), .I1(x1678), .I2(x1679), .I3(n6867), .I4(n6868), .O(n6871));
  LUT5 #(.INIT(32'hFF969600)) lut_n6872 (.I0(x1683), .I1(x1684), .I2(x1685), .I3(n6870), .I4(n6871), .O(n6872));
  LUT3 #(.INIT(8'h96)) lut_n6873 (.I0(n6847), .I1(n6850), .I2(n6851), .O(n6873));
  LUT3 #(.INIT(8'hE8)) lut_n6874 (.I0(n6869), .I1(n6872), .I2(n6873), .O(n6874));
  LUT3 #(.INIT(8'h96)) lut_n6875 (.I0(x1692), .I1(x1693), .I2(x1694), .O(n6875));
  LUT5 #(.INIT(32'h96696996)) lut_n6876 (.I0(x1683), .I1(x1684), .I2(x1685), .I3(n6870), .I4(n6871), .O(n6876));
  LUT5 #(.INIT(32'hFF969600)) lut_n6877 (.I0(x1689), .I1(x1690), .I2(x1691), .I3(n6875), .I4(n6876), .O(n6877));
  LUT3 #(.INIT(8'h96)) lut_n6878 (.I0(x1698), .I1(x1699), .I2(x1700), .O(n6878));
  LUT5 #(.INIT(32'h96696996)) lut_n6879 (.I0(x1689), .I1(x1690), .I2(x1691), .I3(n6875), .I4(n6876), .O(n6879));
  LUT5 #(.INIT(32'hFF969600)) lut_n6880 (.I0(x1695), .I1(x1696), .I2(x1697), .I3(n6878), .I4(n6879), .O(n6880));
  LUT3 #(.INIT(8'h96)) lut_n6881 (.I0(n6869), .I1(n6872), .I2(n6873), .O(n6881));
  LUT3 #(.INIT(8'hE8)) lut_n6882 (.I0(n6877), .I1(n6880), .I2(n6881), .O(n6882));
  LUT3 #(.INIT(8'h96)) lut_n6883 (.I0(n6844), .I1(n6852), .I2(n6853), .O(n6883));
  LUT3 #(.INIT(8'hE8)) lut_n6884 (.I0(n6874), .I1(n6882), .I2(n6883), .O(n6884));
  LUT3 #(.INIT(8'h96)) lut_n6885 (.I0(x1704), .I1(x1705), .I2(x1706), .O(n6885));
  LUT5 #(.INIT(32'h96696996)) lut_n6886 (.I0(x1695), .I1(x1696), .I2(x1697), .I3(n6878), .I4(n6879), .O(n6886));
  LUT5 #(.INIT(32'hFF969600)) lut_n6887 (.I0(x1701), .I1(x1702), .I2(x1703), .I3(n6885), .I4(n6886), .O(n6887));
  LUT3 #(.INIT(8'h96)) lut_n6888 (.I0(x1710), .I1(x1711), .I2(x1712), .O(n6888));
  LUT5 #(.INIT(32'h96696996)) lut_n6889 (.I0(x1701), .I1(x1702), .I2(x1703), .I3(n6885), .I4(n6886), .O(n6889));
  LUT5 #(.INIT(32'hFF969600)) lut_n6890 (.I0(x1707), .I1(x1708), .I2(x1709), .I3(n6888), .I4(n6889), .O(n6890));
  LUT3 #(.INIT(8'h96)) lut_n6891 (.I0(n6877), .I1(n6880), .I2(n6881), .O(n6891));
  LUT3 #(.INIT(8'hE8)) lut_n6892 (.I0(n6887), .I1(n6890), .I2(n6891), .O(n6892));
  LUT3 #(.INIT(8'h96)) lut_n6893 (.I0(x1716), .I1(x1717), .I2(x1718), .O(n6893));
  LUT5 #(.INIT(32'h96696996)) lut_n6894 (.I0(x1707), .I1(x1708), .I2(x1709), .I3(n6888), .I4(n6889), .O(n6894));
  LUT5 #(.INIT(32'hFF969600)) lut_n6895 (.I0(x1713), .I1(x1714), .I2(x1715), .I3(n6893), .I4(n6894), .O(n6895));
  LUT3 #(.INIT(8'h96)) lut_n6896 (.I0(x1722), .I1(x1723), .I2(x1724), .O(n6896));
  LUT5 #(.INIT(32'h96696996)) lut_n6897 (.I0(x1713), .I1(x1714), .I2(x1715), .I3(n6893), .I4(n6894), .O(n6897));
  LUT5 #(.INIT(32'hFF969600)) lut_n6898 (.I0(x1719), .I1(x1720), .I2(x1721), .I3(n6896), .I4(n6897), .O(n6898));
  LUT3 #(.INIT(8'h96)) lut_n6899 (.I0(n6887), .I1(n6890), .I2(n6891), .O(n6899));
  LUT3 #(.INIT(8'hE8)) lut_n6900 (.I0(n6895), .I1(n6898), .I2(n6899), .O(n6900));
  LUT3 #(.INIT(8'h96)) lut_n6901 (.I0(n6874), .I1(n6882), .I2(n6883), .O(n6901));
  LUT3 #(.INIT(8'hE8)) lut_n6902 (.I0(n6892), .I1(n6900), .I2(n6901), .O(n6902));
  LUT3 #(.INIT(8'h96)) lut_n6903 (.I0(n6836), .I1(n6854), .I2(n6855), .O(n6903));
  LUT3 #(.INIT(8'hE8)) lut_n6904 (.I0(n6884), .I1(n6902), .I2(n6903), .O(n6904));
  LUT3 #(.INIT(8'h96)) lut_n6905 (.I0(x1728), .I1(x1729), .I2(x1730), .O(n6905));
  LUT5 #(.INIT(32'h96696996)) lut_n6906 (.I0(x1719), .I1(x1720), .I2(x1721), .I3(n6896), .I4(n6897), .O(n6906));
  LUT5 #(.INIT(32'hFF969600)) lut_n6907 (.I0(x1725), .I1(x1726), .I2(x1727), .I3(n6905), .I4(n6906), .O(n6907));
  LUT3 #(.INIT(8'h96)) lut_n6908 (.I0(x1734), .I1(x1735), .I2(x1736), .O(n6908));
  LUT5 #(.INIT(32'h96696996)) lut_n6909 (.I0(x1725), .I1(x1726), .I2(x1727), .I3(n6905), .I4(n6906), .O(n6909));
  LUT5 #(.INIT(32'hFF969600)) lut_n6910 (.I0(x1731), .I1(x1732), .I2(x1733), .I3(n6908), .I4(n6909), .O(n6910));
  LUT3 #(.INIT(8'h96)) lut_n6911 (.I0(n6895), .I1(n6898), .I2(n6899), .O(n6911));
  LUT3 #(.INIT(8'hE8)) lut_n6912 (.I0(n6907), .I1(n6910), .I2(n6911), .O(n6912));
  LUT3 #(.INIT(8'h96)) lut_n6913 (.I0(x1740), .I1(x1741), .I2(x1742), .O(n6913));
  LUT5 #(.INIT(32'h96696996)) lut_n6914 (.I0(x1731), .I1(x1732), .I2(x1733), .I3(n6908), .I4(n6909), .O(n6914));
  LUT5 #(.INIT(32'hFF969600)) lut_n6915 (.I0(x1737), .I1(x1738), .I2(x1739), .I3(n6913), .I4(n6914), .O(n6915));
  LUT3 #(.INIT(8'h96)) lut_n6916 (.I0(x1746), .I1(x1747), .I2(x1748), .O(n6916));
  LUT5 #(.INIT(32'h96696996)) lut_n6917 (.I0(x1737), .I1(x1738), .I2(x1739), .I3(n6913), .I4(n6914), .O(n6917));
  LUT5 #(.INIT(32'hFF969600)) lut_n6918 (.I0(x1743), .I1(x1744), .I2(x1745), .I3(n6916), .I4(n6917), .O(n6918));
  LUT3 #(.INIT(8'h96)) lut_n6919 (.I0(n6907), .I1(n6910), .I2(n6911), .O(n6919));
  LUT3 #(.INIT(8'hE8)) lut_n6920 (.I0(n6915), .I1(n6918), .I2(n6919), .O(n6920));
  LUT3 #(.INIT(8'h96)) lut_n6921 (.I0(n6892), .I1(n6900), .I2(n6901), .O(n6921));
  LUT3 #(.INIT(8'hE8)) lut_n6922 (.I0(n6912), .I1(n6920), .I2(n6921), .O(n6922));
  LUT3 #(.INIT(8'h96)) lut_n6923 (.I0(x1752), .I1(x1753), .I2(x1754), .O(n6923));
  LUT5 #(.INIT(32'h96696996)) lut_n6924 (.I0(x1743), .I1(x1744), .I2(x1745), .I3(n6916), .I4(n6917), .O(n6924));
  LUT5 #(.INIT(32'hFF969600)) lut_n6925 (.I0(x1749), .I1(x1750), .I2(x1751), .I3(n6923), .I4(n6924), .O(n6925));
  LUT3 #(.INIT(8'h96)) lut_n6926 (.I0(x1758), .I1(x1759), .I2(x1760), .O(n6926));
  LUT5 #(.INIT(32'h96696996)) lut_n6927 (.I0(x1749), .I1(x1750), .I2(x1751), .I3(n6923), .I4(n6924), .O(n6927));
  LUT5 #(.INIT(32'hFF969600)) lut_n6928 (.I0(x1755), .I1(x1756), .I2(x1757), .I3(n6926), .I4(n6927), .O(n6928));
  LUT3 #(.INIT(8'h96)) lut_n6929 (.I0(n6915), .I1(n6918), .I2(n6919), .O(n6929));
  LUT3 #(.INIT(8'hE8)) lut_n6930 (.I0(n6925), .I1(n6928), .I2(n6929), .O(n6930));
  LUT3 #(.INIT(8'h96)) lut_n6931 (.I0(x1764), .I1(x1765), .I2(x1766), .O(n6931));
  LUT5 #(.INIT(32'h96696996)) lut_n6932 (.I0(x1755), .I1(x1756), .I2(x1757), .I3(n6926), .I4(n6927), .O(n6932));
  LUT5 #(.INIT(32'hFF969600)) lut_n6933 (.I0(x1761), .I1(x1762), .I2(x1763), .I3(n6931), .I4(n6932), .O(n6933));
  LUT3 #(.INIT(8'h96)) lut_n6934 (.I0(x1770), .I1(x1771), .I2(x1772), .O(n6934));
  LUT5 #(.INIT(32'h96696996)) lut_n6935 (.I0(x1761), .I1(x1762), .I2(x1763), .I3(n6931), .I4(n6932), .O(n6935));
  LUT5 #(.INIT(32'hFF969600)) lut_n6936 (.I0(x1767), .I1(x1768), .I2(x1769), .I3(n6934), .I4(n6935), .O(n6936));
  LUT3 #(.INIT(8'h96)) lut_n6937 (.I0(n6925), .I1(n6928), .I2(n6929), .O(n6937));
  LUT3 #(.INIT(8'hE8)) lut_n6938 (.I0(n6933), .I1(n6936), .I2(n6937), .O(n6938));
  LUT3 #(.INIT(8'h96)) lut_n6939 (.I0(n6912), .I1(n6920), .I2(n6921), .O(n6939));
  LUT3 #(.INIT(8'hE8)) lut_n6940 (.I0(n6930), .I1(n6938), .I2(n6939), .O(n6940));
  LUT3 #(.INIT(8'h96)) lut_n6941 (.I0(n6884), .I1(n6902), .I2(n6903), .O(n6941));
  LUT3 #(.INIT(8'hE8)) lut_n6942 (.I0(n6922), .I1(n6940), .I2(n6941), .O(n6942));
  LUT3 #(.INIT(8'h96)) lut_n6943 (.I0(n6818), .I1(n6856), .I2(n6857), .O(n6943));
  LUT3 #(.INIT(8'hE8)) lut_n6944 (.I0(n6904), .I1(n6942), .I2(n6943), .O(n6944));
  LUT3 #(.INIT(8'h96)) lut_n6945 (.I0(x1776), .I1(x1777), .I2(x1778), .O(n6945));
  LUT5 #(.INIT(32'h96696996)) lut_n6946 (.I0(x1767), .I1(x1768), .I2(x1769), .I3(n6934), .I4(n6935), .O(n6946));
  LUT5 #(.INIT(32'hFF969600)) lut_n6947 (.I0(x1773), .I1(x1774), .I2(x1775), .I3(n6945), .I4(n6946), .O(n6947));
  LUT3 #(.INIT(8'h96)) lut_n6948 (.I0(x1782), .I1(x1783), .I2(x1784), .O(n6948));
  LUT5 #(.INIT(32'h96696996)) lut_n6949 (.I0(x1773), .I1(x1774), .I2(x1775), .I3(n6945), .I4(n6946), .O(n6949));
  LUT5 #(.INIT(32'hFF969600)) lut_n6950 (.I0(x1779), .I1(x1780), .I2(x1781), .I3(n6948), .I4(n6949), .O(n6950));
  LUT3 #(.INIT(8'h96)) lut_n6951 (.I0(n6933), .I1(n6936), .I2(n6937), .O(n6951));
  LUT3 #(.INIT(8'hE8)) lut_n6952 (.I0(n6947), .I1(n6950), .I2(n6951), .O(n6952));
  LUT3 #(.INIT(8'h96)) lut_n6953 (.I0(x1788), .I1(x1789), .I2(x1790), .O(n6953));
  LUT5 #(.INIT(32'h96696996)) lut_n6954 (.I0(x1779), .I1(x1780), .I2(x1781), .I3(n6948), .I4(n6949), .O(n6954));
  LUT5 #(.INIT(32'hFF969600)) lut_n6955 (.I0(x1785), .I1(x1786), .I2(x1787), .I3(n6953), .I4(n6954), .O(n6955));
  LUT3 #(.INIT(8'h96)) lut_n6956 (.I0(x1794), .I1(x1795), .I2(x1796), .O(n6956));
  LUT5 #(.INIT(32'h96696996)) lut_n6957 (.I0(x1785), .I1(x1786), .I2(x1787), .I3(n6953), .I4(n6954), .O(n6957));
  LUT5 #(.INIT(32'hFF969600)) lut_n6958 (.I0(x1791), .I1(x1792), .I2(x1793), .I3(n6956), .I4(n6957), .O(n6958));
  LUT3 #(.INIT(8'h96)) lut_n6959 (.I0(n6947), .I1(n6950), .I2(n6951), .O(n6959));
  LUT3 #(.INIT(8'hE8)) lut_n6960 (.I0(n6955), .I1(n6958), .I2(n6959), .O(n6960));
  LUT3 #(.INIT(8'h96)) lut_n6961 (.I0(n6930), .I1(n6938), .I2(n6939), .O(n6961));
  LUT3 #(.INIT(8'hE8)) lut_n6962 (.I0(n6952), .I1(n6960), .I2(n6961), .O(n6962));
  LUT3 #(.INIT(8'h96)) lut_n6963 (.I0(x1800), .I1(x1801), .I2(x1802), .O(n6963));
  LUT5 #(.INIT(32'h96696996)) lut_n6964 (.I0(x1791), .I1(x1792), .I2(x1793), .I3(n6956), .I4(n6957), .O(n6964));
  LUT5 #(.INIT(32'hFF969600)) lut_n6965 (.I0(x1797), .I1(x1798), .I2(x1799), .I3(n6963), .I4(n6964), .O(n6965));
  LUT3 #(.INIT(8'h96)) lut_n6966 (.I0(x1806), .I1(x1807), .I2(x1808), .O(n6966));
  LUT5 #(.INIT(32'h96696996)) lut_n6967 (.I0(x1797), .I1(x1798), .I2(x1799), .I3(n6963), .I4(n6964), .O(n6967));
  LUT5 #(.INIT(32'hFF969600)) lut_n6968 (.I0(x1803), .I1(x1804), .I2(x1805), .I3(n6966), .I4(n6967), .O(n6968));
  LUT3 #(.INIT(8'h96)) lut_n6969 (.I0(n6955), .I1(n6958), .I2(n6959), .O(n6969));
  LUT3 #(.INIT(8'hE8)) lut_n6970 (.I0(n6965), .I1(n6968), .I2(n6969), .O(n6970));
  LUT3 #(.INIT(8'h96)) lut_n6971 (.I0(x1812), .I1(x1813), .I2(x1814), .O(n6971));
  LUT5 #(.INIT(32'h96696996)) lut_n6972 (.I0(x1803), .I1(x1804), .I2(x1805), .I3(n6966), .I4(n6967), .O(n6972));
  LUT5 #(.INIT(32'hFF969600)) lut_n6973 (.I0(x1809), .I1(x1810), .I2(x1811), .I3(n6971), .I4(n6972), .O(n6973));
  LUT3 #(.INIT(8'h96)) lut_n6974 (.I0(x1818), .I1(x1819), .I2(x1820), .O(n6974));
  LUT5 #(.INIT(32'h96696996)) lut_n6975 (.I0(x1809), .I1(x1810), .I2(x1811), .I3(n6971), .I4(n6972), .O(n6975));
  LUT5 #(.INIT(32'hFF969600)) lut_n6976 (.I0(x1815), .I1(x1816), .I2(x1817), .I3(n6974), .I4(n6975), .O(n6976));
  LUT3 #(.INIT(8'h96)) lut_n6977 (.I0(n6965), .I1(n6968), .I2(n6969), .O(n6977));
  LUT3 #(.INIT(8'hE8)) lut_n6978 (.I0(n6973), .I1(n6976), .I2(n6977), .O(n6978));
  LUT3 #(.INIT(8'h96)) lut_n6979 (.I0(n6952), .I1(n6960), .I2(n6961), .O(n6979));
  LUT3 #(.INIT(8'hE8)) lut_n6980 (.I0(n6970), .I1(n6978), .I2(n6979), .O(n6980));
  LUT3 #(.INIT(8'h96)) lut_n6981 (.I0(n6922), .I1(n6940), .I2(n6941), .O(n6981));
  LUT3 #(.INIT(8'hE8)) lut_n6982 (.I0(n6962), .I1(n6980), .I2(n6981), .O(n6982));
  LUT3 #(.INIT(8'h96)) lut_n6983 (.I0(x1824), .I1(x1825), .I2(x1826), .O(n6983));
  LUT5 #(.INIT(32'h96696996)) lut_n6984 (.I0(x1815), .I1(x1816), .I2(x1817), .I3(n6974), .I4(n6975), .O(n6984));
  LUT5 #(.INIT(32'hFF969600)) lut_n6985 (.I0(x1821), .I1(x1822), .I2(x1823), .I3(n6983), .I4(n6984), .O(n6985));
  LUT3 #(.INIT(8'h96)) lut_n6986 (.I0(x1830), .I1(x1831), .I2(x1832), .O(n6986));
  LUT5 #(.INIT(32'h96696996)) lut_n6987 (.I0(x1821), .I1(x1822), .I2(x1823), .I3(n6983), .I4(n6984), .O(n6987));
  LUT5 #(.INIT(32'hFF969600)) lut_n6988 (.I0(x1827), .I1(x1828), .I2(x1829), .I3(n6986), .I4(n6987), .O(n6988));
  LUT3 #(.INIT(8'h96)) lut_n6989 (.I0(n6973), .I1(n6976), .I2(n6977), .O(n6989));
  LUT3 #(.INIT(8'hE8)) lut_n6990 (.I0(n6985), .I1(n6988), .I2(n6989), .O(n6990));
  LUT3 #(.INIT(8'h96)) lut_n6991 (.I0(x1836), .I1(x1837), .I2(x1838), .O(n6991));
  LUT5 #(.INIT(32'h96696996)) lut_n6992 (.I0(x1827), .I1(x1828), .I2(x1829), .I3(n6986), .I4(n6987), .O(n6992));
  LUT5 #(.INIT(32'hFF969600)) lut_n6993 (.I0(x1833), .I1(x1834), .I2(x1835), .I3(n6991), .I4(n6992), .O(n6993));
  LUT3 #(.INIT(8'h96)) lut_n6994 (.I0(x1842), .I1(x1843), .I2(x1844), .O(n6994));
  LUT5 #(.INIT(32'h96696996)) lut_n6995 (.I0(x1833), .I1(x1834), .I2(x1835), .I3(n6991), .I4(n6992), .O(n6995));
  LUT5 #(.INIT(32'hFF969600)) lut_n6996 (.I0(x1839), .I1(x1840), .I2(x1841), .I3(n6994), .I4(n6995), .O(n6996));
  LUT3 #(.INIT(8'h96)) lut_n6997 (.I0(n6985), .I1(n6988), .I2(n6989), .O(n6997));
  LUT3 #(.INIT(8'hE8)) lut_n6998 (.I0(n6993), .I1(n6996), .I2(n6997), .O(n6998));
  LUT3 #(.INIT(8'h96)) lut_n6999 (.I0(n6970), .I1(n6978), .I2(n6979), .O(n6999));
  LUT3 #(.INIT(8'hE8)) lut_n7000 (.I0(n6990), .I1(n6998), .I2(n6999), .O(n7000));
  LUT3 #(.INIT(8'h96)) lut_n7001 (.I0(x1848), .I1(x1849), .I2(x1850), .O(n7001));
  LUT5 #(.INIT(32'h96696996)) lut_n7002 (.I0(x1839), .I1(x1840), .I2(x1841), .I3(n6994), .I4(n6995), .O(n7002));
  LUT5 #(.INIT(32'hFF969600)) lut_n7003 (.I0(x1845), .I1(x1846), .I2(x1847), .I3(n7001), .I4(n7002), .O(n7003));
  LUT3 #(.INIT(8'h96)) lut_n7004 (.I0(x1854), .I1(x1855), .I2(x1856), .O(n7004));
  LUT5 #(.INIT(32'h96696996)) lut_n7005 (.I0(x1845), .I1(x1846), .I2(x1847), .I3(n7001), .I4(n7002), .O(n7005));
  LUT5 #(.INIT(32'hFF969600)) lut_n7006 (.I0(x1851), .I1(x1852), .I2(x1853), .I3(n7004), .I4(n7005), .O(n7006));
  LUT3 #(.INIT(8'h96)) lut_n7007 (.I0(n6993), .I1(n6996), .I2(n6997), .O(n7007));
  LUT3 #(.INIT(8'hE8)) lut_n7008 (.I0(n7003), .I1(n7006), .I2(n7007), .O(n7008));
  LUT3 #(.INIT(8'h96)) lut_n7009 (.I0(x1860), .I1(x1861), .I2(x1862), .O(n7009));
  LUT5 #(.INIT(32'h96696996)) lut_n7010 (.I0(x1851), .I1(x1852), .I2(x1853), .I3(n7004), .I4(n7005), .O(n7010));
  LUT5 #(.INIT(32'hFF969600)) lut_n7011 (.I0(x1857), .I1(x1858), .I2(x1859), .I3(n7009), .I4(n7010), .O(n7011));
  LUT3 #(.INIT(8'h96)) lut_n7012 (.I0(x1866), .I1(x1867), .I2(x1868), .O(n7012));
  LUT5 #(.INIT(32'h96696996)) lut_n7013 (.I0(x1857), .I1(x1858), .I2(x1859), .I3(n7009), .I4(n7010), .O(n7013));
  LUT5 #(.INIT(32'hFF969600)) lut_n7014 (.I0(x1863), .I1(x1864), .I2(x1865), .I3(n7012), .I4(n7013), .O(n7014));
  LUT3 #(.INIT(8'h96)) lut_n7015 (.I0(n7003), .I1(n7006), .I2(n7007), .O(n7015));
  LUT3 #(.INIT(8'hE8)) lut_n7016 (.I0(n7011), .I1(n7014), .I2(n7015), .O(n7016));
  LUT3 #(.INIT(8'h96)) lut_n7017 (.I0(n6990), .I1(n6998), .I2(n6999), .O(n7017));
  LUT3 #(.INIT(8'hE8)) lut_n7018 (.I0(n7008), .I1(n7016), .I2(n7017), .O(n7018));
  LUT3 #(.INIT(8'h96)) lut_n7019 (.I0(n6962), .I1(n6980), .I2(n6981), .O(n7019));
  LUT3 #(.INIT(8'hE8)) lut_n7020 (.I0(n7000), .I1(n7018), .I2(n7019), .O(n7020));
  LUT3 #(.INIT(8'h96)) lut_n7021 (.I0(n6904), .I1(n6942), .I2(n6943), .O(n7021));
  LUT3 #(.INIT(8'hE8)) lut_n7022 (.I0(n6982), .I1(n7020), .I2(n7021), .O(n7022));
  LUT3 #(.INIT(8'h96)) lut_n7023 (.I0(n6780), .I1(n6858), .I2(n6859), .O(n7023));
  LUT3 #(.INIT(8'hE8)) lut_n7024 (.I0(n6944), .I1(n7022), .I2(n7023), .O(n7024));
  LUT3 #(.INIT(8'h96)) lut_n7025 (.I0(x1872), .I1(x1873), .I2(x1874), .O(n7025));
  LUT5 #(.INIT(32'h96696996)) lut_n7026 (.I0(x1863), .I1(x1864), .I2(x1865), .I3(n7012), .I4(n7013), .O(n7026));
  LUT5 #(.INIT(32'hFF969600)) lut_n7027 (.I0(x1869), .I1(x1870), .I2(x1871), .I3(n7025), .I4(n7026), .O(n7027));
  LUT3 #(.INIT(8'h96)) lut_n7028 (.I0(x1878), .I1(x1879), .I2(x1880), .O(n7028));
  LUT5 #(.INIT(32'h96696996)) lut_n7029 (.I0(x1869), .I1(x1870), .I2(x1871), .I3(n7025), .I4(n7026), .O(n7029));
  LUT5 #(.INIT(32'hFF969600)) lut_n7030 (.I0(x1875), .I1(x1876), .I2(x1877), .I3(n7028), .I4(n7029), .O(n7030));
  LUT3 #(.INIT(8'h96)) lut_n7031 (.I0(n7011), .I1(n7014), .I2(n7015), .O(n7031));
  LUT3 #(.INIT(8'hE8)) lut_n7032 (.I0(n7027), .I1(n7030), .I2(n7031), .O(n7032));
  LUT3 #(.INIT(8'h96)) lut_n7033 (.I0(x1884), .I1(x1885), .I2(x1886), .O(n7033));
  LUT5 #(.INIT(32'h96696996)) lut_n7034 (.I0(x1875), .I1(x1876), .I2(x1877), .I3(n7028), .I4(n7029), .O(n7034));
  LUT5 #(.INIT(32'hFF969600)) lut_n7035 (.I0(x1881), .I1(x1882), .I2(x1883), .I3(n7033), .I4(n7034), .O(n7035));
  LUT3 #(.INIT(8'h96)) lut_n7036 (.I0(x1890), .I1(x1891), .I2(x1892), .O(n7036));
  LUT5 #(.INIT(32'h96696996)) lut_n7037 (.I0(x1881), .I1(x1882), .I2(x1883), .I3(n7033), .I4(n7034), .O(n7037));
  LUT5 #(.INIT(32'hFF969600)) lut_n7038 (.I0(x1887), .I1(x1888), .I2(x1889), .I3(n7036), .I4(n7037), .O(n7038));
  LUT3 #(.INIT(8'h96)) lut_n7039 (.I0(n7027), .I1(n7030), .I2(n7031), .O(n7039));
  LUT3 #(.INIT(8'hE8)) lut_n7040 (.I0(n7035), .I1(n7038), .I2(n7039), .O(n7040));
  LUT3 #(.INIT(8'h96)) lut_n7041 (.I0(n7008), .I1(n7016), .I2(n7017), .O(n7041));
  LUT3 #(.INIT(8'hE8)) lut_n7042 (.I0(n7032), .I1(n7040), .I2(n7041), .O(n7042));
  LUT3 #(.INIT(8'h96)) lut_n7043 (.I0(x1896), .I1(x1897), .I2(x1898), .O(n7043));
  LUT5 #(.INIT(32'h96696996)) lut_n7044 (.I0(x1887), .I1(x1888), .I2(x1889), .I3(n7036), .I4(n7037), .O(n7044));
  LUT5 #(.INIT(32'hFF969600)) lut_n7045 (.I0(x1893), .I1(x1894), .I2(x1895), .I3(n7043), .I4(n7044), .O(n7045));
  LUT3 #(.INIT(8'h96)) lut_n7046 (.I0(x1902), .I1(x1903), .I2(x1904), .O(n7046));
  LUT5 #(.INIT(32'h96696996)) lut_n7047 (.I0(x1893), .I1(x1894), .I2(x1895), .I3(n7043), .I4(n7044), .O(n7047));
  LUT5 #(.INIT(32'hFF969600)) lut_n7048 (.I0(x1899), .I1(x1900), .I2(x1901), .I3(n7046), .I4(n7047), .O(n7048));
  LUT3 #(.INIT(8'h96)) lut_n7049 (.I0(n7035), .I1(n7038), .I2(n7039), .O(n7049));
  LUT3 #(.INIT(8'hE8)) lut_n7050 (.I0(n7045), .I1(n7048), .I2(n7049), .O(n7050));
  LUT3 #(.INIT(8'h96)) lut_n7051 (.I0(x1908), .I1(x1909), .I2(x1910), .O(n7051));
  LUT5 #(.INIT(32'h96696996)) lut_n7052 (.I0(x1899), .I1(x1900), .I2(x1901), .I3(n7046), .I4(n7047), .O(n7052));
  LUT5 #(.INIT(32'hFF969600)) lut_n7053 (.I0(x1905), .I1(x1906), .I2(x1907), .I3(n7051), .I4(n7052), .O(n7053));
  LUT3 #(.INIT(8'h96)) lut_n7054 (.I0(x1914), .I1(x1915), .I2(x1916), .O(n7054));
  LUT5 #(.INIT(32'h96696996)) lut_n7055 (.I0(x1905), .I1(x1906), .I2(x1907), .I3(n7051), .I4(n7052), .O(n7055));
  LUT5 #(.INIT(32'hFF969600)) lut_n7056 (.I0(x1911), .I1(x1912), .I2(x1913), .I3(n7054), .I4(n7055), .O(n7056));
  LUT3 #(.INIT(8'h96)) lut_n7057 (.I0(n7045), .I1(n7048), .I2(n7049), .O(n7057));
  LUT3 #(.INIT(8'hE8)) lut_n7058 (.I0(n7053), .I1(n7056), .I2(n7057), .O(n7058));
  LUT3 #(.INIT(8'h96)) lut_n7059 (.I0(n7032), .I1(n7040), .I2(n7041), .O(n7059));
  LUT3 #(.INIT(8'hE8)) lut_n7060 (.I0(n7050), .I1(n7058), .I2(n7059), .O(n7060));
  LUT3 #(.INIT(8'h96)) lut_n7061 (.I0(n7000), .I1(n7018), .I2(n7019), .O(n7061));
  LUT3 #(.INIT(8'hE8)) lut_n7062 (.I0(n7042), .I1(n7060), .I2(n7061), .O(n7062));
  LUT3 #(.INIT(8'h96)) lut_n7063 (.I0(x1920), .I1(x1921), .I2(x1922), .O(n7063));
  LUT5 #(.INIT(32'h96696996)) lut_n7064 (.I0(x1911), .I1(x1912), .I2(x1913), .I3(n7054), .I4(n7055), .O(n7064));
  LUT5 #(.INIT(32'hFF969600)) lut_n7065 (.I0(x1917), .I1(x1918), .I2(x1919), .I3(n7063), .I4(n7064), .O(n7065));
  LUT3 #(.INIT(8'h96)) lut_n7066 (.I0(x1926), .I1(x1927), .I2(x1928), .O(n7066));
  LUT5 #(.INIT(32'h96696996)) lut_n7067 (.I0(x1917), .I1(x1918), .I2(x1919), .I3(n7063), .I4(n7064), .O(n7067));
  LUT5 #(.INIT(32'hFF969600)) lut_n7068 (.I0(x1923), .I1(x1924), .I2(x1925), .I3(n7066), .I4(n7067), .O(n7068));
  LUT3 #(.INIT(8'h96)) lut_n7069 (.I0(n7053), .I1(n7056), .I2(n7057), .O(n7069));
  LUT3 #(.INIT(8'hE8)) lut_n7070 (.I0(n7065), .I1(n7068), .I2(n7069), .O(n7070));
  LUT3 #(.INIT(8'h96)) lut_n7071 (.I0(x1932), .I1(x1933), .I2(x1934), .O(n7071));
  LUT5 #(.INIT(32'h96696996)) lut_n7072 (.I0(x1923), .I1(x1924), .I2(x1925), .I3(n7066), .I4(n7067), .O(n7072));
  LUT5 #(.INIT(32'hFF969600)) lut_n7073 (.I0(x1929), .I1(x1930), .I2(x1931), .I3(n7071), .I4(n7072), .O(n7073));
  LUT3 #(.INIT(8'h96)) lut_n7074 (.I0(x1938), .I1(x1939), .I2(x1940), .O(n7074));
  LUT5 #(.INIT(32'h96696996)) lut_n7075 (.I0(x1929), .I1(x1930), .I2(x1931), .I3(n7071), .I4(n7072), .O(n7075));
  LUT5 #(.INIT(32'hFF969600)) lut_n7076 (.I0(x1935), .I1(x1936), .I2(x1937), .I3(n7074), .I4(n7075), .O(n7076));
  LUT3 #(.INIT(8'h96)) lut_n7077 (.I0(n7065), .I1(n7068), .I2(n7069), .O(n7077));
  LUT3 #(.INIT(8'hE8)) lut_n7078 (.I0(n7073), .I1(n7076), .I2(n7077), .O(n7078));
  LUT3 #(.INIT(8'h96)) lut_n7079 (.I0(n7050), .I1(n7058), .I2(n7059), .O(n7079));
  LUT3 #(.INIT(8'hE8)) lut_n7080 (.I0(n7070), .I1(n7078), .I2(n7079), .O(n7080));
  LUT3 #(.INIT(8'h96)) lut_n7081 (.I0(x1944), .I1(x1945), .I2(x1946), .O(n7081));
  LUT5 #(.INIT(32'h96696996)) lut_n7082 (.I0(x1935), .I1(x1936), .I2(x1937), .I3(n7074), .I4(n7075), .O(n7082));
  LUT5 #(.INIT(32'hFF969600)) lut_n7083 (.I0(x1941), .I1(x1942), .I2(x1943), .I3(n7081), .I4(n7082), .O(n7083));
  LUT3 #(.INIT(8'h96)) lut_n7084 (.I0(x1950), .I1(x1951), .I2(x1952), .O(n7084));
  LUT5 #(.INIT(32'h96696996)) lut_n7085 (.I0(x1941), .I1(x1942), .I2(x1943), .I3(n7081), .I4(n7082), .O(n7085));
  LUT5 #(.INIT(32'hFF969600)) lut_n7086 (.I0(x1947), .I1(x1948), .I2(x1949), .I3(n7084), .I4(n7085), .O(n7086));
  LUT3 #(.INIT(8'h96)) lut_n7087 (.I0(n7073), .I1(n7076), .I2(n7077), .O(n7087));
  LUT3 #(.INIT(8'hE8)) lut_n7088 (.I0(n7083), .I1(n7086), .I2(n7087), .O(n7088));
  LUT3 #(.INIT(8'h96)) lut_n7089 (.I0(x1956), .I1(x1957), .I2(x1958), .O(n7089));
  LUT5 #(.INIT(32'h96696996)) lut_n7090 (.I0(x1947), .I1(x1948), .I2(x1949), .I3(n7084), .I4(n7085), .O(n7090));
  LUT5 #(.INIT(32'hFF969600)) lut_n7091 (.I0(x1953), .I1(x1954), .I2(x1955), .I3(n7089), .I4(n7090), .O(n7091));
  LUT3 #(.INIT(8'h96)) lut_n7092 (.I0(x1962), .I1(x1963), .I2(x1964), .O(n7092));
  LUT5 #(.INIT(32'h96696996)) lut_n7093 (.I0(x1953), .I1(x1954), .I2(x1955), .I3(n7089), .I4(n7090), .O(n7093));
  LUT5 #(.INIT(32'hFF969600)) lut_n7094 (.I0(x1959), .I1(x1960), .I2(x1961), .I3(n7092), .I4(n7093), .O(n7094));
  LUT3 #(.INIT(8'h96)) lut_n7095 (.I0(n7083), .I1(n7086), .I2(n7087), .O(n7095));
  LUT3 #(.INIT(8'hE8)) lut_n7096 (.I0(n7091), .I1(n7094), .I2(n7095), .O(n7096));
  LUT3 #(.INIT(8'h96)) lut_n7097 (.I0(n7070), .I1(n7078), .I2(n7079), .O(n7097));
  LUT3 #(.INIT(8'hE8)) lut_n7098 (.I0(n7088), .I1(n7096), .I2(n7097), .O(n7098));
  LUT3 #(.INIT(8'h96)) lut_n7099 (.I0(n7042), .I1(n7060), .I2(n7061), .O(n7099));
  LUT3 #(.INIT(8'hE8)) lut_n7100 (.I0(n7080), .I1(n7098), .I2(n7099), .O(n7100));
  LUT3 #(.INIT(8'h96)) lut_n7101 (.I0(n6982), .I1(n7020), .I2(n7021), .O(n7101));
  LUT3 #(.INIT(8'hE8)) lut_n7102 (.I0(n7062), .I1(n7100), .I2(n7101), .O(n7102));
  LUT3 #(.INIT(8'h96)) lut_n7103 (.I0(x1968), .I1(x1969), .I2(x1970), .O(n7103));
  LUT5 #(.INIT(32'h96696996)) lut_n7104 (.I0(x1959), .I1(x1960), .I2(x1961), .I3(n7092), .I4(n7093), .O(n7104));
  LUT5 #(.INIT(32'hFF969600)) lut_n7105 (.I0(x1965), .I1(x1966), .I2(x1967), .I3(n7103), .I4(n7104), .O(n7105));
  LUT3 #(.INIT(8'h96)) lut_n7106 (.I0(x1974), .I1(x1975), .I2(x1976), .O(n7106));
  LUT5 #(.INIT(32'h96696996)) lut_n7107 (.I0(x1965), .I1(x1966), .I2(x1967), .I3(n7103), .I4(n7104), .O(n7107));
  LUT5 #(.INIT(32'hFF969600)) lut_n7108 (.I0(x1971), .I1(x1972), .I2(x1973), .I3(n7106), .I4(n7107), .O(n7108));
  LUT3 #(.INIT(8'h96)) lut_n7109 (.I0(n7091), .I1(n7094), .I2(n7095), .O(n7109));
  LUT3 #(.INIT(8'hE8)) lut_n7110 (.I0(n7105), .I1(n7108), .I2(n7109), .O(n7110));
  LUT3 #(.INIT(8'h96)) lut_n7111 (.I0(x1980), .I1(x1981), .I2(x1982), .O(n7111));
  LUT5 #(.INIT(32'h96696996)) lut_n7112 (.I0(x1971), .I1(x1972), .I2(x1973), .I3(n7106), .I4(n7107), .O(n7112));
  LUT5 #(.INIT(32'hFF969600)) lut_n7113 (.I0(x1977), .I1(x1978), .I2(x1979), .I3(n7111), .I4(n7112), .O(n7113));
  LUT3 #(.INIT(8'h96)) lut_n7114 (.I0(x1986), .I1(x1987), .I2(x1988), .O(n7114));
  LUT5 #(.INIT(32'h96696996)) lut_n7115 (.I0(x1977), .I1(x1978), .I2(x1979), .I3(n7111), .I4(n7112), .O(n7115));
  LUT5 #(.INIT(32'hFF969600)) lut_n7116 (.I0(x1983), .I1(x1984), .I2(x1985), .I3(n7114), .I4(n7115), .O(n7116));
  LUT3 #(.INIT(8'h96)) lut_n7117 (.I0(n7105), .I1(n7108), .I2(n7109), .O(n7117));
  LUT3 #(.INIT(8'hE8)) lut_n7118 (.I0(n7113), .I1(n7116), .I2(n7117), .O(n7118));
  LUT3 #(.INIT(8'h96)) lut_n7119 (.I0(n7088), .I1(n7096), .I2(n7097), .O(n7119));
  LUT3 #(.INIT(8'hE8)) lut_n7120 (.I0(n7110), .I1(n7118), .I2(n7119), .O(n7120));
  LUT3 #(.INIT(8'h96)) lut_n7121 (.I0(x1992), .I1(x1993), .I2(x1994), .O(n7121));
  LUT5 #(.INIT(32'h96696996)) lut_n7122 (.I0(x1983), .I1(x1984), .I2(x1985), .I3(n7114), .I4(n7115), .O(n7122));
  LUT5 #(.INIT(32'hFF969600)) lut_n7123 (.I0(x1989), .I1(x1990), .I2(x1991), .I3(n7121), .I4(n7122), .O(n7123));
  LUT3 #(.INIT(8'h96)) lut_n7124 (.I0(x1998), .I1(x1999), .I2(x2000), .O(n7124));
  LUT5 #(.INIT(32'h96696996)) lut_n7125 (.I0(x1989), .I1(x1990), .I2(x1991), .I3(n7121), .I4(n7122), .O(n7125));
  LUT5 #(.INIT(32'hFF969600)) lut_n7126 (.I0(x1995), .I1(x1996), .I2(x1997), .I3(n7124), .I4(n7125), .O(n7126));
  LUT3 #(.INIT(8'h96)) lut_n7127 (.I0(n7113), .I1(n7116), .I2(n7117), .O(n7127));
  LUT3 #(.INIT(8'hE8)) lut_n7128 (.I0(n7123), .I1(n7126), .I2(n7127), .O(n7128));
  LUT3 #(.INIT(8'h96)) lut_n7129 (.I0(x2004), .I1(x2005), .I2(x2006), .O(n7129));
  LUT5 #(.INIT(32'h96696996)) lut_n7130 (.I0(x1995), .I1(x1996), .I2(x1997), .I3(n7124), .I4(n7125), .O(n7130));
  LUT5 #(.INIT(32'hFF969600)) lut_n7131 (.I0(x2001), .I1(x2002), .I2(x2003), .I3(n7129), .I4(n7130), .O(n7131));
  LUT3 #(.INIT(8'h96)) lut_n7132 (.I0(x2010), .I1(x2011), .I2(x2012), .O(n7132));
  LUT5 #(.INIT(32'h96696996)) lut_n7133 (.I0(x2001), .I1(x2002), .I2(x2003), .I3(n7129), .I4(n7130), .O(n7133));
  LUT5 #(.INIT(32'hFF969600)) lut_n7134 (.I0(x2007), .I1(x2008), .I2(x2009), .I3(n7132), .I4(n7133), .O(n7134));
  LUT3 #(.INIT(8'h96)) lut_n7135 (.I0(n7123), .I1(n7126), .I2(n7127), .O(n7135));
  LUT3 #(.INIT(8'hE8)) lut_n7136 (.I0(n7131), .I1(n7134), .I2(n7135), .O(n7136));
  LUT3 #(.INIT(8'h96)) lut_n7137 (.I0(n7110), .I1(n7118), .I2(n7119), .O(n7137));
  LUT3 #(.INIT(8'hE8)) lut_n7138 (.I0(n7128), .I1(n7136), .I2(n7137), .O(n7138));
  LUT3 #(.INIT(8'h96)) lut_n7139 (.I0(n7080), .I1(n7098), .I2(n7099), .O(n7139));
  LUT3 #(.INIT(8'hE8)) lut_n7140 (.I0(n7120), .I1(n7138), .I2(n7139), .O(n7140));
  LUT3 #(.INIT(8'h96)) lut_n7141 (.I0(x2016), .I1(x2017), .I2(x2018), .O(n7141));
  LUT5 #(.INIT(32'h96696996)) lut_n7142 (.I0(x2007), .I1(x2008), .I2(x2009), .I3(n7132), .I4(n7133), .O(n7142));
  LUT5 #(.INIT(32'hFF969600)) lut_n7143 (.I0(x2013), .I1(x2014), .I2(x2015), .I3(n7141), .I4(n7142), .O(n7143));
  LUT3 #(.INIT(8'h96)) lut_n7144 (.I0(x2022), .I1(x2023), .I2(x2024), .O(n7144));
  LUT5 #(.INIT(32'h96696996)) lut_n7145 (.I0(x2013), .I1(x2014), .I2(x2015), .I3(n7141), .I4(n7142), .O(n7145));
  LUT5 #(.INIT(32'hFF969600)) lut_n7146 (.I0(x2019), .I1(x2020), .I2(x2021), .I3(n7144), .I4(n7145), .O(n7146));
  LUT3 #(.INIT(8'h96)) lut_n7147 (.I0(n7131), .I1(n7134), .I2(n7135), .O(n7147));
  LUT3 #(.INIT(8'hE8)) lut_n7148 (.I0(n7143), .I1(n7146), .I2(n7147), .O(n7148));
  LUT3 #(.INIT(8'h96)) lut_n7149 (.I0(x2028), .I1(x2029), .I2(x2030), .O(n7149));
  LUT5 #(.INIT(32'h96696996)) lut_n7150 (.I0(x2019), .I1(x2020), .I2(x2021), .I3(n7144), .I4(n7145), .O(n7150));
  LUT5 #(.INIT(32'hFF969600)) lut_n7151 (.I0(x2025), .I1(x2026), .I2(x2027), .I3(n7149), .I4(n7150), .O(n7151));
  LUT3 #(.INIT(8'h96)) lut_n7152 (.I0(x2034), .I1(x2035), .I2(x2036), .O(n7152));
  LUT5 #(.INIT(32'h96696996)) lut_n7153 (.I0(x2025), .I1(x2026), .I2(x2027), .I3(n7149), .I4(n7150), .O(n7153));
  LUT5 #(.INIT(32'hFF969600)) lut_n7154 (.I0(x2031), .I1(x2032), .I2(x2033), .I3(n7152), .I4(n7153), .O(n7154));
  LUT3 #(.INIT(8'h96)) lut_n7155 (.I0(n7143), .I1(n7146), .I2(n7147), .O(n7155));
  LUT3 #(.INIT(8'hE8)) lut_n7156 (.I0(n7151), .I1(n7154), .I2(n7155), .O(n7156));
  LUT3 #(.INIT(8'h96)) lut_n7157 (.I0(n7128), .I1(n7136), .I2(n7137), .O(n7157));
  LUT3 #(.INIT(8'hE8)) lut_n7158 (.I0(n7148), .I1(n7156), .I2(n7157), .O(n7158));
  LUT3 #(.INIT(8'h96)) lut_n7159 (.I0(x2040), .I1(x2041), .I2(x2042), .O(n7159));
  LUT5 #(.INIT(32'h96696996)) lut_n7160 (.I0(x2031), .I1(x2032), .I2(x2033), .I3(n7152), .I4(n7153), .O(n7160));
  LUT5 #(.INIT(32'hFF969600)) lut_n7161 (.I0(x2037), .I1(x2038), .I2(x2039), .I3(n7159), .I4(n7160), .O(n7161));
  LUT3 #(.INIT(8'h96)) lut_n7162 (.I0(x2046), .I1(x2047), .I2(x2048), .O(n7162));
  LUT5 #(.INIT(32'h96696996)) lut_n7163 (.I0(x2037), .I1(x2038), .I2(x2039), .I3(n7159), .I4(n7160), .O(n7163));
  LUT5 #(.INIT(32'hFF969600)) lut_n7164 (.I0(x2043), .I1(x2044), .I2(x2045), .I3(n7162), .I4(n7163), .O(n7164));
  LUT3 #(.INIT(8'h96)) lut_n7165 (.I0(n7151), .I1(n7154), .I2(n7155), .O(n7165));
  LUT3 #(.INIT(8'hE8)) lut_n7166 (.I0(n7161), .I1(n7164), .I2(n7165), .O(n7166));
  LUT3 #(.INIT(8'h96)) lut_n7167 (.I0(x2052), .I1(x2053), .I2(x2054), .O(n7167));
  LUT5 #(.INIT(32'h96696996)) lut_n7168 (.I0(x2043), .I1(x2044), .I2(x2045), .I3(n7162), .I4(n7163), .O(n7168));
  LUT5 #(.INIT(32'hFF969600)) lut_n7169 (.I0(x2049), .I1(x2050), .I2(x2051), .I3(n7167), .I4(n7168), .O(n7169));
  LUT3 #(.INIT(8'h96)) lut_n7170 (.I0(x2058), .I1(x2059), .I2(x2060), .O(n7170));
  LUT5 #(.INIT(32'h96696996)) lut_n7171 (.I0(x2049), .I1(x2050), .I2(x2051), .I3(n7167), .I4(n7168), .O(n7171));
  LUT5 #(.INIT(32'hFF969600)) lut_n7172 (.I0(x2055), .I1(x2056), .I2(x2057), .I3(n7170), .I4(n7171), .O(n7172));
  LUT3 #(.INIT(8'h96)) lut_n7173 (.I0(n7161), .I1(n7164), .I2(n7165), .O(n7173));
  LUT3 #(.INIT(8'hE8)) lut_n7174 (.I0(n7169), .I1(n7172), .I2(n7173), .O(n7174));
  LUT3 #(.INIT(8'h96)) lut_n7175 (.I0(n7148), .I1(n7156), .I2(n7157), .O(n7175));
  LUT3 #(.INIT(8'hE8)) lut_n7176 (.I0(n7166), .I1(n7174), .I2(n7175), .O(n7176));
  LUT3 #(.INIT(8'h96)) lut_n7177 (.I0(n7120), .I1(n7138), .I2(n7139), .O(n7177));
  LUT3 #(.INIT(8'hE8)) lut_n7178 (.I0(n7158), .I1(n7176), .I2(n7177), .O(n7178));
  LUT3 #(.INIT(8'h96)) lut_n7179 (.I0(n7062), .I1(n7100), .I2(n7101), .O(n7179));
  LUT3 #(.INIT(8'hE8)) lut_n7180 (.I0(n7140), .I1(n7178), .I2(n7179), .O(n7180));
  LUT3 #(.INIT(8'h96)) lut_n7181 (.I0(n6944), .I1(n7022), .I2(n7023), .O(n7181));
  LUT3 #(.INIT(8'hE8)) lut_n7182 (.I0(n7102), .I1(n7180), .I2(n7181), .O(n7182));
  LUT3 #(.INIT(8'h96)) lut_n7183 (.I0(n6702), .I1(n6860), .I2(n6861), .O(n7183));
  LUT3 #(.INIT(8'hE8)) lut_n7184 (.I0(n7024), .I1(n7182), .I2(n7183), .O(n7184));
  LUT3 #(.INIT(8'h96)) lut_n7185 (.I0(x2064), .I1(x2065), .I2(x2066), .O(n7185));
  LUT5 #(.INIT(32'h96696996)) lut_n7186 (.I0(x2055), .I1(x2056), .I2(x2057), .I3(n7170), .I4(n7171), .O(n7186));
  LUT5 #(.INIT(32'hFF969600)) lut_n7187 (.I0(x2061), .I1(x2062), .I2(x2063), .I3(n7185), .I4(n7186), .O(n7187));
  LUT3 #(.INIT(8'h96)) lut_n7188 (.I0(x2070), .I1(x2071), .I2(x2072), .O(n7188));
  LUT5 #(.INIT(32'h96696996)) lut_n7189 (.I0(x2061), .I1(x2062), .I2(x2063), .I3(n7185), .I4(n7186), .O(n7189));
  LUT5 #(.INIT(32'hFF969600)) lut_n7190 (.I0(x2067), .I1(x2068), .I2(x2069), .I3(n7188), .I4(n7189), .O(n7190));
  LUT3 #(.INIT(8'h96)) lut_n7191 (.I0(n7169), .I1(n7172), .I2(n7173), .O(n7191));
  LUT3 #(.INIT(8'hE8)) lut_n7192 (.I0(n7187), .I1(n7190), .I2(n7191), .O(n7192));
  LUT3 #(.INIT(8'h96)) lut_n7193 (.I0(x2076), .I1(x2077), .I2(x2078), .O(n7193));
  LUT5 #(.INIT(32'h96696996)) lut_n7194 (.I0(x2067), .I1(x2068), .I2(x2069), .I3(n7188), .I4(n7189), .O(n7194));
  LUT5 #(.INIT(32'hFF969600)) lut_n7195 (.I0(x2073), .I1(x2074), .I2(x2075), .I3(n7193), .I4(n7194), .O(n7195));
  LUT3 #(.INIT(8'h96)) lut_n7196 (.I0(x2082), .I1(x2083), .I2(x2084), .O(n7196));
  LUT5 #(.INIT(32'h96696996)) lut_n7197 (.I0(x2073), .I1(x2074), .I2(x2075), .I3(n7193), .I4(n7194), .O(n7197));
  LUT5 #(.INIT(32'hFF969600)) lut_n7198 (.I0(x2079), .I1(x2080), .I2(x2081), .I3(n7196), .I4(n7197), .O(n7198));
  LUT3 #(.INIT(8'h96)) lut_n7199 (.I0(n7187), .I1(n7190), .I2(n7191), .O(n7199));
  LUT3 #(.INIT(8'hE8)) lut_n7200 (.I0(n7195), .I1(n7198), .I2(n7199), .O(n7200));
  LUT3 #(.INIT(8'h96)) lut_n7201 (.I0(n7166), .I1(n7174), .I2(n7175), .O(n7201));
  LUT3 #(.INIT(8'hE8)) lut_n7202 (.I0(n7192), .I1(n7200), .I2(n7201), .O(n7202));
  LUT3 #(.INIT(8'h96)) lut_n7203 (.I0(x2088), .I1(x2089), .I2(x2090), .O(n7203));
  LUT5 #(.INIT(32'h96696996)) lut_n7204 (.I0(x2079), .I1(x2080), .I2(x2081), .I3(n7196), .I4(n7197), .O(n7204));
  LUT5 #(.INIT(32'hFF969600)) lut_n7205 (.I0(x2085), .I1(x2086), .I2(x2087), .I3(n7203), .I4(n7204), .O(n7205));
  LUT3 #(.INIT(8'h96)) lut_n7206 (.I0(x2094), .I1(x2095), .I2(x2096), .O(n7206));
  LUT5 #(.INIT(32'h96696996)) lut_n7207 (.I0(x2085), .I1(x2086), .I2(x2087), .I3(n7203), .I4(n7204), .O(n7207));
  LUT5 #(.INIT(32'hFF969600)) lut_n7208 (.I0(x2091), .I1(x2092), .I2(x2093), .I3(n7206), .I4(n7207), .O(n7208));
  LUT3 #(.INIT(8'h96)) lut_n7209 (.I0(n7195), .I1(n7198), .I2(n7199), .O(n7209));
  LUT3 #(.INIT(8'hE8)) lut_n7210 (.I0(n7205), .I1(n7208), .I2(n7209), .O(n7210));
  LUT3 #(.INIT(8'h96)) lut_n7211 (.I0(x2100), .I1(x2101), .I2(x2102), .O(n7211));
  LUT5 #(.INIT(32'h96696996)) lut_n7212 (.I0(x2091), .I1(x2092), .I2(x2093), .I3(n7206), .I4(n7207), .O(n7212));
  LUT5 #(.INIT(32'hFF969600)) lut_n7213 (.I0(x2097), .I1(x2098), .I2(x2099), .I3(n7211), .I4(n7212), .O(n7213));
  LUT3 #(.INIT(8'h96)) lut_n7214 (.I0(x2106), .I1(x2107), .I2(x2108), .O(n7214));
  LUT5 #(.INIT(32'h96696996)) lut_n7215 (.I0(x2097), .I1(x2098), .I2(x2099), .I3(n7211), .I4(n7212), .O(n7215));
  LUT5 #(.INIT(32'hFF969600)) lut_n7216 (.I0(x2103), .I1(x2104), .I2(x2105), .I3(n7214), .I4(n7215), .O(n7216));
  LUT3 #(.INIT(8'h96)) lut_n7217 (.I0(n7205), .I1(n7208), .I2(n7209), .O(n7217));
  LUT3 #(.INIT(8'hE8)) lut_n7218 (.I0(n7213), .I1(n7216), .I2(n7217), .O(n7218));
  LUT3 #(.INIT(8'h96)) lut_n7219 (.I0(n7192), .I1(n7200), .I2(n7201), .O(n7219));
  LUT3 #(.INIT(8'hE8)) lut_n7220 (.I0(n7210), .I1(n7218), .I2(n7219), .O(n7220));
  LUT3 #(.INIT(8'h96)) lut_n7221 (.I0(n7158), .I1(n7176), .I2(n7177), .O(n7221));
  LUT3 #(.INIT(8'hE8)) lut_n7222 (.I0(n7202), .I1(n7220), .I2(n7221), .O(n7222));
  LUT3 #(.INIT(8'h96)) lut_n7223 (.I0(x2112), .I1(x2113), .I2(x2114), .O(n7223));
  LUT5 #(.INIT(32'h96696996)) lut_n7224 (.I0(x2103), .I1(x2104), .I2(x2105), .I3(n7214), .I4(n7215), .O(n7224));
  LUT5 #(.INIT(32'hFF969600)) lut_n7225 (.I0(x2109), .I1(x2110), .I2(x2111), .I3(n7223), .I4(n7224), .O(n7225));
  LUT3 #(.INIT(8'h96)) lut_n7226 (.I0(x2118), .I1(x2119), .I2(x2120), .O(n7226));
  LUT5 #(.INIT(32'h96696996)) lut_n7227 (.I0(x2109), .I1(x2110), .I2(x2111), .I3(n7223), .I4(n7224), .O(n7227));
  LUT5 #(.INIT(32'hFF969600)) lut_n7228 (.I0(x2115), .I1(x2116), .I2(x2117), .I3(n7226), .I4(n7227), .O(n7228));
  LUT3 #(.INIT(8'h96)) lut_n7229 (.I0(n7213), .I1(n7216), .I2(n7217), .O(n7229));
  LUT3 #(.INIT(8'hE8)) lut_n7230 (.I0(n7225), .I1(n7228), .I2(n7229), .O(n7230));
  LUT3 #(.INIT(8'h96)) lut_n7231 (.I0(x2124), .I1(x2125), .I2(x2126), .O(n7231));
  LUT5 #(.INIT(32'h96696996)) lut_n7232 (.I0(x2115), .I1(x2116), .I2(x2117), .I3(n7226), .I4(n7227), .O(n7232));
  LUT5 #(.INIT(32'hFF969600)) lut_n7233 (.I0(x2121), .I1(x2122), .I2(x2123), .I3(n7231), .I4(n7232), .O(n7233));
  LUT3 #(.INIT(8'h96)) lut_n7234 (.I0(x2130), .I1(x2131), .I2(x2132), .O(n7234));
  LUT5 #(.INIT(32'h96696996)) lut_n7235 (.I0(x2121), .I1(x2122), .I2(x2123), .I3(n7231), .I4(n7232), .O(n7235));
  LUT5 #(.INIT(32'hFF969600)) lut_n7236 (.I0(x2127), .I1(x2128), .I2(x2129), .I3(n7234), .I4(n7235), .O(n7236));
  LUT3 #(.INIT(8'h96)) lut_n7237 (.I0(n7225), .I1(n7228), .I2(n7229), .O(n7237));
  LUT3 #(.INIT(8'hE8)) lut_n7238 (.I0(n7233), .I1(n7236), .I2(n7237), .O(n7238));
  LUT3 #(.INIT(8'h96)) lut_n7239 (.I0(n7210), .I1(n7218), .I2(n7219), .O(n7239));
  LUT3 #(.INIT(8'hE8)) lut_n7240 (.I0(n7230), .I1(n7238), .I2(n7239), .O(n7240));
  LUT3 #(.INIT(8'h96)) lut_n7241 (.I0(x2136), .I1(x2137), .I2(x2138), .O(n7241));
  LUT5 #(.INIT(32'h96696996)) lut_n7242 (.I0(x2127), .I1(x2128), .I2(x2129), .I3(n7234), .I4(n7235), .O(n7242));
  LUT5 #(.INIT(32'hFF969600)) lut_n7243 (.I0(x2133), .I1(x2134), .I2(x2135), .I3(n7241), .I4(n7242), .O(n7243));
  LUT3 #(.INIT(8'h96)) lut_n7244 (.I0(x2142), .I1(x2143), .I2(x2144), .O(n7244));
  LUT5 #(.INIT(32'h96696996)) lut_n7245 (.I0(x2133), .I1(x2134), .I2(x2135), .I3(n7241), .I4(n7242), .O(n7245));
  LUT5 #(.INIT(32'hFF969600)) lut_n7246 (.I0(x2139), .I1(x2140), .I2(x2141), .I3(n7244), .I4(n7245), .O(n7246));
  LUT3 #(.INIT(8'h96)) lut_n7247 (.I0(n7233), .I1(n7236), .I2(n7237), .O(n7247));
  LUT3 #(.INIT(8'hE8)) lut_n7248 (.I0(n7243), .I1(n7246), .I2(n7247), .O(n7248));
  LUT3 #(.INIT(8'h96)) lut_n7249 (.I0(x2148), .I1(x2149), .I2(x2150), .O(n7249));
  LUT5 #(.INIT(32'h96696996)) lut_n7250 (.I0(x2139), .I1(x2140), .I2(x2141), .I3(n7244), .I4(n7245), .O(n7250));
  LUT5 #(.INIT(32'hFF969600)) lut_n7251 (.I0(x2145), .I1(x2146), .I2(x2147), .I3(n7249), .I4(n7250), .O(n7251));
  LUT3 #(.INIT(8'h96)) lut_n7252 (.I0(x2154), .I1(x2155), .I2(x2156), .O(n7252));
  LUT5 #(.INIT(32'h96696996)) lut_n7253 (.I0(x2145), .I1(x2146), .I2(x2147), .I3(n7249), .I4(n7250), .O(n7253));
  LUT5 #(.INIT(32'hFF969600)) lut_n7254 (.I0(x2151), .I1(x2152), .I2(x2153), .I3(n7252), .I4(n7253), .O(n7254));
  LUT3 #(.INIT(8'h96)) lut_n7255 (.I0(n7243), .I1(n7246), .I2(n7247), .O(n7255));
  LUT3 #(.INIT(8'hE8)) lut_n7256 (.I0(n7251), .I1(n7254), .I2(n7255), .O(n7256));
  LUT3 #(.INIT(8'h96)) lut_n7257 (.I0(n7230), .I1(n7238), .I2(n7239), .O(n7257));
  LUT3 #(.INIT(8'hE8)) lut_n7258 (.I0(n7248), .I1(n7256), .I2(n7257), .O(n7258));
  LUT3 #(.INIT(8'h96)) lut_n7259 (.I0(n7202), .I1(n7220), .I2(n7221), .O(n7259));
  LUT3 #(.INIT(8'hE8)) lut_n7260 (.I0(n7240), .I1(n7258), .I2(n7259), .O(n7260));
  LUT3 #(.INIT(8'h96)) lut_n7261 (.I0(n7140), .I1(n7178), .I2(n7179), .O(n7261));
  LUT3 #(.INIT(8'hE8)) lut_n7262 (.I0(n7222), .I1(n7260), .I2(n7261), .O(n7262));
  LUT3 #(.INIT(8'h96)) lut_n7263 (.I0(x2160), .I1(x2161), .I2(x2162), .O(n7263));
  LUT5 #(.INIT(32'h96696996)) lut_n7264 (.I0(x2151), .I1(x2152), .I2(x2153), .I3(n7252), .I4(n7253), .O(n7264));
  LUT5 #(.INIT(32'hFF969600)) lut_n7265 (.I0(x2157), .I1(x2158), .I2(x2159), .I3(n7263), .I4(n7264), .O(n7265));
  LUT3 #(.INIT(8'h96)) lut_n7266 (.I0(x2166), .I1(x2167), .I2(x2168), .O(n7266));
  LUT5 #(.INIT(32'h96696996)) lut_n7267 (.I0(x2157), .I1(x2158), .I2(x2159), .I3(n7263), .I4(n7264), .O(n7267));
  LUT5 #(.INIT(32'hFF969600)) lut_n7268 (.I0(x2163), .I1(x2164), .I2(x2165), .I3(n7266), .I4(n7267), .O(n7268));
  LUT3 #(.INIT(8'h96)) lut_n7269 (.I0(n7251), .I1(n7254), .I2(n7255), .O(n7269));
  LUT3 #(.INIT(8'hE8)) lut_n7270 (.I0(n7265), .I1(n7268), .I2(n7269), .O(n7270));
  LUT3 #(.INIT(8'h96)) lut_n7271 (.I0(x2172), .I1(x2173), .I2(x2174), .O(n7271));
  LUT5 #(.INIT(32'h96696996)) lut_n7272 (.I0(x2163), .I1(x2164), .I2(x2165), .I3(n7266), .I4(n7267), .O(n7272));
  LUT5 #(.INIT(32'hFF969600)) lut_n7273 (.I0(x2169), .I1(x2170), .I2(x2171), .I3(n7271), .I4(n7272), .O(n7273));
  LUT3 #(.INIT(8'h96)) lut_n7274 (.I0(x2178), .I1(x2179), .I2(x2180), .O(n7274));
  LUT5 #(.INIT(32'h96696996)) lut_n7275 (.I0(x2169), .I1(x2170), .I2(x2171), .I3(n7271), .I4(n7272), .O(n7275));
  LUT5 #(.INIT(32'hFF969600)) lut_n7276 (.I0(x2175), .I1(x2176), .I2(x2177), .I3(n7274), .I4(n7275), .O(n7276));
  LUT3 #(.INIT(8'h96)) lut_n7277 (.I0(n7265), .I1(n7268), .I2(n7269), .O(n7277));
  LUT3 #(.INIT(8'hE8)) lut_n7278 (.I0(n7273), .I1(n7276), .I2(n7277), .O(n7278));
  LUT3 #(.INIT(8'h96)) lut_n7279 (.I0(n7248), .I1(n7256), .I2(n7257), .O(n7279));
  LUT3 #(.INIT(8'hE8)) lut_n7280 (.I0(n7270), .I1(n7278), .I2(n7279), .O(n7280));
  LUT3 #(.INIT(8'h96)) lut_n7281 (.I0(x2184), .I1(x2185), .I2(x2186), .O(n7281));
  LUT5 #(.INIT(32'h96696996)) lut_n7282 (.I0(x2175), .I1(x2176), .I2(x2177), .I3(n7274), .I4(n7275), .O(n7282));
  LUT5 #(.INIT(32'hFF969600)) lut_n7283 (.I0(x2181), .I1(x2182), .I2(x2183), .I3(n7281), .I4(n7282), .O(n7283));
  LUT3 #(.INIT(8'h96)) lut_n7284 (.I0(x2190), .I1(x2191), .I2(x2192), .O(n7284));
  LUT5 #(.INIT(32'h96696996)) lut_n7285 (.I0(x2181), .I1(x2182), .I2(x2183), .I3(n7281), .I4(n7282), .O(n7285));
  LUT5 #(.INIT(32'hFF969600)) lut_n7286 (.I0(x2187), .I1(x2188), .I2(x2189), .I3(n7284), .I4(n7285), .O(n7286));
  LUT3 #(.INIT(8'h96)) lut_n7287 (.I0(n7273), .I1(n7276), .I2(n7277), .O(n7287));
  LUT3 #(.INIT(8'hE8)) lut_n7288 (.I0(n7283), .I1(n7286), .I2(n7287), .O(n7288));
  LUT3 #(.INIT(8'h96)) lut_n7289 (.I0(x2196), .I1(x2197), .I2(x2198), .O(n7289));
  LUT5 #(.INIT(32'h96696996)) lut_n7290 (.I0(x2187), .I1(x2188), .I2(x2189), .I3(n7284), .I4(n7285), .O(n7290));
  LUT5 #(.INIT(32'hFF969600)) lut_n7291 (.I0(x2193), .I1(x2194), .I2(x2195), .I3(n7289), .I4(n7290), .O(n7291));
  LUT3 #(.INIT(8'h96)) lut_n7292 (.I0(x2202), .I1(x2203), .I2(x2204), .O(n7292));
  LUT5 #(.INIT(32'h96696996)) lut_n7293 (.I0(x2193), .I1(x2194), .I2(x2195), .I3(n7289), .I4(n7290), .O(n7293));
  LUT5 #(.INIT(32'hFF969600)) lut_n7294 (.I0(x2199), .I1(x2200), .I2(x2201), .I3(n7292), .I4(n7293), .O(n7294));
  LUT3 #(.INIT(8'h96)) lut_n7295 (.I0(n7283), .I1(n7286), .I2(n7287), .O(n7295));
  LUT3 #(.INIT(8'hE8)) lut_n7296 (.I0(n7291), .I1(n7294), .I2(n7295), .O(n7296));
  LUT3 #(.INIT(8'h96)) lut_n7297 (.I0(n7270), .I1(n7278), .I2(n7279), .O(n7297));
  LUT3 #(.INIT(8'hE8)) lut_n7298 (.I0(n7288), .I1(n7296), .I2(n7297), .O(n7298));
  LUT3 #(.INIT(8'h96)) lut_n7299 (.I0(n7240), .I1(n7258), .I2(n7259), .O(n7299));
  LUT3 #(.INIT(8'hE8)) lut_n7300 (.I0(n7280), .I1(n7298), .I2(n7299), .O(n7300));
  LUT3 #(.INIT(8'h96)) lut_n7301 (.I0(x2208), .I1(x2209), .I2(x2210), .O(n7301));
  LUT5 #(.INIT(32'h96696996)) lut_n7302 (.I0(x2199), .I1(x2200), .I2(x2201), .I3(n7292), .I4(n7293), .O(n7302));
  LUT5 #(.INIT(32'hFF969600)) lut_n7303 (.I0(x2205), .I1(x2206), .I2(x2207), .I3(n7301), .I4(n7302), .O(n7303));
  LUT3 #(.INIT(8'h96)) lut_n7304 (.I0(x2214), .I1(x2215), .I2(x2216), .O(n7304));
  LUT5 #(.INIT(32'h96696996)) lut_n7305 (.I0(x2205), .I1(x2206), .I2(x2207), .I3(n7301), .I4(n7302), .O(n7305));
  LUT5 #(.INIT(32'hFF969600)) lut_n7306 (.I0(x2211), .I1(x2212), .I2(x2213), .I3(n7304), .I4(n7305), .O(n7306));
  LUT3 #(.INIT(8'h96)) lut_n7307 (.I0(n7291), .I1(n7294), .I2(n7295), .O(n7307));
  LUT3 #(.INIT(8'hE8)) lut_n7308 (.I0(n7303), .I1(n7306), .I2(n7307), .O(n7308));
  LUT3 #(.INIT(8'h96)) lut_n7309 (.I0(x2220), .I1(x2221), .I2(x2222), .O(n7309));
  LUT5 #(.INIT(32'h96696996)) lut_n7310 (.I0(x2211), .I1(x2212), .I2(x2213), .I3(n7304), .I4(n7305), .O(n7310));
  LUT5 #(.INIT(32'hFF969600)) lut_n7311 (.I0(x2217), .I1(x2218), .I2(x2219), .I3(n7309), .I4(n7310), .O(n7311));
  LUT3 #(.INIT(8'h96)) lut_n7312 (.I0(x2226), .I1(x2227), .I2(x2228), .O(n7312));
  LUT5 #(.INIT(32'h96696996)) lut_n7313 (.I0(x2217), .I1(x2218), .I2(x2219), .I3(n7309), .I4(n7310), .O(n7313));
  LUT5 #(.INIT(32'hFF969600)) lut_n7314 (.I0(x2223), .I1(x2224), .I2(x2225), .I3(n7312), .I4(n7313), .O(n7314));
  LUT3 #(.INIT(8'h96)) lut_n7315 (.I0(n7303), .I1(n7306), .I2(n7307), .O(n7315));
  LUT3 #(.INIT(8'hE8)) lut_n7316 (.I0(n7311), .I1(n7314), .I2(n7315), .O(n7316));
  LUT3 #(.INIT(8'h96)) lut_n7317 (.I0(n7288), .I1(n7296), .I2(n7297), .O(n7317));
  LUT3 #(.INIT(8'hE8)) lut_n7318 (.I0(n7308), .I1(n7316), .I2(n7317), .O(n7318));
  LUT3 #(.INIT(8'h96)) lut_n7319 (.I0(x2232), .I1(x2233), .I2(x2234), .O(n7319));
  LUT5 #(.INIT(32'h96696996)) lut_n7320 (.I0(x2223), .I1(x2224), .I2(x2225), .I3(n7312), .I4(n7313), .O(n7320));
  LUT5 #(.INIT(32'hFF969600)) lut_n7321 (.I0(x2229), .I1(x2230), .I2(x2231), .I3(n7319), .I4(n7320), .O(n7321));
  LUT3 #(.INIT(8'h96)) lut_n7322 (.I0(x2238), .I1(x2239), .I2(x2240), .O(n7322));
  LUT5 #(.INIT(32'h96696996)) lut_n7323 (.I0(x2229), .I1(x2230), .I2(x2231), .I3(n7319), .I4(n7320), .O(n7323));
  LUT5 #(.INIT(32'hFF969600)) lut_n7324 (.I0(x2235), .I1(x2236), .I2(x2237), .I3(n7322), .I4(n7323), .O(n7324));
  LUT3 #(.INIT(8'h96)) lut_n7325 (.I0(n7311), .I1(n7314), .I2(n7315), .O(n7325));
  LUT3 #(.INIT(8'hE8)) lut_n7326 (.I0(n7321), .I1(n7324), .I2(n7325), .O(n7326));
  LUT3 #(.INIT(8'h96)) lut_n7327 (.I0(x2244), .I1(x2245), .I2(x2246), .O(n7327));
  LUT5 #(.INIT(32'h96696996)) lut_n7328 (.I0(x2235), .I1(x2236), .I2(x2237), .I3(n7322), .I4(n7323), .O(n7328));
  LUT5 #(.INIT(32'hFF969600)) lut_n7329 (.I0(x2241), .I1(x2242), .I2(x2243), .I3(n7327), .I4(n7328), .O(n7329));
  LUT3 #(.INIT(8'h96)) lut_n7330 (.I0(x2250), .I1(x2251), .I2(x2252), .O(n7330));
  LUT5 #(.INIT(32'h96696996)) lut_n7331 (.I0(x2241), .I1(x2242), .I2(x2243), .I3(n7327), .I4(n7328), .O(n7331));
  LUT5 #(.INIT(32'hFF969600)) lut_n7332 (.I0(x2247), .I1(x2248), .I2(x2249), .I3(n7330), .I4(n7331), .O(n7332));
  LUT3 #(.INIT(8'h96)) lut_n7333 (.I0(n7321), .I1(n7324), .I2(n7325), .O(n7333));
  LUT3 #(.INIT(8'hE8)) lut_n7334 (.I0(n7329), .I1(n7332), .I2(n7333), .O(n7334));
  LUT3 #(.INIT(8'h96)) lut_n7335 (.I0(n7308), .I1(n7316), .I2(n7317), .O(n7335));
  LUT3 #(.INIT(8'hE8)) lut_n7336 (.I0(n7326), .I1(n7334), .I2(n7335), .O(n7336));
  LUT3 #(.INIT(8'h96)) lut_n7337 (.I0(n7280), .I1(n7298), .I2(n7299), .O(n7337));
  LUT3 #(.INIT(8'hE8)) lut_n7338 (.I0(n7318), .I1(n7336), .I2(n7337), .O(n7338));
  LUT3 #(.INIT(8'h96)) lut_n7339 (.I0(n7222), .I1(n7260), .I2(n7261), .O(n7339));
  LUT3 #(.INIT(8'hE8)) lut_n7340 (.I0(n7300), .I1(n7338), .I2(n7339), .O(n7340));
  LUT3 #(.INIT(8'h96)) lut_n7341 (.I0(n7102), .I1(n7180), .I2(n7181), .O(n7341));
  LUT3 #(.INIT(8'hE8)) lut_n7342 (.I0(n7262), .I1(n7340), .I2(n7341), .O(n7342));
  LUT3 #(.INIT(8'h96)) lut_n7343 (.I0(x2256), .I1(x2257), .I2(x2258), .O(n7343));
  LUT5 #(.INIT(32'h96696996)) lut_n7344 (.I0(x2247), .I1(x2248), .I2(x2249), .I3(n7330), .I4(n7331), .O(n7344));
  LUT5 #(.INIT(32'hFF969600)) lut_n7345 (.I0(x2253), .I1(x2254), .I2(x2255), .I3(n7343), .I4(n7344), .O(n7345));
  LUT3 #(.INIT(8'h96)) lut_n7346 (.I0(x2262), .I1(x2263), .I2(x2264), .O(n7346));
  LUT5 #(.INIT(32'h96696996)) lut_n7347 (.I0(x2253), .I1(x2254), .I2(x2255), .I3(n7343), .I4(n7344), .O(n7347));
  LUT5 #(.INIT(32'hFF969600)) lut_n7348 (.I0(x2259), .I1(x2260), .I2(x2261), .I3(n7346), .I4(n7347), .O(n7348));
  LUT3 #(.INIT(8'h96)) lut_n7349 (.I0(n7329), .I1(n7332), .I2(n7333), .O(n7349));
  LUT3 #(.INIT(8'hE8)) lut_n7350 (.I0(n7345), .I1(n7348), .I2(n7349), .O(n7350));
  LUT3 #(.INIT(8'h96)) lut_n7351 (.I0(x2268), .I1(x2269), .I2(x2270), .O(n7351));
  LUT5 #(.INIT(32'h96696996)) lut_n7352 (.I0(x2259), .I1(x2260), .I2(x2261), .I3(n7346), .I4(n7347), .O(n7352));
  LUT5 #(.INIT(32'hFF969600)) lut_n7353 (.I0(x2265), .I1(x2266), .I2(x2267), .I3(n7351), .I4(n7352), .O(n7353));
  LUT3 #(.INIT(8'h96)) lut_n7354 (.I0(x2274), .I1(x2275), .I2(x2276), .O(n7354));
  LUT5 #(.INIT(32'h96696996)) lut_n7355 (.I0(x2265), .I1(x2266), .I2(x2267), .I3(n7351), .I4(n7352), .O(n7355));
  LUT5 #(.INIT(32'hFF969600)) lut_n7356 (.I0(x2271), .I1(x2272), .I2(x2273), .I3(n7354), .I4(n7355), .O(n7356));
  LUT3 #(.INIT(8'h96)) lut_n7357 (.I0(n7345), .I1(n7348), .I2(n7349), .O(n7357));
  LUT3 #(.INIT(8'hE8)) lut_n7358 (.I0(n7353), .I1(n7356), .I2(n7357), .O(n7358));
  LUT3 #(.INIT(8'h96)) lut_n7359 (.I0(n7326), .I1(n7334), .I2(n7335), .O(n7359));
  LUT3 #(.INIT(8'hE8)) lut_n7360 (.I0(n7350), .I1(n7358), .I2(n7359), .O(n7360));
  LUT3 #(.INIT(8'h96)) lut_n7361 (.I0(x2280), .I1(x2281), .I2(x2282), .O(n7361));
  LUT5 #(.INIT(32'h96696996)) lut_n7362 (.I0(x2271), .I1(x2272), .I2(x2273), .I3(n7354), .I4(n7355), .O(n7362));
  LUT5 #(.INIT(32'hFF969600)) lut_n7363 (.I0(x2277), .I1(x2278), .I2(x2279), .I3(n7361), .I4(n7362), .O(n7363));
  LUT3 #(.INIT(8'h96)) lut_n7364 (.I0(x2286), .I1(x2287), .I2(x2288), .O(n7364));
  LUT5 #(.INIT(32'h96696996)) lut_n7365 (.I0(x2277), .I1(x2278), .I2(x2279), .I3(n7361), .I4(n7362), .O(n7365));
  LUT5 #(.INIT(32'hFF969600)) lut_n7366 (.I0(x2283), .I1(x2284), .I2(x2285), .I3(n7364), .I4(n7365), .O(n7366));
  LUT3 #(.INIT(8'h96)) lut_n7367 (.I0(n7353), .I1(n7356), .I2(n7357), .O(n7367));
  LUT3 #(.INIT(8'hE8)) lut_n7368 (.I0(n7363), .I1(n7366), .I2(n7367), .O(n7368));
  LUT3 #(.INIT(8'h96)) lut_n7369 (.I0(x2292), .I1(x2293), .I2(x2294), .O(n7369));
  LUT5 #(.INIT(32'h96696996)) lut_n7370 (.I0(x2283), .I1(x2284), .I2(x2285), .I3(n7364), .I4(n7365), .O(n7370));
  LUT5 #(.INIT(32'hFF969600)) lut_n7371 (.I0(x2289), .I1(x2290), .I2(x2291), .I3(n7369), .I4(n7370), .O(n7371));
  LUT3 #(.INIT(8'h96)) lut_n7372 (.I0(x2298), .I1(x2299), .I2(x2300), .O(n7372));
  LUT5 #(.INIT(32'h96696996)) lut_n7373 (.I0(x2289), .I1(x2290), .I2(x2291), .I3(n7369), .I4(n7370), .O(n7373));
  LUT5 #(.INIT(32'hFF969600)) lut_n7374 (.I0(x2295), .I1(x2296), .I2(x2297), .I3(n7372), .I4(n7373), .O(n7374));
  LUT3 #(.INIT(8'h96)) lut_n7375 (.I0(n7363), .I1(n7366), .I2(n7367), .O(n7375));
  LUT3 #(.INIT(8'hE8)) lut_n7376 (.I0(n7371), .I1(n7374), .I2(n7375), .O(n7376));
  LUT3 #(.INIT(8'h96)) lut_n7377 (.I0(n7350), .I1(n7358), .I2(n7359), .O(n7377));
  LUT3 #(.INIT(8'hE8)) lut_n7378 (.I0(n7368), .I1(n7376), .I2(n7377), .O(n7378));
  LUT3 #(.INIT(8'h96)) lut_n7379 (.I0(n7318), .I1(n7336), .I2(n7337), .O(n7379));
  LUT3 #(.INIT(8'hE8)) lut_n7380 (.I0(n7360), .I1(n7378), .I2(n7379), .O(n7380));
  LUT3 #(.INIT(8'h96)) lut_n7381 (.I0(x2304), .I1(x2305), .I2(x2306), .O(n7381));
  LUT5 #(.INIT(32'h96696996)) lut_n7382 (.I0(x2295), .I1(x2296), .I2(x2297), .I3(n7372), .I4(n7373), .O(n7382));
  LUT5 #(.INIT(32'hFF969600)) lut_n7383 (.I0(x2301), .I1(x2302), .I2(x2303), .I3(n7381), .I4(n7382), .O(n7383));
  LUT3 #(.INIT(8'h96)) lut_n7384 (.I0(x2310), .I1(x2311), .I2(x2312), .O(n7384));
  LUT5 #(.INIT(32'h96696996)) lut_n7385 (.I0(x2301), .I1(x2302), .I2(x2303), .I3(n7381), .I4(n7382), .O(n7385));
  LUT5 #(.INIT(32'hFF969600)) lut_n7386 (.I0(x2307), .I1(x2308), .I2(x2309), .I3(n7384), .I4(n7385), .O(n7386));
  LUT3 #(.INIT(8'h96)) lut_n7387 (.I0(n7371), .I1(n7374), .I2(n7375), .O(n7387));
  LUT3 #(.INIT(8'hE8)) lut_n7388 (.I0(n7383), .I1(n7386), .I2(n7387), .O(n7388));
  LUT3 #(.INIT(8'h96)) lut_n7389 (.I0(x2316), .I1(x2317), .I2(x2318), .O(n7389));
  LUT5 #(.INIT(32'h96696996)) lut_n7390 (.I0(x2307), .I1(x2308), .I2(x2309), .I3(n7384), .I4(n7385), .O(n7390));
  LUT5 #(.INIT(32'hFF969600)) lut_n7391 (.I0(x2313), .I1(x2314), .I2(x2315), .I3(n7389), .I4(n7390), .O(n7391));
  LUT3 #(.INIT(8'h96)) lut_n7392 (.I0(x2322), .I1(x2323), .I2(x2324), .O(n7392));
  LUT5 #(.INIT(32'h96696996)) lut_n7393 (.I0(x2313), .I1(x2314), .I2(x2315), .I3(n7389), .I4(n7390), .O(n7393));
  LUT5 #(.INIT(32'hFF969600)) lut_n7394 (.I0(x2319), .I1(x2320), .I2(x2321), .I3(n7392), .I4(n7393), .O(n7394));
  LUT3 #(.INIT(8'h96)) lut_n7395 (.I0(n7383), .I1(n7386), .I2(n7387), .O(n7395));
  LUT3 #(.INIT(8'hE8)) lut_n7396 (.I0(n7391), .I1(n7394), .I2(n7395), .O(n7396));
  LUT3 #(.INIT(8'h96)) lut_n7397 (.I0(n7368), .I1(n7376), .I2(n7377), .O(n7397));
  LUT3 #(.INIT(8'hE8)) lut_n7398 (.I0(n7388), .I1(n7396), .I2(n7397), .O(n7398));
  LUT3 #(.INIT(8'h96)) lut_n7399 (.I0(x2328), .I1(x2329), .I2(x2330), .O(n7399));
  LUT5 #(.INIT(32'h96696996)) lut_n7400 (.I0(x2319), .I1(x2320), .I2(x2321), .I3(n7392), .I4(n7393), .O(n7400));
  LUT5 #(.INIT(32'hFF969600)) lut_n7401 (.I0(x2325), .I1(x2326), .I2(x2327), .I3(n7399), .I4(n7400), .O(n7401));
  LUT3 #(.INIT(8'h96)) lut_n7402 (.I0(x2334), .I1(x2335), .I2(x2336), .O(n7402));
  LUT5 #(.INIT(32'h96696996)) lut_n7403 (.I0(x2325), .I1(x2326), .I2(x2327), .I3(n7399), .I4(n7400), .O(n7403));
  LUT5 #(.INIT(32'hFF969600)) lut_n7404 (.I0(x2331), .I1(x2332), .I2(x2333), .I3(n7402), .I4(n7403), .O(n7404));
  LUT3 #(.INIT(8'h96)) lut_n7405 (.I0(n7391), .I1(n7394), .I2(n7395), .O(n7405));
  LUT3 #(.INIT(8'hE8)) lut_n7406 (.I0(n7401), .I1(n7404), .I2(n7405), .O(n7406));
  LUT3 #(.INIT(8'h96)) lut_n7407 (.I0(x2340), .I1(x2341), .I2(x2342), .O(n7407));
  LUT5 #(.INIT(32'h96696996)) lut_n7408 (.I0(x2331), .I1(x2332), .I2(x2333), .I3(n7402), .I4(n7403), .O(n7408));
  LUT5 #(.INIT(32'hFF969600)) lut_n7409 (.I0(x2337), .I1(x2338), .I2(x2339), .I3(n7407), .I4(n7408), .O(n7409));
  LUT3 #(.INIT(8'h96)) lut_n7410 (.I0(x2346), .I1(x2347), .I2(x2348), .O(n7410));
  LUT5 #(.INIT(32'h96696996)) lut_n7411 (.I0(x2337), .I1(x2338), .I2(x2339), .I3(n7407), .I4(n7408), .O(n7411));
  LUT5 #(.INIT(32'hFF969600)) lut_n7412 (.I0(x2343), .I1(x2344), .I2(x2345), .I3(n7410), .I4(n7411), .O(n7412));
  LUT3 #(.INIT(8'h96)) lut_n7413 (.I0(n7401), .I1(n7404), .I2(n7405), .O(n7413));
  LUT3 #(.INIT(8'hE8)) lut_n7414 (.I0(n7409), .I1(n7412), .I2(n7413), .O(n7414));
  LUT3 #(.INIT(8'h96)) lut_n7415 (.I0(n7388), .I1(n7396), .I2(n7397), .O(n7415));
  LUT3 #(.INIT(8'hE8)) lut_n7416 (.I0(n7406), .I1(n7414), .I2(n7415), .O(n7416));
  LUT3 #(.INIT(8'h96)) lut_n7417 (.I0(n7360), .I1(n7378), .I2(n7379), .O(n7417));
  LUT3 #(.INIT(8'hE8)) lut_n7418 (.I0(n7398), .I1(n7416), .I2(n7417), .O(n7418));
  LUT3 #(.INIT(8'h96)) lut_n7419 (.I0(n7300), .I1(n7338), .I2(n7339), .O(n7419));
  LUT3 #(.INIT(8'hE8)) lut_n7420 (.I0(n7380), .I1(n7418), .I2(n7419), .O(n7420));
  LUT3 #(.INIT(8'h96)) lut_n7421 (.I0(x2352), .I1(x2353), .I2(x2354), .O(n7421));
  LUT5 #(.INIT(32'h96696996)) lut_n7422 (.I0(x2343), .I1(x2344), .I2(x2345), .I3(n7410), .I4(n7411), .O(n7422));
  LUT5 #(.INIT(32'hFF969600)) lut_n7423 (.I0(x2349), .I1(x2350), .I2(x2351), .I3(n7421), .I4(n7422), .O(n7423));
  LUT3 #(.INIT(8'h96)) lut_n7424 (.I0(x2358), .I1(x2359), .I2(x2360), .O(n7424));
  LUT5 #(.INIT(32'h96696996)) lut_n7425 (.I0(x2349), .I1(x2350), .I2(x2351), .I3(n7421), .I4(n7422), .O(n7425));
  LUT5 #(.INIT(32'hFF969600)) lut_n7426 (.I0(x2355), .I1(x2356), .I2(x2357), .I3(n7424), .I4(n7425), .O(n7426));
  LUT3 #(.INIT(8'h96)) lut_n7427 (.I0(n7409), .I1(n7412), .I2(n7413), .O(n7427));
  LUT3 #(.INIT(8'hE8)) lut_n7428 (.I0(n7423), .I1(n7426), .I2(n7427), .O(n7428));
  LUT3 #(.INIT(8'h96)) lut_n7429 (.I0(x2364), .I1(x2365), .I2(x2366), .O(n7429));
  LUT5 #(.INIT(32'h96696996)) lut_n7430 (.I0(x2355), .I1(x2356), .I2(x2357), .I3(n7424), .I4(n7425), .O(n7430));
  LUT5 #(.INIT(32'hFF969600)) lut_n7431 (.I0(x2361), .I1(x2362), .I2(x2363), .I3(n7429), .I4(n7430), .O(n7431));
  LUT3 #(.INIT(8'h96)) lut_n7432 (.I0(x2370), .I1(x2371), .I2(x2372), .O(n7432));
  LUT5 #(.INIT(32'h96696996)) lut_n7433 (.I0(x2361), .I1(x2362), .I2(x2363), .I3(n7429), .I4(n7430), .O(n7433));
  LUT5 #(.INIT(32'hFF969600)) lut_n7434 (.I0(x2367), .I1(x2368), .I2(x2369), .I3(n7432), .I4(n7433), .O(n7434));
  LUT3 #(.INIT(8'h96)) lut_n7435 (.I0(n7423), .I1(n7426), .I2(n7427), .O(n7435));
  LUT3 #(.INIT(8'hE8)) lut_n7436 (.I0(n7431), .I1(n7434), .I2(n7435), .O(n7436));
  LUT3 #(.INIT(8'h96)) lut_n7437 (.I0(n7406), .I1(n7414), .I2(n7415), .O(n7437));
  LUT3 #(.INIT(8'hE8)) lut_n7438 (.I0(n7428), .I1(n7436), .I2(n7437), .O(n7438));
  LUT3 #(.INIT(8'h96)) lut_n7439 (.I0(x2376), .I1(x2377), .I2(x2378), .O(n7439));
  LUT5 #(.INIT(32'h96696996)) lut_n7440 (.I0(x2367), .I1(x2368), .I2(x2369), .I3(n7432), .I4(n7433), .O(n7440));
  LUT5 #(.INIT(32'hFF969600)) lut_n7441 (.I0(x2373), .I1(x2374), .I2(x2375), .I3(n7439), .I4(n7440), .O(n7441));
  LUT3 #(.INIT(8'h96)) lut_n7442 (.I0(x2382), .I1(x2383), .I2(x2384), .O(n7442));
  LUT5 #(.INIT(32'h96696996)) lut_n7443 (.I0(x2373), .I1(x2374), .I2(x2375), .I3(n7439), .I4(n7440), .O(n7443));
  LUT5 #(.INIT(32'hFF969600)) lut_n7444 (.I0(x2379), .I1(x2380), .I2(x2381), .I3(n7442), .I4(n7443), .O(n7444));
  LUT3 #(.INIT(8'h96)) lut_n7445 (.I0(n7431), .I1(n7434), .I2(n7435), .O(n7445));
  LUT3 #(.INIT(8'hE8)) lut_n7446 (.I0(n7441), .I1(n7444), .I2(n7445), .O(n7446));
  LUT3 #(.INIT(8'h96)) lut_n7447 (.I0(x2388), .I1(x2389), .I2(x2390), .O(n7447));
  LUT5 #(.INIT(32'h96696996)) lut_n7448 (.I0(x2379), .I1(x2380), .I2(x2381), .I3(n7442), .I4(n7443), .O(n7448));
  LUT5 #(.INIT(32'hFF969600)) lut_n7449 (.I0(x2385), .I1(x2386), .I2(x2387), .I3(n7447), .I4(n7448), .O(n7449));
  LUT3 #(.INIT(8'h96)) lut_n7450 (.I0(x2394), .I1(x2395), .I2(x2396), .O(n7450));
  LUT5 #(.INIT(32'h96696996)) lut_n7451 (.I0(x2385), .I1(x2386), .I2(x2387), .I3(n7447), .I4(n7448), .O(n7451));
  LUT5 #(.INIT(32'hFF969600)) lut_n7452 (.I0(x2391), .I1(x2392), .I2(x2393), .I3(n7450), .I4(n7451), .O(n7452));
  LUT3 #(.INIT(8'h96)) lut_n7453 (.I0(n7441), .I1(n7444), .I2(n7445), .O(n7453));
  LUT3 #(.INIT(8'hE8)) lut_n7454 (.I0(n7449), .I1(n7452), .I2(n7453), .O(n7454));
  LUT3 #(.INIT(8'h96)) lut_n7455 (.I0(n7428), .I1(n7436), .I2(n7437), .O(n7455));
  LUT3 #(.INIT(8'hE8)) lut_n7456 (.I0(n7446), .I1(n7454), .I2(n7455), .O(n7456));
  LUT3 #(.INIT(8'h96)) lut_n7457 (.I0(n7398), .I1(n7416), .I2(n7417), .O(n7457));
  LUT3 #(.INIT(8'hE8)) lut_n7458 (.I0(n7438), .I1(n7456), .I2(n7457), .O(n7458));
  LUT3 #(.INIT(8'h96)) lut_n7459 (.I0(x2400), .I1(x2401), .I2(x2402), .O(n7459));
  LUT5 #(.INIT(32'h96696996)) lut_n7460 (.I0(x2391), .I1(x2392), .I2(x2393), .I3(n7450), .I4(n7451), .O(n7460));
  LUT5 #(.INIT(32'hFF969600)) lut_n7461 (.I0(x2397), .I1(x2398), .I2(x2399), .I3(n7459), .I4(n7460), .O(n7461));
  LUT3 #(.INIT(8'h96)) lut_n7462 (.I0(x2406), .I1(x2407), .I2(x2408), .O(n7462));
  LUT5 #(.INIT(32'h96696996)) lut_n7463 (.I0(x2397), .I1(x2398), .I2(x2399), .I3(n7459), .I4(n7460), .O(n7463));
  LUT5 #(.INIT(32'hFF969600)) lut_n7464 (.I0(x2403), .I1(x2404), .I2(x2405), .I3(n7462), .I4(n7463), .O(n7464));
  LUT3 #(.INIT(8'h96)) lut_n7465 (.I0(n7449), .I1(n7452), .I2(n7453), .O(n7465));
  LUT3 #(.INIT(8'hE8)) lut_n7466 (.I0(n7461), .I1(n7464), .I2(n7465), .O(n7466));
  LUT3 #(.INIT(8'h96)) lut_n7467 (.I0(x2412), .I1(x2413), .I2(x2414), .O(n7467));
  LUT5 #(.INIT(32'h96696996)) lut_n7468 (.I0(x2403), .I1(x2404), .I2(x2405), .I3(n7462), .I4(n7463), .O(n7468));
  LUT5 #(.INIT(32'hFF969600)) lut_n7469 (.I0(x2409), .I1(x2410), .I2(x2411), .I3(n7467), .I4(n7468), .O(n7469));
  LUT3 #(.INIT(8'h96)) lut_n7470 (.I0(x2418), .I1(x2419), .I2(x2420), .O(n7470));
  LUT5 #(.INIT(32'h96696996)) lut_n7471 (.I0(x2409), .I1(x2410), .I2(x2411), .I3(n7467), .I4(n7468), .O(n7471));
  LUT5 #(.INIT(32'hFF969600)) lut_n7472 (.I0(x2415), .I1(x2416), .I2(x2417), .I3(n7470), .I4(n7471), .O(n7472));
  LUT3 #(.INIT(8'h96)) lut_n7473 (.I0(n7461), .I1(n7464), .I2(n7465), .O(n7473));
  LUT3 #(.INIT(8'hE8)) lut_n7474 (.I0(n7469), .I1(n7472), .I2(n7473), .O(n7474));
  LUT3 #(.INIT(8'h96)) lut_n7475 (.I0(n7446), .I1(n7454), .I2(n7455), .O(n7475));
  LUT3 #(.INIT(8'hE8)) lut_n7476 (.I0(n7466), .I1(n7474), .I2(n7475), .O(n7476));
  LUT3 #(.INIT(8'h96)) lut_n7477 (.I0(x2424), .I1(x2425), .I2(x2426), .O(n7477));
  LUT5 #(.INIT(32'h96696996)) lut_n7478 (.I0(x2415), .I1(x2416), .I2(x2417), .I3(n7470), .I4(n7471), .O(n7478));
  LUT5 #(.INIT(32'hFF969600)) lut_n7479 (.I0(x2421), .I1(x2422), .I2(x2423), .I3(n7477), .I4(n7478), .O(n7479));
  LUT3 #(.INIT(8'h96)) lut_n7480 (.I0(x2430), .I1(x2431), .I2(x2432), .O(n7480));
  LUT5 #(.INIT(32'h96696996)) lut_n7481 (.I0(x2421), .I1(x2422), .I2(x2423), .I3(n7477), .I4(n7478), .O(n7481));
  LUT5 #(.INIT(32'hFF969600)) lut_n7482 (.I0(x2427), .I1(x2428), .I2(x2429), .I3(n7480), .I4(n7481), .O(n7482));
  LUT3 #(.INIT(8'h96)) lut_n7483 (.I0(n7469), .I1(n7472), .I2(n7473), .O(n7483));
  LUT3 #(.INIT(8'hE8)) lut_n7484 (.I0(n7479), .I1(n7482), .I2(n7483), .O(n7484));
  LUT3 #(.INIT(8'h96)) lut_n7485 (.I0(x2436), .I1(x2437), .I2(x2438), .O(n7485));
  LUT5 #(.INIT(32'h96696996)) lut_n7486 (.I0(x2427), .I1(x2428), .I2(x2429), .I3(n7480), .I4(n7481), .O(n7486));
  LUT5 #(.INIT(32'hFF969600)) lut_n7487 (.I0(x2433), .I1(x2434), .I2(x2435), .I3(n7485), .I4(n7486), .O(n7487));
  LUT3 #(.INIT(8'h96)) lut_n7488 (.I0(x2442), .I1(x2443), .I2(x2444), .O(n7488));
  LUT5 #(.INIT(32'h96696996)) lut_n7489 (.I0(x2433), .I1(x2434), .I2(x2435), .I3(n7485), .I4(n7486), .O(n7489));
  LUT5 #(.INIT(32'hFF969600)) lut_n7490 (.I0(x2439), .I1(x2440), .I2(x2441), .I3(n7488), .I4(n7489), .O(n7490));
  LUT3 #(.INIT(8'h96)) lut_n7491 (.I0(n7479), .I1(n7482), .I2(n7483), .O(n7491));
  LUT3 #(.INIT(8'hE8)) lut_n7492 (.I0(n7487), .I1(n7490), .I2(n7491), .O(n7492));
  LUT3 #(.INIT(8'h96)) lut_n7493 (.I0(n7466), .I1(n7474), .I2(n7475), .O(n7493));
  LUT3 #(.INIT(8'hE8)) lut_n7494 (.I0(n7484), .I1(n7492), .I2(n7493), .O(n7494));
  LUT3 #(.INIT(8'h96)) lut_n7495 (.I0(n7438), .I1(n7456), .I2(n7457), .O(n7495));
  LUT3 #(.INIT(8'hE8)) lut_n7496 (.I0(n7476), .I1(n7494), .I2(n7495), .O(n7496));
  LUT3 #(.INIT(8'h96)) lut_n7497 (.I0(n7380), .I1(n7418), .I2(n7419), .O(n7497));
  LUT3 #(.INIT(8'hE8)) lut_n7498 (.I0(n7458), .I1(n7496), .I2(n7497), .O(n7498));
  LUT3 #(.INIT(8'h96)) lut_n7499 (.I0(n7262), .I1(n7340), .I2(n7341), .O(n7499));
  LUT3 #(.INIT(8'hE8)) lut_n7500 (.I0(n7420), .I1(n7498), .I2(n7499), .O(n7500));
  LUT3 #(.INIT(8'h96)) lut_n7501 (.I0(n7024), .I1(n7182), .I2(n7183), .O(n7501));
  LUT3 #(.INIT(8'hE8)) lut_n7502 (.I0(n7342), .I1(n7500), .I2(n7501), .O(n7502));
  LUT3 #(.INIT(8'h96)) lut_n7503 (.I0(n6544), .I1(n6862), .I2(n6863), .O(n7503));
  LUT3 #(.INIT(8'hE8)) lut_n7504 (.I0(n7184), .I1(n7502), .I2(n7503), .O(n7504));
  LUT3 #(.INIT(8'h96)) lut_n7505 (.I0(x2448), .I1(x2449), .I2(x2450), .O(n7505));
  LUT5 #(.INIT(32'h96696996)) lut_n7506 (.I0(x2439), .I1(x2440), .I2(x2441), .I3(n7488), .I4(n7489), .O(n7506));
  LUT5 #(.INIT(32'hFF969600)) lut_n7507 (.I0(x2445), .I1(x2446), .I2(x2447), .I3(n7505), .I4(n7506), .O(n7507));
  LUT3 #(.INIT(8'h96)) lut_n7508 (.I0(x2454), .I1(x2455), .I2(x2456), .O(n7508));
  LUT5 #(.INIT(32'h96696996)) lut_n7509 (.I0(x2445), .I1(x2446), .I2(x2447), .I3(n7505), .I4(n7506), .O(n7509));
  LUT5 #(.INIT(32'hFF969600)) lut_n7510 (.I0(x2451), .I1(x2452), .I2(x2453), .I3(n7508), .I4(n7509), .O(n7510));
  LUT3 #(.INIT(8'h96)) lut_n7511 (.I0(n7487), .I1(n7490), .I2(n7491), .O(n7511));
  LUT3 #(.INIT(8'hE8)) lut_n7512 (.I0(n7507), .I1(n7510), .I2(n7511), .O(n7512));
  LUT3 #(.INIT(8'h96)) lut_n7513 (.I0(x2460), .I1(x2461), .I2(x2462), .O(n7513));
  LUT5 #(.INIT(32'h96696996)) lut_n7514 (.I0(x2451), .I1(x2452), .I2(x2453), .I3(n7508), .I4(n7509), .O(n7514));
  LUT5 #(.INIT(32'hFF969600)) lut_n7515 (.I0(x2457), .I1(x2458), .I2(x2459), .I3(n7513), .I4(n7514), .O(n7515));
  LUT3 #(.INIT(8'h96)) lut_n7516 (.I0(x2466), .I1(x2467), .I2(x2468), .O(n7516));
  LUT5 #(.INIT(32'h96696996)) lut_n7517 (.I0(x2457), .I1(x2458), .I2(x2459), .I3(n7513), .I4(n7514), .O(n7517));
  LUT5 #(.INIT(32'hFF969600)) lut_n7518 (.I0(x2463), .I1(x2464), .I2(x2465), .I3(n7516), .I4(n7517), .O(n7518));
  LUT3 #(.INIT(8'h96)) lut_n7519 (.I0(n7507), .I1(n7510), .I2(n7511), .O(n7519));
  LUT3 #(.INIT(8'hE8)) lut_n7520 (.I0(n7515), .I1(n7518), .I2(n7519), .O(n7520));
  LUT3 #(.INIT(8'h96)) lut_n7521 (.I0(n7484), .I1(n7492), .I2(n7493), .O(n7521));
  LUT3 #(.INIT(8'hE8)) lut_n7522 (.I0(n7512), .I1(n7520), .I2(n7521), .O(n7522));
  LUT3 #(.INIT(8'h96)) lut_n7523 (.I0(x2472), .I1(x2473), .I2(x2474), .O(n7523));
  LUT5 #(.INIT(32'h96696996)) lut_n7524 (.I0(x2463), .I1(x2464), .I2(x2465), .I3(n7516), .I4(n7517), .O(n7524));
  LUT5 #(.INIT(32'hFF969600)) lut_n7525 (.I0(x2469), .I1(x2470), .I2(x2471), .I3(n7523), .I4(n7524), .O(n7525));
  LUT3 #(.INIT(8'h96)) lut_n7526 (.I0(x2478), .I1(x2479), .I2(x2480), .O(n7526));
  LUT5 #(.INIT(32'h96696996)) lut_n7527 (.I0(x2469), .I1(x2470), .I2(x2471), .I3(n7523), .I4(n7524), .O(n7527));
  LUT5 #(.INIT(32'hFF969600)) lut_n7528 (.I0(x2475), .I1(x2476), .I2(x2477), .I3(n7526), .I4(n7527), .O(n7528));
  LUT3 #(.INIT(8'h96)) lut_n7529 (.I0(n7515), .I1(n7518), .I2(n7519), .O(n7529));
  LUT3 #(.INIT(8'hE8)) lut_n7530 (.I0(n7525), .I1(n7528), .I2(n7529), .O(n7530));
  LUT3 #(.INIT(8'h96)) lut_n7531 (.I0(x2484), .I1(x2485), .I2(x2486), .O(n7531));
  LUT5 #(.INIT(32'h96696996)) lut_n7532 (.I0(x2475), .I1(x2476), .I2(x2477), .I3(n7526), .I4(n7527), .O(n7532));
  LUT5 #(.INIT(32'hFF969600)) lut_n7533 (.I0(x2481), .I1(x2482), .I2(x2483), .I3(n7531), .I4(n7532), .O(n7533));
  LUT3 #(.INIT(8'h96)) lut_n7534 (.I0(x2490), .I1(x2491), .I2(x2492), .O(n7534));
  LUT5 #(.INIT(32'h96696996)) lut_n7535 (.I0(x2481), .I1(x2482), .I2(x2483), .I3(n7531), .I4(n7532), .O(n7535));
  LUT5 #(.INIT(32'hFF969600)) lut_n7536 (.I0(x2487), .I1(x2488), .I2(x2489), .I3(n7534), .I4(n7535), .O(n7536));
  LUT3 #(.INIT(8'h96)) lut_n7537 (.I0(n7525), .I1(n7528), .I2(n7529), .O(n7537));
  LUT3 #(.INIT(8'hE8)) lut_n7538 (.I0(n7533), .I1(n7536), .I2(n7537), .O(n7538));
  LUT3 #(.INIT(8'h96)) lut_n7539 (.I0(n7512), .I1(n7520), .I2(n7521), .O(n7539));
  LUT3 #(.INIT(8'hE8)) lut_n7540 (.I0(n7530), .I1(n7538), .I2(n7539), .O(n7540));
  LUT3 #(.INIT(8'h96)) lut_n7541 (.I0(n7476), .I1(n7494), .I2(n7495), .O(n7541));
  LUT3 #(.INIT(8'hE8)) lut_n7542 (.I0(n7522), .I1(n7540), .I2(n7541), .O(n7542));
  LUT3 #(.INIT(8'h96)) lut_n7543 (.I0(x2496), .I1(x2497), .I2(x2498), .O(n7543));
  LUT5 #(.INIT(32'h96696996)) lut_n7544 (.I0(x2487), .I1(x2488), .I2(x2489), .I3(n7534), .I4(n7535), .O(n7544));
  LUT5 #(.INIT(32'hFF969600)) lut_n7545 (.I0(x2493), .I1(x2494), .I2(x2495), .I3(n7543), .I4(n7544), .O(n7545));
  LUT3 #(.INIT(8'h96)) lut_n7546 (.I0(x2502), .I1(x2503), .I2(x2504), .O(n7546));
  LUT5 #(.INIT(32'h96696996)) lut_n7547 (.I0(x2493), .I1(x2494), .I2(x2495), .I3(n7543), .I4(n7544), .O(n7547));
  LUT5 #(.INIT(32'hFF969600)) lut_n7548 (.I0(x2499), .I1(x2500), .I2(x2501), .I3(n7546), .I4(n7547), .O(n7548));
  LUT3 #(.INIT(8'h96)) lut_n7549 (.I0(n7533), .I1(n7536), .I2(n7537), .O(n7549));
  LUT3 #(.INIT(8'hE8)) lut_n7550 (.I0(n7545), .I1(n7548), .I2(n7549), .O(n7550));
  LUT3 #(.INIT(8'h96)) lut_n7551 (.I0(x2508), .I1(x2509), .I2(x2510), .O(n7551));
  LUT5 #(.INIT(32'h96696996)) lut_n7552 (.I0(x2499), .I1(x2500), .I2(x2501), .I3(n7546), .I4(n7547), .O(n7552));
  LUT5 #(.INIT(32'hFF969600)) lut_n7553 (.I0(x2505), .I1(x2506), .I2(x2507), .I3(n7551), .I4(n7552), .O(n7553));
  LUT3 #(.INIT(8'h96)) lut_n7554 (.I0(x2514), .I1(x2515), .I2(x2516), .O(n7554));
  LUT5 #(.INIT(32'h96696996)) lut_n7555 (.I0(x2505), .I1(x2506), .I2(x2507), .I3(n7551), .I4(n7552), .O(n7555));
  LUT5 #(.INIT(32'hFF969600)) lut_n7556 (.I0(x2511), .I1(x2512), .I2(x2513), .I3(n7554), .I4(n7555), .O(n7556));
  LUT3 #(.INIT(8'h96)) lut_n7557 (.I0(n7545), .I1(n7548), .I2(n7549), .O(n7557));
  LUT3 #(.INIT(8'hE8)) lut_n7558 (.I0(n7553), .I1(n7556), .I2(n7557), .O(n7558));
  LUT3 #(.INIT(8'h96)) lut_n7559 (.I0(n7530), .I1(n7538), .I2(n7539), .O(n7559));
  LUT3 #(.INIT(8'hE8)) lut_n7560 (.I0(n7550), .I1(n7558), .I2(n7559), .O(n7560));
  LUT3 #(.INIT(8'h96)) lut_n7561 (.I0(x2520), .I1(x2521), .I2(x2522), .O(n7561));
  LUT5 #(.INIT(32'h96696996)) lut_n7562 (.I0(x2511), .I1(x2512), .I2(x2513), .I3(n7554), .I4(n7555), .O(n7562));
  LUT5 #(.INIT(32'hFF969600)) lut_n7563 (.I0(x2517), .I1(x2518), .I2(x2519), .I3(n7561), .I4(n7562), .O(n7563));
  LUT3 #(.INIT(8'h96)) lut_n7564 (.I0(x2526), .I1(x2527), .I2(x2528), .O(n7564));
  LUT5 #(.INIT(32'h96696996)) lut_n7565 (.I0(x2517), .I1(x2518), .I2(x2519), .I3(n7561), .I4(n7562), .O(n7565));
  LUT5 #(.INIT(32'hFF969600)) lut_n7566 (.I0(x2523), .I1(x2524), .I2(x2525), .I3(n7564), .I4(n7565), .O(n7566));
  LUT3 #(.INIT(8'h96)) lut_n7567 (.I0(n7553), .I1(n7556), .I2(n7557), .O(n7567));
  LUT3 #(.INIT(8'hE8)) lut_n7568 (.I0(n7563), .I1(n7566), .I2(n7567), .O(n7568));
  LUT3 #(.INIT(8'h96)) lut_n7569 (.I0(x2532), .I1(x2533), .I2(x2534), .O(n7569));
  LUT5 #(.INIT(32'h96696996)) lut_n7570 (.I0(x2523), .I1(x2524), .I2(x2525), .I3(n7564), .I4(n7565), .O(n7570));
  LUT5 #(.INIT(32'hFF969600)) lut_n7571 (.I0(x2529), .I1(x2530), .I2(x2531), .I3(n7569), .I4(n7570), .O(n7571));
  LUT3 #(.INIT(8'h96)) lut_n7572 (.I0(x2538), .I1(x2539), .I2(x2540), .O(n7572));
  LUT5 #(.INIT(32'h96696996)) lut_n7573 (.I0(x2529), .I1(x2530), .I2(x2531), .I3(n7569), .I4(n7570), .O(n7573));
  LUT5 #(.INIT(32'hFF969600)) lut_n7574 (.I0(x2535), .I1(x2536), .I2(x2537), .I3(n7572), .I4(n7573), .O(n7574));
  LUT3 #(.INIT(8'h96)) lut_n7575 (.I0(n7563), .I1(n7566), .I2(n7567), .O(n7575));
  LUT3 #(.INIT(8'hE8)) lut_n7576 (.I0(n7571), .I1(n7574), .I2(n7575), .O(n7576));
  LUT3 #(.INIT(8'h96)) lut_n7577 (.I0(n7550), .I1(n7558), .I2(n7559), .O(n7577));
  LUT3 #(.INIT(8'hE8)) lut_n7578 (.I0(n7568), .I1(n7576), .I2(n7577), .O(n7578));
  LUT3 #(.INIT(8'h96)) lut_n7579 (.I0(n7522), .I1(n7540), .I2(n7541), .O(n7579));
  LUT3 #(.INIT(8'hE8)) lut_n7580 (.I0(n7560), .I1(n7578), .I2(n7579), .O(n7580));
  LUT3 #(.INIT(8'h96)) lut_n7581 (.I0(n7458), .I1(n7496), .I2(n7497), .O(n7581));
  LUT3 #(.INIT(8'hE8)) lut_n7582 (.I0(n7542), .I1(n7580), .I2(n7581), .O(n7582));
  LUT3 #(.INIT(8'h96)) lut_n7583 (.I0(x2544), .I1(x2545), .I2(x2546), .O(n7583));
  LUT5 #(.INIT(32'h96696996)) lut_n7584 (.I0(x2535), .I1(x2536), .I2(x2537), .I3(n7572), .I4(n7573), .O(n7584));
  LUT5 #(.INIT(32'hFF969600)) lut_n7585 (.I0(x2541), .I1(x2542), .I2(x2543), .I3(n7583), .I4(n7584), .O(n7585));
  LUT3 #(.INIT(8'h96)) lut_n7586 (.I0(x2550), .I1(x2551), .I2(x2552), .O(n7586));
  LUT5 #(.INIT(32'h96696996)) lut_n7587 (.I0(x2541), .I1(x2542), .I2(x2543), .I3(n7583), .I4(n7584), .O(n7587));
  LUT5 #(.INIT(32'hFF969600)) lut_n7588 (.I0(x2547), .I1(x2548), .I2(x2549), .I3(n7586), .I4(n7587), .O(n7588));
  LUT3 #(.INIT(8'h96)) lut_n7589 (.I0(n7571), .I1(n7574), .I2(n7575), .O(n7589));
  LUT3 #(.INIT(8'hE8)) lut_n7590 (.I0(n7585), .I1(n7588), .I2(n7589), .O(n7590));
  LUT3 #(.INIT(8'h96)) lut_n7591 (.I0(x2556), .I1(x2557), .I2(x2558), .O(n7591));
  LUT5 #(.INIT(32'h96696996)) lut_n7592 (.I0(x2547), .I1(x2548), .I2(x2549), .I3(n7586), .I4(n7587), .O(n7592));
  LUT5 #(.INIT(32'hFF969600)) lut_n7593 (.I0(x2553), .I1(x2554), .I2(x2555), .I3(n7591), .I4(n7592), .O(n7593));
  LUT3 #(.INIT(8'h96)) lut_n7594 (.I0(x2562), .I1(x2563), .I2(x2564), .O(n7594));
  LUT5 #(.INIT(32'h96696996)) lut_n7595 (.I0(x2553), .I1(x2554), .I2(x2555), .I3(n7591), .I4(n7592), .O(n7595));
  LUT5 #(.INIT(32'hFF969600)) lut_n7596 (.I0(x2559), .I1(x2560), .I2(x2561), .I3(n7594), .I4(n7595), .O(n7596));
  LUT3 #(.INIT(8'h96)) lut_n7597 (.I0(n7585), .I1(n7588), .I2(n7589), .O(n7597));
  LUT3 #(.INIT(8'hE8)) lut_n7598 (.I0(n7593), .I1(n7596), .I2(n7597), .O(n7598));
  LUT3 #(.INIT(8'h96)) lut_n7599 (.I0(n7568), .I1(n7576), .I2(n7577), .O(n7599));
  LUT3 #(.INIT(8'hE8)) lut_n7600 (.I0(n7590), .I1(n7598), .I2(n7599), .O(n7600));
  LUT3 #(.INIT(8'h96)) lut_n7601 (.I0(x2568), .I1(x2569), .I2(x2570), .O(n7601));
  LUT5 #(.INIT(32'h96696996)) lut_n7602 (.I0(x2559), .I1(x2560), .I2(x2561), .I3(n7594), .I4(n7595), .O(n7602));
  LUT5 #(.INIT(32'hFF969600)) lut_n7603 (.I0(x2565), .I1(x2566), .I2(x2567), .I3(n7601), .I4(n7602), .O(n7603));
  LUT3 #(.INIT(8'h96)) lut_n7604 (.I0(x2574), .I1(x2575), .I2(x2576), .O(n7604));
  LUT5 #(.INIT(32'h96696996)) lut_n7605 (.I0(x2565), .I1(x2566), .I2(x2567), .I3(n7601), .I4(n7602), .O(n7605));
  LUT5 #(.INIT(32'hFF969600)) lut_n7606 (.I0(x2571), .I1(x2572), .I2(x2573), .I3(n7604), .I4(n7605), .O(n7606));
  LUT3 #(.INIT(8'h96)) lut_n7607 (.I0(n7593), .I1(n7596), .I2(n7597), .O(n7607));
  LUT3 #(.INIT(8'hE8)) lut_n7608 (.I0(n7603), .I1(n7606), .I2(n7607), .O(n7608));
  LUT3 #(.INIT(8'h96)) lut_n7609 (.I0(x2580), .I1(x2581), .I2(x2582), .O(n7609));
  LUT5 #(.INIT(32'h96696996)) lut_n7610 (.I0(x2571), .I1(x2572), .I2(x2573), .I3(n7604), .I4(n7605), .O(n7610));
  LUT5 #(.INIT(32'hFF969600)) lut_n7611 (.I0(x2577), .I1(x2578), .I2(x2579), .I3(n7609), .I4(n7610), .O(n7611));
  LUT3 #(.INIT(8'h96)) lut_n7612 (.I0(x2586), .I1(x2587), .I2(x2588), .O(n7612));
  LUT5 #(.INIT(32'h96696996)) lut_n7613 (.I0(x2577), .I1(x2578), .I2(x2579), .I3(n7609), .I4(n7610), .O(n7613));
  LUT5 #(.INIT(32'hFF969600)) lut_n7614 (.I0(x2583), .I1(x2584), .I2(x2585), .I3(n7612), .I4(n7613), .O(n7614));
  LUT3 #(.INIT(8'h96)) lut_n7615 (.I0(n7603), .I1(n7606), .I2(n7607), .O(n7615));
  LUT3 #(.INIT(8'hE8)) lut_n7616 (.I0(n7611), .I1(n7614), .I2(n7615), .O(n7616));
  LUT3 #(.INIT(8'h96)) lut_n7617 (.I0(n7590), .I1(n7598), .I2(n7599), .O(n7617));
  LUT3 #(.INIT(8'hE8)) lut_n7618 (.I0(n7608), .I1(n7616), .I2(n7617), .O(n7618));
  LUT3 #(.INIT(8'h96)) lut_n7619 (.I0(n7560), .I1(n7578), .I2(n7579), .O(n7619));
  LUT3 #(.INIT(8'hE8)) lut_n7620 (.I0(n7600), .I1(n7618), .I2(n7619), .O(n7620));
  LUT3 #(.INIT(8'h96)) lut_n7621 (.I0(x2592), .I1(x2593), .I2(x2594), .O(n7621));
  LUT5 #(.INIT(32'h96696996)) lut_n7622 (.I0(x2583), .I1(x2584), .I2(x2585), .I3(n7612), .I4(n7613), .O(n7622));
  LUT5 #(.INIT(32'hFF969600)) lut_n7623 (.I0(x2589), .I1(x2590), .I2(x2591), .I3(n7621), .I4(n7622), .O(n7623));
  LUT3 #(.INIT(8'h96)) lut_n7624 (.I0(x2598), .I1(x2599), .I2(x2600), .O(n7624));
  LUT5 #(.INIT(32'h96696996)) lut_n7625 (.I0(x2589), .I1(x2590), .I2(x2591), .I3(n7621), .I4(n7622), .O(n7625));
  LUT5 #(.INIT(32'hFF969600)) lut_n7626 (.I0(x2595), .I1(x2596), .I2(x2597), .I3(n7624), .I4(n7625), .O(n7626));
  LUT3 #(.INIT(8'h96)) lut_n7627 (.I0(n7611), .I1(n7614), .I2(n7615), .O(n7627));
  LUT3 #(.INIT(8'hE8)) lut_n7628 (.I0(n7623), .I1(n7626), .I2(n7627), .O(n7628));
  LUT3 #(.INIT(8'h96)) lut_n7629 (.I0(x2604), .I1(x2605), .I2(x2606), .O(n7629));
  LUT5 #(.INIT(32'h96696996)) lut_n7630 (.I0(x2595), .I1(x2596), .I2(x2597), .I3(n7624), .I4(n7625), .O(n7630));
  LUT5 #(.INIT(32'hFF969600)) lut_n7631 (.I0(x2601), .I1(x2602), .I2(x2603), .I3(n7629), .I4(n7630), .O(n7631));
  LUT3 #(.INIT(8'h96)) lut_n7632 (.I0(x2610), .I1(x2611), .I2(x2612), .O(n7632));
  LUT5 #(.INIT(32'h96696996)) lut_n7633 (.I0(x2601), .I1(x2602), .I2(x2603), .I3(n7629), .I4(n7630), .O(n7633));
  LUT5 #(.INIT(32'hFF969600)) lut_n7634 (.I0(x2607), .I1(x2608), .I2(x2609), .I3(n7632), .I4(n7633), .O(n7634));
  LUT3 #(.INIT(8'h96)) lut_n7635 (.I0(n7623), .I1(n7626), .I2(n7627), .O(n7635));
  LUT3 #(.INIT(8'hE8)) lut_n7636 (.I0(n7631), .I1(n7634), .I2(n7635), .O(n7636));
  LUT3 #(.INIT(8'h96)) lut_n7637 (.I0(n7608), .I1(n7616), .I2(n7617), .O(n7637));
  LUT3 #(.INIT(8'hE8)) lut_n7638 (.I0(n7628), .I1(n7636), .I2(n7637), .O(n7638));
  LUT3 #(.INIT(8'h96)) lut_n7639 (.I0(x2616), .I1(x2617), .I2(x2618), .O(n7639));
  LUT5 #(.INIT(32'h96696996)) lut_n7640 (.I0(x2607), .I1(x2608), .I2(x2609), .I3(n7632), .I4(n7633), .O(n7640));
  LUT5 #(.INIT(32'hFF969600)) lut_n7641 (.I0(x2613), .I1(x2614), .I2(x2615), .I3(n7639), .I4(n7640), .O(n7641));
  LUT3 #(.INIT(8'h96)) lut_n7642 (.I0(x2622), .I1(x2623), .I2(x2624), .O(n7642));
  LUT5 #(.INIT(32'h96696996)) lut_n7643 (.I0(x2613), .I1(x2614), .I2(x2615), .I3(n7639), .I4(n7640), .O(n7643));
  LUT5 #(.INIT(32'hFF969600)) lut_n7644 (.I0(x2619), .I1(x2620), .I2(x2621), .I3(n7642), .I4(n7643), .O(n7644));
  LUT3 #(.INIT(8'h96)) lut_n7645 (.I0(n7631), .I1(n7634), .I2(n7635), .O(n7645));
  LUT3 #(.INIT(8'hE8)) lut_n7646 (.I0(n7641), .I1(n7644), .I2(n7645), .O(n7646));
  LUT3 #(.INIT(8'h96)) lut_n7647 (.I0(x2628), .I1(x2629), .I2(x2630), .O(n7647));
  LUT5 #(.INIT(32'h96696996)) lut_n7648 (.I0(x2619), .I1(x2620), .I2(x2621), .I3(n7642), .I4(n7643), .O(n7648));
  LUT5 #(.INIT(32'hFF969600)) lut_n7649 (.I0(x2625), .I1(x2626), .I2(x2627), .I3(n7647), .I4(n7648), .O(n7649));
  LUT3 #(.INIT(8'h96)) lut_n7650 (.I0(x2634), .I1(x2635), .I2(x2636), .O(n7650));
  LUT5 #(.INIT(32'h96696996)) lut_n7651 (.I0(x2625), .I1(x2626), .I2(x2627), .I3(n7647), .I4(n7648), .O(n7651));
  LUT5 #(.INIT(32'hFF969600)) lut_n7652 (.I0(x2631), .I1(x2632), .I2(x2633), .I3(n7650), .I4(n7651), .O(n7652));
  LUT3 #(.INIT(8'h96)) lut_n7653 (.I0(n7641), .I1(n7644), .I2(n7645), .O(n7653));
  LUT3 #(.INIT(8'hE8)) lut_n7654 (.I0(n7649), .I1(n7652), .I2(n7653), .O(n7654));
  LUT3 #(.INIT(8'h96)) lut_n7655 (.I0(n7628), .I1(n7636), .I2(n7637), .O(n7655));
  LUT3 #(.INIT(8'hE8)) lut_n7656 (.I0(n7646), .I1(n7654), .I2(n7655), .O(n7656));
  LUT3 #(.INIT(8'h96)) lut_n7657 (.I0(n7600), .I1(n7618), .I2(n7619), .O(n7657));
  LUT3 #(.INIT(8'hE8)) lut_n7658 (.I0(n7638), .I1(n7656), .I2(n7657), .O(n7658));
  LUT3 #(.INIT(8'h96)) lut_n7659 (.I0(n7542), .I1(n7580), .I2(n7581), .O(n7659));
  LUT3 #(.INIT(8'hE8)) lut_n7660 (.I0(n7620), .I1(n7658), .I2(n7659), .O(n7660));
  LUT3 #(.INIT(8'h96)) lut_n7661 (.I0(n7420), .I1(n7498), .I2(n7499), .O(n7661));
  LUT3 #(.INIT(8'hE8)) lut_n7662 (.I0(n7582), .I1(n7660), .I2(n7661), .O(n7662));
  LUT3 #(.INIT(8'h96)) lut_n7663 (.I0(x2640), .I1(x2641), .I2(x2642), .O(n7663));
  LUT5 #(.INIT(32'h96696996)) lut_n7664 (.I0(x2631), .I1(x2632), .I2(x2633), .I3(n7650), .I4(n7651), .O(n7664));
  LUT5 #(.INIT(32'hFF969600)) lut_n7665 (.I0(x2637), .I1(x2638), .I2(x2639), .I3(n7663), .I4(n7664), .O(n7665));
  LUT3 #(.INIT(8'h96)) lut_n7666 (.I0(x2646), .I1(x2647), .I2(x2648), .O(n7666));
  LUT5 #(.INIT(32'h96696996)) lut_n7667 (.I0(x2637), .I1(x2638), .I2(x2639), .I3(n7663), .I4(n7664), .O(n7667));
  LUT5 #(.INIT(32'hFF969600)) lut_n7668 (.I0(x2643), .I1(x2644), .I2(x2645), .I3(n7666), .I4(n7667), .O(n7668));
  LUT3 #(.INIT(8'h96)) lut_n7669 (.I0(n7649), .I1(n7652), .I2(n7653), .O(n7669));
  LUT3 #(.INIT(8'hE8)) lut_n7670 (.I0(n7665), .I1(n7668), .I2(n7669), .O(n7670));
  LUT3 #(.INIT(8'h96)) lut_n7671 (.I0(x2652), .I1(x2653), .I2(x2654), .O(n7671));
  LUT5 #(.INIT(32'h96696996)) lut_n7672 (.I0(x2643), .I1(x2644), .I2(x2645), .I3(n7666), .I4(n7667), .O(n7672));
  LUT5 #(.INIT(32'hFF969600)) lut_n7673 (.I0(x2649), .I1(x2650), .I2(x2651), .I3(n7671), .I4(n7672), .O(n7673));
  LUT3 #(.INIT(8'h96)) lut_n7674 (.I0(x2658), .I1(x2659), .I2(x2660), .O(n7674));
  LUT5 #(.INIT(32'h96696996)) lut_n7675 (.I0(x2649), .I1(x2650), .I2(x2651), .I3(n7671), .I4(n7672), .O(n7675));
  LUT5 #(.INIT(32'hFF969600)) lut_n7676 (.I0(x2655), .I1(x2656), .I2(x2657), .I3(n7674), .I4(n7675), .O(n7676));
  LUT3 #(.INIT(8'h96)) lut_n7677 (.I0(n7665), .I1(n7668), .I2(n7669), .O(n7677));
  LUT3 #(.INIT(8'hE8)) lut_n7678 (.I0(n7673), .I1(n7676), .I2(n7677), .O(n7678));
  LUT3 #(.INIT(8'h96)) lut_n7679 (.I0(n7646), .I1(n7654), .I2(n7655), .O(n7679));
  LUT3 #(.INIT(8'hE8)) lut_n7680 (.I0(n7670), .I1(n7678), .I2(n7679), .O(n7680));
  LUT3 #(.INIT(8'h96)) lut_n7681 (.I0(x2664), .I1(x2665), .I2(x2666), .O(n7681));
  LUT5 #(.INIT(32'h96696996)) lut_n7682 (.I0(x2655), .I1(x2656), .I2(x2657), .I3(n7674), .I4(n7675), .O(n7682));
  LUT5 #(.INIT(32'hFF969600)) lut_n7683 (.I0(x2661), .I1(x2662), .I2(x2663), .I3(n7681), .I4(n7682), .O(n7683));
  LUT3 #(.INIT(8'h96)) lut_n7684 (.I0(x2670), .I1(x2671), .I2(x2672), .O(n7684));
  LUT5 #(.INIT(32'h96696996)) lut_n7685 (.I0(x2661), .I1(x2662), .I2(x2663), .I3(n7681), .I4(n7682), .O(n7685));
  LUT5 #(.INIT(32'hFF969600)) lut_n7686 (.I0(x2667), .I1(x2668), .I2(x2669), .I3(n7684), .I4(n7685), .O(n7686));
  LUT3 #(.INIT(8'h96)) lut_n7687 (.I0(n7673), .I1(n7676), .I2(n7677), .O(n7687));
  LUT3 #(.INIT(8'hE8)) lut_n7688 (.I0(n7683), .I1(n7686), .I2(n7687), .O(n7688));
  LUT3 #(.INIT(8'h96)) lut_n7689 (.I0(x2676), .I1(x2677), .I2(x2678), .O(n7689));
  LUT5 #(.INIT(32'h96696996)) lut_n7690 (.I0(x2667), .I1(x2668), .I2(x2669), .I3(n7684), .I4(n7685), .O(n7690));
  LUT5 #(.INIT(32'hFF969600)) lut_n7691 (.I0(x2673), .I1(x2674), .I2(x2675), .I3(n7689), .I4(n7690), .O(n7691));
  LUT3 #(.INIT(8'h96)) lut_n7692 (.I0(x2682), .I1(x2683), .I2(x2684), .O(n7692));
  LUT5 #(.INIT(32'h96696996)) lut_n7693 (.I0(x2673), .I1(x2674), .I2(x2675), .I3(n7689), .I4(n7690), .O(n7693));
  LUT5 #(.INIT(32'hFF969600)) lut_n7694 (.I0(x2679), .I1(x2680), .I2(x2681), .I3(n7692), .I4(n7693), .O(n7694));
  LUT3 #(.INIT(8'h96)) lut_n7695 (.I0(n7683), .I1(n7686), .I2(n7687), .O(n7695));
  LUT3 #(.INIT(8'hE8)) lut_n7696 (.I0(n7691), .I1(n7694), .I2(n7695), .O(n7696));
  LUT3 #(.INIT(8'h96)) lut_n7697 (.I0(n7670), .I1(n7678), .I2(n7679), .O(n7697));
  LUT3 #(.INIT(8'hE8)) lut_n7698 (.I0(n7688), .I1(n7696), .I2(n7697), .O(n7698));
  LUT3 #(.INIT(8'h96)) lut_n7699 (.I0(n7638), .I1(n7656), .I2(n7657), .O(n7699));
  LUT3 #(.INIT(8'hE8)) lut_n7700 (.I0(n7680), .I1(n7698), .I2(n7699), .O(n7700));
  LUT3 #(.INIT(8'h96)) lut_n7701 (.I0(x2688), .I1(x2689), .I2(x2690), .O(n7701));
  LUT5 #(.INIT(32'h96696996)) lut_n7702 (.I0(x2679), .I1(x2680), .I2(x2681), .I3(n7692), .I4(n7693), .O(n7702));
  LUT5 #(.INIT(32'hFF969600)) lut_n7703 (.I0(x2685), .I1(x2686), .I2(x2687), .I3(n7701), .I4(n7702), .O(n7703));
  LUT3 #(.INIT(8'h96)) lut_n7704 (.I0(x2694), .I1(x2695), .I2(x2696), .O(n7704));
  LUT5 #(.INIT(32'h96696996)) lut_n7705 (.I0(x2685), .I1(x2686), .I2(x2687), .I3(n7701), .I4(n7702), .O(n7705));
  LUT5 #(.INIT(32'hFF969600)) lut_n7706 (.I0(x2691), .I1(x2692), .I2(x2693), .I3(n7704), .I4(n7705), .O(n7706));
  LUT3 #(.INIT(8'h96)) lut_n7707 (.I0(n7691), .I1(n7694), .I2(n7695), .O(n7707));
  LUT3 #(.INIT(8'hE8)) lut_n7708 (.I0(n7703), .I1(n7706), .I2(n7707), .O(n7708));
  LUT3 #(.INIT(8'h96)) lut_n7709 (.I0(x2700), .I1(x2701), .I2(x2702), .O(n7709));
  LUT5 #(.INIT(32'h96696996)) lut_n7710 (.I0(x2691), .I1(x2692), .I2(x2693), .I3(n7704), .I4(n7705), .O(n7710));
  LUT5 #(.INIT(32'hFF969600)) lut_n7711 (.I0(x2697), .I1(x2698), .I2(x2699), .I3(n7709), .I4(n7710), .O(n7711));
  LUT3 #(.INIT(8'h96)) lut_n7712 (.I0(x2706), .I1(x2707), .I2(x2708), .O(n7712));
  LUT5 #(.INIT(32'h96696996)) lut_n7713 (.I0(x2697), .I1(x2698), .I2(x2699), .I3(n7709), .I4(n7710), .O(n7713));
  LUT5 #(.INIT(32'hFF969600)) lut_n7714 (.I0(x2703), .I1(x2704), .I2(x2705), .I3(n7712), .I4(n7713), .O(n7714));
  LUT3 #(.INIT(8'h96)) lut_n7715 (.I0(n7703), .I1(n7706), .I2(n7707), .O(n7715));
  LUT3 #(.INIT(8'hE8)) lut_n7716 (.I0(n7711), .I1(n7714), .I2(n7715), .O(n7716));
  LUT3 #(.INIT(8'h96)) lut_n7717 (.I0(n7688), .I1(n7696), .I2(n7697), .O(n7717));
  LUT3 #(.INIT(8'hE8)) lut_n7718 (.I0(n7708), .I1(n7716), .I2(n7717), .O(n7718));
  LUT3 #(.INIT(8'h96)) lut_n7719 (.I0(x2712), .I1(x2713), .I2(x2714), .O(n7719));
  LUT5 #(.INIT(32'h96696996)) lut_n7720 (.I0(x2703), .I1(x2704), .I2(x2705), .I3(n7712), .I4(n7713), .O(n7720));
  LUT5 #(.INIT(32'hFF969600)) lut_n7721 (.I0(x2709), .I1(x2710), .I2(x2711), .I3(n7719), .I4(n7720), .O(n7721));
  LUT3 #(.INIT(8'h96)) lut_n7722 (.I0(x2718), .I1(x2719), .I2(x2720), .O(n7722));
  LUT5 #(.INIT(32'h96696996)) lut_n7723 (.I0(x2709), .I1(x2710), .I2(x2711), .I3(n7719), .I4(n7720), .O(n7723));
  LUT5 #(.INIT(32'hFF969600)) lut_n7724 (.I0(x2715), .I1(x2716), .I2(x2717), .I3(n7722), .I4(n7723), .O(n7724));
  LUT3 #(.INIT(8'h96)) lut_n7725 (.I0(n7711), .I1(n7714), .I2(n7715), .O(n7725));
  LUT3 #(.INIT(8'hE8)) lut_n7726 (.I0(n7721), .I1(n7724), .I2(n7725), .O(n7726));
  LUT3 #(.INIT(8'h96)) lut_n7727 (.I0(x2724), .I1(x2725), .I2(x2726), .O(n7727));
  LUT5 #(.INIT(32'h96696996)) lut_n7728 (.I0(x2715), .I1(x2716), .I2(x2717), .I3(n7722), .I4(n7723), .O(n7728));
  LUT5 #(.INIT(32'hFF969600)) lut_n7729 (.I0(x2721), .I1(x2722), .I2(x2723), .I3(n7727), .I4(n7728), .O(n7729));
  LUT3 #(.INIT(8'h96)) lut_n7730 (.I0(x2730), .I1(x2731), .I2(x2732), .O(n7730));
  LUT5 #(.INIT(32'h96696996)) lut_n7731 (.I0(x2721), .I1(x2722), .I2(x2723), .I3(n7727), .I4(n7728), .O(n7731));
  LUT5 #(.INIT(32'hFF969600)) lut_n7732 (.I0(x2727), .I1(x2728), .I2(x2729), .I3(n7730), .I4(n7731), .O(n7732));
  LUT3 #(.INIT(8'h96)) lut_n7733 (.I0(n7721), .I1(n7724), .I2(n7725), .O(n7733));
  LUT3 #(.INIT(8'hE8)) lut_n7734 (.I0(n7729), .I1(n7732), .I2(n7733), .O(n7734));
  LUT3 #(.INIT(8'h96)) lut_n7735 (.I0(n7708), .I1(n7716), .I2(n7717), .O(n7735));
  LUT3 #(.INIT(8'hE8)) lut_n7736 (.I0(n7726), .I1(n7734), .I2(n7735), .O(n7736));
  LUT3 #(.INIT(8'h96)) lut_n7737 (.I0(n7680), .I1(n7698), .I2(n7699), .O(n7737));
  LUT3 #(.INIT(8'hE8)) lut_n7738 (.I0(n7718), .I1(n7736), .I2(n7737), .O(n7738));
  LUT3 #(.INIT(8'h96)) lut_n7739 (.I0(n7620), .I1(n7658), .I2(n7659), .O(n7739));
  LUT3 #(.INIT(8'hE8)) lut_n7740 (.I0(n7700), .I1(n7738), .I2(n7739), .O(n7740));
  LUT3 #(.INIT(8'h96)) lut_n7741 (.I0(x2736), .I1(x2737), .I2(x2738), .O(n7741));
  LUT5 #(.INIT(32'h96696996)) lut_n7742 (.I0(x2727), .I1(x2728), .I2(x2729), .I3(n7730), .I4(n7731), .O(n7742));
  LUT5 #(.INIT(32'hFF969600)) lut_n7743 (.I0(x2733), .I1(x2734), .I2(x2735), .I3(n7741), .I4(n7742), .O(n7743));
  LUT3 #(.INIT(8'h96)) lut_n7744 (.I0(x2742), .I1(x2743), .I2(x2744), .O(n7744));
  LUT5 #(.INIT(32'h96696996)) lut_n7745 (.I0(x2733), .I1(x2734), .I2(x2735), .I3(n7741), .I4(n7742), .O(n7745));
  LUT5 #(.INIT(32'hFF969600)) lut_n7746 (.I0(x2739), .I1(x2740), .I2(x2741), .I3(n7744), .I4(n7745), .O(n7746));
  LUT3 #(.INIT(8'h96)) lut_n7747 (.I0(n7729), .I1(n7732), .I2(n7733), .O(n7747));
  LUT3 #(.INIT(8'hE8)) lut_n7748 (.I0(n7743), .I1(n7746), .I2(n7747), .O(n7748));
  LUT3 #(.INIT(8'h96)) lut_n7749 (.I0(x2748), .I1(x2749), .I2(x2750), .O(n7749));
  LUT5 #(.INIT(32'h96696996)) lut_n7750 (.I0(x2739), .I1(x2740), .I2(x2741), .I3(n7744), .I4(n7745), .O(n7750));
  LUT5 #(.INIT(32'hFF969600)) lut_n7751 (.I0(x2745), .I1(x2746), .I2(x2747), .I3(n7749), .I4(n7750), .O(n7751));
  LUT3 #(.INIT(8'h96)) lut_n7752 (.I0(x2754), .I1(x2755), .I2(x2756), .O(n7752));
  LUT5 #(.INIT(32'h96696996)) lut_n7753 (.I0(x2745), .I1(x2746), .I2(x2747), .I3(n7749), .I4(n7750), .O(n7753));
  LUT5 #(.INIT(32'hFF969600)) lut_n7754 (.I0(x2751), .I1(x2752), .I2(x2753), .I3(n7752), .I4(n7753), .O(n7754));
  LUT3 #(.INIT(8'h96)) lut_n7755 (.I0(n7743), .I1(n7746), .I2(n7747), .O(n7755));
  LUT3 #(.INIT(8'hE8)) lut_n7756 (.I0(n7751), .I1(n7754), .I2(n7755), .O(n7756));
  LUT3 #(.INIT(8'h96)) lut_n7757 (.I0(n7726), .I1(n7734), .I2(n7735), .O(n7757));
  LUT3 #(.INIT(8'hE8)) lut_n7758 (.I0(n7748), .I1(n7756), .I2(n7757), .O(n7758));
  LUT3 #(.INIT(8'h96)) lut_n7759 (.I0(x2760), .I1(x2761), .I2(x2762), .O(n7759));
  LUT5 #(.INIT(32'h96696996)) lut_n7760 (.I0(x2751), .I1(x2752), .I2(x2753), .I3(n7752), .I4(n7753), .O(n7760));
  LUT5 #(.INIT(32'hFF969600)) lut_n7761 (.I0(x2757), .I1(x2758), .I2(x2759), .I3(n7759), .I4(n7760), .O(n7761));
  LUT3 #(.INIT(8'h96)) lut_n7762 (.I0(x2766), .I1(x2767), .I2(x2768), .O(n7762));
  LUT5 #(.INIT(32'h96696996)) lut_n7763 (.I0(x2757), .I1(x2758), .I2(x2759), .I3(n7759), .I4(n7760), .O(n7763));
  LUT5 #(.INIT(32'hFF969600)) lut_n7764 (.I0(x2763), .I1(x2764), .I2(x2765), .I3(n7762), .I4(n7763), .O(n7764));
  LUT3 #(.INIT(8'h96)) lut_n7765 (.I0(n7751), .I1(n7754), .I2(n7755), .O(n7765));
  LUT3 #(.INIT(8'hE8)) lut_n7766 (.I0(n7761), .I1(n7764), .I2(n7765), .O(n7766));
  LUT3 #(.INIT(8'h96)) lut_n7767 (.I0(x2772), .I1(x2773), .I2(x2774), .O(n7767));
  LUT5 #(.INIT(32'h96696996)) lut_n7768 (.I0(x2763), .I1(x2764), .I2(x2765), .I3(n7762), .I4(n7763), .O(n7768));
  LUT5 #(.INIT(32'hFF969600)) lut_n7769 (.I0(x2769), .I1(x2770), .I2(x2771), .I3(n7767), .I4(n7768), .O(n7769));
  LUT3 #(.INIT(8'h96)) lut_n7770 (.I0(x2778), .I1(x2779), .I2(x2780), .O(n7770));
  LUT5 #(.INIT(32'h96696996)) lut_n7771 (.I0(x2769), .I1(x2770), .I2(x2771), .I3(n7767), .I4(n7768), .O(n7771));
  LUT5 #(.INIT(32'hFF969600)) lut_n7772 (.I0(x2775), .I1(x2776), .I2(x2777), .I3(n7770), .I4(n7771), .O(n7772));
  LUT3 #(.INIT(8'h96)) lut_n7773 (.I0(n7761), .I1(n7764), .I2(n7765), .O(n7773));
  LUT3 #(.INIT(8'hE8)) lut_n7774 (.I0(n7769), .I1(n7772), .I2(n7773), .O(n7774));
  LUT3 #(.INIT(8'h96)) lut_n7775 (.I0(n7748), .I1(n7756), .I2(n7757), .O(n7775));
  LUT3 #(.INIT(8'hE8)) lut_n7776 (.I0(n7766), .I1(n7774), .I2(n7775), .O(n7776));
  LUT3 #(.INIT(8'h96)) lut_n7777 (.I0(n7718), .I1(n7736), .I2(n7737), .O(n7777));
  LUT3 #(.INIT(8'hE8)) lut_n7778 (.I0(n7758), .I1(n7776), .I2(n7777), .O(n7778));
  LUT3 #(.INIT(8'h96)) lut_n7779 (.I0(x2784), .I1(x2785), .I2(x2786), .O(n7779));
  LUT5 #(.INIT(32'h96696996)) lut_n7780 (.I0(x2775), .I1(x2776), .I2(x2777), .I3(n7770), .I4(n7771), .O(n7780));
  LUT5 #(.INIT(32'hFF969600)) lut_n7781 (.I0(x2781), .I1(x2782), .I2(x2783), .I3(n7779), .I4(n7780), .O(n7781));
  LUT3 #(.INIT(8'h96)) lut_n7782 (.I0(x2790), .I1(x2791), .I2(x2792), .O(n7782));
  LUT5 #(.INIT(32'h96696996)) lut_n7783 (.I0(x2781), .I1(x2782), .I2(x2783), .I3(n7779), .I4(n7780), .O(n7783));
  LUT5 #(.INIT(32'hFF969600)) lut_n7784 (.I0(x2787), .I1(x2788), .I2(x2789), .I3(n7782), .I4(n7783), .O(n7784));
  LUT3 #(.INIT(8'h96)) lut_n7785 (.I0(n7769), .I1(n7772), .I2(n7773), .O(n7785));
  LUT3 #(.INIT(8'hE8)) lut_n7786 (.I0(n7781), .I1(n7784), .I2(n7785), .O(n7786));
  LUT3 #(.INIT(8'h96)) lut_n7787 (.I0(x2796), .I1(x2797), .I2(x2798), .O(n7787));
  LUT5 #(.INIT(32'h96696996)) lut_n7788 (.I0(x2787), .I1(x2788), .I2(x2789), .I3(n7782), .I4(n7783), .O(n7788));
  LUT5 #(.INIT(32'hFF969600)) lut_n7789 (.I0(x2793), .I1(x2794), .I2(x2795), .I3(n7787), .I4(n7788), .O(n7789));
  LUT3 #(.INIT(8'h96)) lut_n7790 (.I0(x2802), .I1(x2803), .I2(x2804), .O(n7790));
  LUT5 #(.INIT(32'h96696996)) lut_n7791 (.I0(x2793), .I1(x2794), .I2(x2795), .I3(n7787), .I4(n7788), .O(n7791));
  LUT5 #(.INIT(32'hFF969600)) lut_n7792 (.I0(x2799), .I1(x2800), .I2(x2801), .I3(n7790), .I4(n7791), .O(n7792));
  LUT3 #(.INIT(8'h96)) lut_n7793 (.I0(n7781), .I1(n7784), .I2(n7785), .O(n7793));
  LUT3 #(.INIT(8'hE8)) lut_n7794 (.I0(n7789), .I1(n7792), .I2(n7793), .O(n7794));
  LUT3 #(.INIT(8'h96)) lut_n7795 (.I0(n7766), .I1(n7774), .I2(n7775), .O(n7795));
  LUT3 #(.INIT(8'hE8)) lut_n7796 (.I0(n7786), .I1(n7794), .I2(n7795), .O(n7796));
  LUT3 #(.INIT(8'h96)) lut_n7797 (.I0(x2808), .I1(x2809), .I2(x2810), .O(n7797));
  LUT5 #(.INIT(32'h96696996)) lut_n7798 (.I0(x2799), .I1(x2800), .I2(x2801), .I3(n7790), .I4(n7791), .O(n7798));
  LUT5 #(.INIT(32'hFF969600)) lut_n7799 (.I0(x2805), .I1(x2806), .I2(x2807), .I3(n7797), .I4(n7798), .O(n7799));
  LUT3 #(.INIT(8'h96)) lut_n7800 (.I0(x2814), .I1(x2815), .I2(x2816), .O(n7800));
  LUT5 #(.INIT(32'h96696996)) lut_n7801 (.I0(x2805), .I1(x2806), .I2(x2807), .I3(n7797), .I4(n7798), .O(n7801));
  LUT5 #(.INIT(32'hFF969600)) lut_n7802 (.I0(x2811), .I1(x2812), .I2(x2813), .I3(n7800), .I4(n7801), .O(n7802));
  LUT3 #(.INIT(8'h96)) lut_n7803 (.I0(n7789), .I1(n7792), .I2(n7793), .O(n7803));
  LUT3 #(.INIT(8'hE8)) lut_n7804 (.I0(n7799), .I1(n7802), .I2(n7803), .O(n7804));
  LUT3 #(.INIT(8'h96)) lut_n7805 (.I0(x2820), .I1(x2821), .I2(x2822), .O(n7805));
  LUT5 #(.INIT(32'h96696996)) lut_n7806 (.I0(x2811), .I1(x2812), .I2(x2813), .I3(n7800), .I4(n7801), .O(n7806));
  LUT5 #(.INIT(32'hFF969600)) lut_n7807 (.I0(x2817), .I1(x2818), .I2(x2819), .I3(n7805), .I4(n7806), .O(n7807));
  LUT3 #(.INIT(8'h96)) lut_n7808 (.I0(x2826), .I1(x2827), .I2(x2828), .O(n7808));
  LUT5 #(.INIT(32'h96696996)) lut_n7809 (.I0(x2817), .I1(x2818), .I2(x2819), .I3(n7805), .I4(n7806), .O(n7809));
  LUT5 #(.INIT(32'hFF969600)) lut_n7810 (.I0(x2823), .I1(x2824), .I2(x2825), .I3(n7808), .I4(n7809), .O(n7810));
  LUT3 #(.INIT(8'h96)) lut_n7811 (.I0(n7799), .I1(n7802), .I2(n7803), .O(n7811));
  LUT3 #(.INIT(8'hE8)) lut_n7812 (.I0(n7807), .I1(n7810), .I2(n7811), .O(n7812));
  LUT3 #(.INIT(8'h96)) lut_n7813 (.I0(n7786), .I1(n7794), .I2(n7795), .O(n7813));
  LUT3 #(.INIT(8'hE8)) lut_n7814 (.I0(n7804), .I1(n7812), .I2(n7813), .O(n7814));
  LUT3 #(.INIT(8'h96)) lut_n7815 (.I0(n7758), .I1(n7776), .I2(n7777), .O(n7815));
  LUT3 #(.INIT(8'hE8)) lut_n7816 (.I0(n7796), .I1(n7814), .I2(n7815), .O(n7816));
  LUT3 #(.INIT(8'h96)) lut_n7817 (.I0(n7700), .I1(n7738), .I2(n7739), .O(n7817));
  LUT3 #(.INIT(8'hE8)) lut_n7818 (.I0(n7778), .I1(n7816), .I2(n7817), .O(n7818));
  LUT3 #(.INIT(8'h96)) lut_n7819 (.I0(n7582), .I1(n7660), .I2(n7661), .O(n7819));
  LUT3 #(.INIT(8'hE8)) lut_n7820 (.I0(n7740), .I1(n7818), .I2(n7819), .O(n7820));
  LUT3 #(.INIT(8'h96)) lut_n7821 (.I0(n7342), .I1(n7500), .I2(n7501), .O(n7821));
  LUT3 #(.INIT(8'hE8)) lut_n7822 (.I0(n7662), .I1(n7820), .I2(n7821), .O(n7822));
  LUT3 #(.INIT(8'h96)) lut_n7823 (.I0(x2832), .I1(x2833), .I2(x2834), .O(n7823));
  LUT5 #(.INIT(32'h96696996)) lut_n7824 (.I0(x2823), .I1(x2824), .I2(x2825), .I3(n7808), .I4(n7809), .O(n7824));
  LUT5 #(.INIT(32'hFF969600)) lut_n7825 (.I0(x2829), .I1(x2830), .I2(x2831), .I3(n7823), .I4(n7824), .O(n7825));
  LUT3 #(.INIT(8'h96)) lut_n7826 (.I0(x2838), .I1(x2839), .I2(x2840), .O(n7826));
  LUT5 #(.INIT(32'h96696996)) lut_n7827 (.I0(x2829), .I1(x2830), .I2(x2831), .I3(n7823), .I4(n7824), .O(n7827));
  LUT5 #(.INIT(32'hFF969600)) lut_n7828 (.I0(x2835), .I1(x2836), .I2(x2837), .I3(n7826), .I4(n7827), .O(n7828));
  LUT3 #(.INIT(8'h96)) lut_n7829 (.I0(n7807), .I1(n7810), .I2(n7811), .O(n7829));
  LUT3 #(.INIT(8'hE8)) lut_n7830 (.I0(n7825), .I1(n7828), .I2(n7829), .O(n7830));
  LUT3 #(.INIT(8'h96)) lut_n7831 (.I0(x2844), .I1(x2845), .I2(x2846), .O(n7831));
  LUT5 #(.INIT(32'h96696996)) lut_n7832 (.I0(x2835), .I1(x2836), .I2(x2837), .I3(n7826), .I4(n7827), .O(n7832));
  LUT5 #(.INIT(32'hFF969600)) lut_n7833 (.I0(x2841), .I1(x2842), .I2(x2843), .I3(n7831), .I4(n7832), .O(n7833));
  LUT3 #(.INIT(8'h96)) lut_n7834 (.I0(x2850), .I1(x2851), .I2(x2852), .O(n7834));
  LUT5 #(.INIT(32'h96696996)) lut_n7835 (.I0(x2841), .I1(x2842), .I2(x2843), .I3(n7831), .I4(n7832), .O(n7835));
  LUT5 #(.INIT(32'hFF969600)) lut_n7836 (.I0(x2847), .I1(x2848), .I2(x2849), .I3(n7834), .I4(n7835), .O(n7836));
  LUT3 #(.INIT(8'h96)) lut_n7837 (.I0(n7825), .I1(n7828), .I2(n7829), .O(n7837));
  LUT3 #(.INIT(8'hE8)) lut_n7838 (.I0(n7833), .I1(n7836), .I2(n7837), .O(n7838));
  LUT3 #(.INIT(8'h96)) lut_n7839 (.I0(n7804), .I1(n7812), .I2(n7813), .O(n7839));
  LUT3 #(.INIT(8'hE8)) lut_n7840 (.I0(n7830), .I1(n7838), .I2(n7839), .O(n7840));
  LUT3 #(.INIT(8'h96)) lut_n7841 (.I0(x2856), .I1(x2857), .I2(x2858), .O(n7841));
  LUT5 #(.INIT(32'h96696996)) lut_n7842 (.I0(x2847), .I1(x2848), .I2(x2849), .I3(n7834), .I4(n7835), .O(n7842));
  LUT5 #(.INIT(32'hFF969600)) lut_n7843 (.I0(x2853), .I1(x2854), .I2(x2855), .I3(n7841), .I4(n7842), .O(n7843));
  LUT3 #(.INIT(8'h96)) lut_n7844 (.I0(x2862), .I1(x2863), .I2(x2864), .O(n7844));
  LUT5 #(.INIT(32'h96696996)) lut_n7845 (.I0(x2853), .I1(x2854), .I2(x2855), .I3(n7841), .I4(n7842), .O(n7845));
  LUT5 #(.INIT(32'hFF969600)) lut_n7846 (.I0(x2859), .I1(x2860), .I2(x2861), .I3(n7844), .I4(n7845), .O(n7846));
  LUT3 #(.INIT(8'h96)) lut_n7847 (.I0(n7833), .I1(n7836), .I2(n7837), .O(n7847));
  LUT3 #(.INIT(8'hE8)) lut_n7848 (.I0(n7843), .I1(n7846), .I2(n7847), .O(n7848));
  LUT3 #(.INIT(8'h96)) lut_n7849 (.I0(x2868), .I1(x2869), .I2(x2870), .O(n7849));
  LUT5 #(.INIT(32'h96696996)) lut_n7850 (.I0(x2859), .I1(x2860), .I2(x2861), .I3(n7844), .I4(n7845), .O(n7850));
  LUT5 #(.INIT(32'hFF969600)) lut_n7851 (.I0(x2865), .I1(x2866), .I2(x2867), .I3(n7849), .I4(n7850), .O(n7851));
  LUT3 #(.INIT(8'h96)) lut_n7852 (.I0(x2874), .I1(x2875), .I2(x2876), .O(n7852));
  LUT5 #(.INIT(32'h96696996)) lut_n7853 (.I0(x2865), .I1(x2866), .I2(x2867), .I3(n7849), .I4(n7850), .O(n7853));
  LUT5 #(.INIT(32'hFF969600)) lut_n7854 (.I0(x2871), .I1(x2872), .I2(x2873), .I3(n7852), .I4(n7853), .O(n7854));
  LUT3 #(.INIT(8'h96)) lut_n7855 (.I0(n7843), .I1(n7846), .I2(n7847), .O(n7855));
  LUT3 #(.INIT(8'hE8)) lut_n7856 (.I0(n7851), .I1(n7854), .I2(n7855), .O(n7856));
  LUT3 #(.INIT(8'h96)) lut_n7857 (.I0(n7830), .I1(n7838), .I2(n7839), .O(n7857));
  LUT3 #(.INIT(8'hE8)) lut_n7858 (.I0(n7848), .I1(n7856), .I2(n7857), .O(n7858));
  LUT3 #(.INIT(8'h96)) lut_n7859 (.I0(n7796), .I1(n7814), .I2(n7815), .O(n7859));
  LUT3 #(.INIT(8'hE8)) lut_n7860 (.I0(n7840), .I1(n7858), .I2(n7859), .O(n7860));
  LUT3 #(.INIT(8'h96)) lut_n7861 (.I0(x2880), .I1(x2881), .I2(x2882), .O(n7861));
  LUT5 #(.INIT(32'h96696996)) lut_n7862 (.I0(x2871), .I1(x2872), .I2(x2873), .I3(n7852), .I4(n7853), .O(n7862));
  LUT5 #(.INIT(32'hFF969600)) lut_n7863 (.I0(x2877), .I1(x2878), .I2(x2879), .I3(n7861), .I4(n7862), .O(n7863));
  LUT3 #(.INIT(8'h96)) lut_n7864 (.I0(x2886), .I1(x2887), .I2(x2888), .O(n7864));
  LUT5 #(.INIT(32'h96696996)) lut_n7865 (.I0(x2877), .I1(x2878), .I2(x2879), .I3(n7861), .I4(n7862), .O(n7865));
  LUT5 #(.INIT(32'hFF969600)) lut_n7866 (.I0(x2883), .I1(x2884), .I2(x2885), .I3(n7864), .I4(n7865), .O(n7866));
  LUT3 #(.INIT(8'h96)) lut_n7867 (.I0(n7851), .I1(n7854), .I2(n7855), .O(n7867));
  LUT3 #(.INIT(8'hE8)) lut_n7868 (.I0(n7863), .I1(n7866), .I2(n7867), .O(n7868));
  LUT3 #(.INIT(8'h96)) lut_n7869 (.I0(x2892), .I1(x2893), .I2(x2894), .O(n7869));
  LUT5 #(.INIT(32'h96696996)) lut_n7870 (.I0(x2883), .I1(x2884), .I2(x2885), .I3(n7864), .I4(n7865), .O(n7870));
  LUT5 #(.INIT(32'hFF969600)) lut_n7871 (.I0(x2889), .I1(x2890), .I2(x2891), .I3(n7869), .I4(n7870), .O(n7871));
  LUT3 #(.INIT(8'h96)) lut_n7872 (.I0(x2898), .I1(x2899), .I2(x2900), .O(n7872));
  LUT5 #(.INIT(32'h96696996)) lut_n7873 (.I0(x2889), .I1(x2890), .I2(x2891), .I3(n7869), .I4(n7870), .O(n7873));
  LUT5 #(.INIT(32'hFF969600)) lut_n7874 (.I0(x2895), .I1(x2896), .I2(x2897), .I3(n7872), .I4(n7873), .O(n7874));
  LUT3 #(.INIT(8'h96)) lut_n7875 (.I0(n7863), .I1(n7866), .I2(n7867), .O(n7875));
  LUT3 #(.INIT(8'hE8)) lut_n7876 (.I0(n7871), .I1(n7874), .I2(n7875), .O(n7876));
  LUT3 #(.INIT(8'h96)) lut_n7877 (.I0(n7848), .I1(n7856), .I2(n7857), .O(n7877));
  LUT3 #(.INIT(8'hE8)) lut_n7878 (.I0(n7868), .I1(n7876), .I2(n7877), .O(n7878));
  LUT3 #(.INIT(8'h96)) lut_n7879 (.I0(x2904), .I1(x2905), .I2(x2906), .O(n7879));
  LUT5 #(.INIT(32'h96696996)) lut_n7880 (.I0(x2895), .I1(x2896), .I2(x2897), .I3(n7872), .I4(n7873), .O(n7880));
  LUT5 #(.INIT(32'hFF969600)) lut_n7881 (.I0(x2901), .I1(x2902), .I2(x2903), .I3(n7879), .I4(n7880), .O(n7881));
  LUT3 #(.INIT(8'h96)) lut_n7882 (.I0(x2910), .I1(x2911), .I2(x2912), .O(n7882));
  LUT5 #(.INIT(32'h96696996)) lut_n7883 (.I0(x2901), .I1(x2902), .I2(x2903), .I3(n7879), .I4(n7880), .O(n7883));
  LUT5 #(.INIT(32'hFF969600)) lut_n7884 (.I0(x2907), .I1(x2908), .I2(x2909), .I3(n7882), .I4(n7883), .O(n7884));
  LUT3 #(.INIT(8'h96)) lut_n7885 (.I0(n7871), .I1(n7874), .I2(n7875), .O(n7885));
  LUT3 #(.INIT(8'hE8)) lut_n7886 (.I0(n7881), .I1(n7884), .I2(n7885), .O(n7886));
  LUT3 #(.INIT(8'h96)) lut_n7887 (.I0(x2916), .I1(x2917), .I2(x2918), .O(n7887));
  LUT5 #(.INIT(32'h96696996)) lut_n7888 (.I0(x2907), .I1(x2908), .I2(x2909), .I3(n7882), .I4(n7883), .O(n7888));
  LUT5 #(.INIT(32'hFF969600)) lut_n7889 (.I0(x2913), .I1(x2914), .I2(x2915), .I3(n7887), .I4(n7888), .O(n7889));
  LUT3 #(.INIT(8'h96)) lut_n7890 (.I0(x2922), .I1(x2923), .I2(x2924), .O(n7890));
  LUT5 #(.INIT(32'h96696996)) lut_n7891 (.I0(x2913), .I1(x2914), .I2(x2915), .I3(n7887), .I4(n7888), .O(n7891));
  LUT5 #(.INIT(32'hFF969600)) lut_n7892 (.I0(x2919), .I1(x2920), .I2(x2921), .I3(n7890), .I4(n7891), .O(n7892));
  LUT3 #(.INIT(8'h96)) lut_n7893 (.I0(n7881), .I1(n7884), .I2(n7885), .O(n7893));
  LUT3 #(.INIT(8'hE8)) lut_n7894 (.I0(n7889), .I1(n7892), .I2(n7893), .O(n7894));
  LUT3 #(.INIT(8'h96)) lut_n7895 (.I0(n7868), .I1(n7876), .I2(n7877), .O(n7895));
  LUT3 #(.INIT(8'hE8)) lut_n7896 (.I0(n7886), .I1(n7894), .I2(n7895), .O(n7896));
  LUT3 #(.INIT(8'h96)) lut_n7897 (.I0(n7840), .I1(n7858), .I2(n7859), .O(n7897));
  LUT3 #(.INIT(8'hE8)) lut_n7898 (.I0(n7878), .I1(n7896), .I2(n7897), .O(n7898));
  LUT3 #(.INIT(8'h96)) lut_n7899 (.I0(n7778), .I1(n7816), .I2(n7817), .O(n7899));
  LUT3 #(.INIT(8'hE8)) lut_n7900 (.I0(n7860), .I1(n7898), .I2(n7899), .O(n7900));
  LUT3 #(.INIT(8'h96)) lut_n7901 (.I0(x2928), .I1(x2929), .I2(x2930), .O(n7901));
  LUT5 #(.INIT(32'h96696996)) lut_n7902 (.I0(x2919), .I1(x2920), .I2(x2921), .I3(n7890), .I4(n7891), .O(n7902));
  LUT5 #(.INIT(32'hFF969600)) lut_n7903 (.I0(x2925), .I1(x2926), .I2(x2927), .I3(n7901), .I4(n7902), .O(n7903));
  LUT3 #(.INIT(8'h96)) lut_n7904 (.I0(x2934), .I1(x2935), .I2(x2936), .O(n7904));
  LUT5 #(.INIT(32'h96696996)) lut_n7905 (.I0(x2925), .I1(x2926), .I2(x2927), .I3(n7901), .I4(n7902), .O(n7905));
  LUT5 #(.INIT(32'hFF969600)) lut_n7906 (.I0(x2931), .I1(x2932), .I2(x2933), .I3(n7904), .I4(n7905), .O(n7906));
  LUT3 #(.INIT(8'h96)) lut_n7907 (.I0(n7889), .I1(n7892), .I2(n7893), .O(n7907));
  LUT3 #(.INIT(8'hE8)) lut_n7908 (.I0(n7903), .I1(n7906), .I2(n7907), .O(n7908));
  LUT3 #(.INIT(8'h96)) lut_n7909 (.I0(x2940), .I1(x2941), .I2(x2942), .O(n7909));
  LUT5 #(.INIT(32'h96696996)) lut_n7910 (.I0(x2931), .I1(x2932), .I2(x2933), .I3(n7904), .I4(n7905), .O(n7910));
  LUT5 #(.INIT(32'hFF969600)) lut_n7911 (.I0(x2937), .I1(x2938), .I2(x2939), .I3(n7909), .I4(n7910), .O(n7911));
  LUT3 #(.INIT(8'h96)) lut_n7912 (.I0(x2946), .I1(x2947), .I2(x2948), .O(n7912));
  LUT5 #(.INIT(32'h96696996)) lut_n7913 (.I0(x2937), .I1(x2938), .I2(x2939), .I3(n7909), .I4(n7910), .O(n7913));
  LUT5 #(.INIT(32'hFF969600)) lut_n7914 (.I0(x2943), .I1(x2944), .I2(x2945), .I3(n7912), .I4(n7913), .O(n7914));
  LUT3 #(.INIT(8'h96)) lut_n7915 (.I0(n7903), .I1(n7906), .I2(n7907), .O(n7915));
  LUT3 #(.INIT(8'hE8)) lut_n7916 (.I0(n7911), .I1(n7914), .I2(n7915), .O(n7916));
  LUT3 #(.INIT(8'h96)) lut_n7917 (.I0(n7886), .I1(n7894), .I2(n7895), .O(n7917));
  LUT3 #(.INIT(8'hE8)) lut_n7918 (.I0(n7908), .I1(n7916), .I2(n7917), .O(n7918));
  LUT3 #(.INIT(8'h96)) lut_n7919 (.I0(x2952), .I1(x2953), .I2(x2954), .O(n7919));
  LUT5 #(.INIT(32'h96696996)) lut_n7920 (.I0(x2943), .I1(x2944), .I2(x2945), .I3(n7912), .I4(n7913), .O(n7920));
  LUT5 #(.INIT(32'hFF969600)) lut_n7921 (.I0(x2949), .I1(x2950), .I2(x2951), .I3(n7919), .I4(n7920), .O(n7921));
  LUT3 #(.INIT(8'h96)) lut_n7922 (.I0(x2958), .I1(x2959), .I2(x2960), .O(n7922));
  LUT5 #(.INIT(32'h96696996)) lut_n7923 (.I0(x2949), .I1(x2950), .I2(x2951), .I3(n7919), .I4(n7920), .O(n7923));
  LUT5 #(.INIT(32'hFF969600)) lut_n7924 (.I0(x2955), .I1(x2956), .I2(x2957), .I3(n7922), .I4(n7923), .O(n7924));
  LUT3 #(.INIT(8'h96)) lut_n7925 (.I0(n7911), .I1(n7914), .I2(n7915), .O(n7925));
  LUT3 #(.INIT(8'hE8)) lut_n7926 (.I0(n7921), .I1(n7924), .I2(n7925), .O(n7926));
  LUT3 #(.INIT(8'h96)) lut_n7927 (.I0(x2964), .I1(x2965), .I2(x2966), .O(n7927));
  LUT5 #(.INIT(32'h96696996)) lut_n7928 (.I0(x2955), .I1(x2956), .I2(x2957), .I3(n7922), .I4(n7923), .O(n7928));
  LUT5 #(.INIT(32'hFF969600)) lut_n7929 (.I0(x2961), .I1(x2962), .I2(x2963), .I3(n7927), .I4(n7928), .O(n7929));
  LUT3 #(.INIT(8'h96)) lut_n7930 (.I0(x2970), .I1(x2971), .I2(x2972), .O(n7930));
  LUT5 #(.INIT(32'h96696996)) lut_n7931 (.I0(x2961), .I1(x2962), .I2(x2963), .I3(n7927), .I4(n7928), .O(n7931));
  LUT5 #(.INIT(32'hFF969600)) lut_n7932 (.I0(x2967), .I1(x2968), .I2(x2969), .I3(n7930), .I4(n7931), .O(n7932));
  LUT3 #(.INIT(8'h96)) lut_n7933 (.I0(n7921), .I1(n7924), .I2(n7925), .O(n7933));
  LUT3 #(.INIT(8'hE8)) lut_n7934 (.I0(n7929), .I1(n7932), .I2(n7933), .O(n7934));
  LUT3 #(.INIT(8'h96)) lut_n7935 (.I0(n7908), .I1(n7916), .I2(n7917), .O(n7935));
  LUT3 #(.INIT(8'hE8)) lut_n7936 (.I0(n7926), .I1(n7934), .I2(n7935), .O(n7936));
  LUT3 #(.INIT(8'h96)) lut_n7937 (.I0(n7878), .I1(n7896), .I2(n7897), .O(n7937));
  LUT3 #(.INIT(8'h96)) lut_n7938 (.I0(x2976), .I1(x2977), .I2(x2978), .O(n7938));
  LUT5 #(.INIT(32'h96696996)) lut_n7939 (.I0(x2967), .I1(x2968), .I2(x2969), .I3(n7930), .I4(n7931), .O(n7939));
  LUT5 #(.INIT(32'hFF969600)) lut_n7940 (.I0(x2973), .I1(x2974), .I2(x2975), .I3(n7938), .I4(n7939), .O(n7940));
  LUT3 #(.INIT(8'h96)) lut_n7941 (.I0(x2982), .I1(x2983), .I2(x2984), .O(n7941));
  LUT5 #(.INIT(32'h96696996)) lut_n7942 (.I0(x2973), .I1(x2974), .I2(x2975), .I3(n7938), .I4(n7939), .O(n7942));
  LUT5 #(.INIT(32'hFF969600)) lut_n7943 (.I0(x2979), .I1(x2980), .I2(x2981), .I3(n7941), .I4(n7942), .O(n7943));
  LUT3 #(.INIT(8'h96)) lut_n7944 (.I0(n7929), .I1(n7932), .I2(n7933), .O(n7944));
  LUT3 #(.INIT(8'hE8)) lut_n7945 (.I0(n7940), .I1(n7943), .I2(n7944), .O(n7945));
  LUT3 #(.INIT(8'h96)) lut_n7946 (.I0(x2988), .I1(x2989), .I2(x2990), .O(n7946));
  LUT5 #(.INIT(32'h96696996)) lut_n7947 (.I0(x2979), .I1(x2980), .I2(x2981), .I3(n7941), .I4(n7942), .O(n7947));
  LUT5 #(.INIT(32'hFF969600)) lut_n7948 (.I0(x2985), .I1(x2986), .I2(x2987), .I3(n7946), .I4(n7947), .O(n7948));
  LUT3 #(.INIT(8'h96)) lut_n7949 (.I0(x2994), .I1(x2995), .I2(x2996), .O(n7949));
  LUT5 #(.INIT(32'h96696996)) lut_n7950 (.I0(x2985), .I1(x2986), .I2(x2987), .I3(n7946), .I4(n7947), .O(n7950));
  LUT5 #(.INIT(32'hFF969600)) lut_n7951 (.I0(x2991), .I1(x2992), .I2(x2993), .I3(n7949), .I4(n7950), .O(n7951));
  LUT3 #(.INIT(8'h96)) lut_n7952 (.I0(n7940), .I1(n7943), .I2(n7944), .O(n7952));
  LUT3 #(.INIT(8'hE8)) lut_n7953 (.I0(n7948), .I1(n7951), .I2(n7952), .O(n7953));
  LUT3 #(.INIT(8'h96)) lut_n7954 (.I0(n7926), .I1(n7934), .I2(n7935), .O(n7954));
  LUT3 #(.INIT(8'hE8)) lut_n7955 (.I0(n7945), .I1(n7953), .I2(n7954), .O(n7955));
  LUT5 #(.INIT(32'h96696996)) lut_n7956 (.I0(x2991), .I1(x2992), .I2(x2993), .I3(n7949), .I4(n7950), .O(n7956));
  LUT5 #(.INIT(32'hFF969600)) lut_n7957 (.I0(x2997), .I1(x2998), .I2(x2999), .I3(x3000), .I4(n7956), .O(n7957));
  LUT5 #(.INIT(32'h96696996)) lut_n7958 (.I0(x2997), .I1(x2998), .I2(x2999), .I3(x3000), .I4(n7956), .O(n7958));
  LUT3 #(.INIT(8'h96)) lut_n7959 (.I0(n7948), .I1(n7951), .I2(n7952), .O(n7959));
  LUT6 #(.INIT(64'hFF96969696969600)) lut_n7960 (.I0(n7945), .I1(n7953), .I2(n7954), .I3(n7957), .I4(n7958), .I5(n7959), .O(n7960));
  LUT3 #(.INIT(8'h96)) lut_n7961 (.I0(n7860), .I1(n7898), .I2(n7899), .O(n7961));
  LUT6 #(.INIT(64'hFFFEFEE8E8808000)) lut_n7962 (.I0(n7918), .I1(n7936), .I2(n7937), .I3(n7955), .I4(n7960), .I5(n7961), .O(n7962));
  LUT3 #(.INIT(8'h96)) lut_n7963 (.I0(n7740), .I1(n7818), .I2(n7819), .O(n7963));
  LUT6 #(.INIT(64'hFF96969696969600)) lut_n7964 (.I0(n7662), .I1(n7820), .I2(n7821), .I3(n7900), .I4(n7962), .I5(n7963), .O(n7964));
  LUT5 #(.INIT(32'hFF969600)) lut_n7965 (.I0(n7184), .I1(n7502), .I2(n7503), .I3(n7822), .I4(n7964), .O(n7965));
  LUT5 #(.INIT(32'hFF969600)) lut_n7966 (.I0(n6226), .I1(n6864), .I2(n6865), .I3(n7504), .I4(n7965), .O(n7966));
  LUT5 #(.INIT(32'hFF969600)) lut_n7967 (.I0(n4254), .I1(n4892), .I2(n5587), .I3(n6866), .I4(n7966), .O(n7967));
  LUT5 #(.INIT(32'h96696996)) lut_n7968 (.I0(n4254), .I1(n4892), .I2(n5587), .I3(n6866), .I4(n7966), .O(n7968));
  LUT3 #(.INIT(8'hE8)) lut_n7969 (.I0(n5588), .I1(n7967), .I2(n7968), .O(n7969));
  assign y0 = n7969;
endmodule
