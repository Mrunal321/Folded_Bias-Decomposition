module top (x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, y0);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64;
  output y0;
  wire n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161;
  LUT3 #(.INIT(8'hE8)) lut_n67 (.I0(x0), .I1(x1), .I2(x2), .O(n67));
  LUT3 #(.INIT(8'hE8)) lut_n68 (.I0(x6), .I1(x7), .I2(x8), .O(n68));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n69 (.I0(x3), .I1(x4), .I2(x5), .I3(n67), .I4(n68), .O(n69));
  LUT3 #(.INIT(8'hE8)) lut_n70 (.I0(x12), .I1(x13), .I2(x14), .O(n70));
  LUT5 #(.INIT(32'hE81717E8)) lut_n71 (.I0(x3), .I1(x4), .I2(x5), .I3(n67), .I4(n68), .O(n71));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n72 (.I0(x9), .I1(x10), .I2(x11), .I3(n70), .I4(n71), .O(n72));
  LUT3 #(.INIT(8'hE8)) lut_n73 (.I0(x18), .I1(x19), .I2(x20), .O(n73));
  LUT5 #(.INIT(32'hE81717E8)) lut_n74 (.I0(x9), .I1(x10), .I2(x11), .I3(n70), .I4(n71), .O(n74));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n75 (.I0(x15), .I1(x16), .I2(x17), .I3(n73), .I4(n74), .O(n75));
  LUT3 #(.INIT(8'hE8)) lut_n76 (.I0(n69), .I1(n72), .I2(n75), .O(n76));
  LUT3 #(.INIT(8'hE8)) lut_n77 (.I0(x24), .I1(x25), .I2(x26), .O(n77));
  LUT5 #(.INIT(32'hE81717E8)) lut_n78 (.I0(x15), .I1(x16), .I2(x17), .I3(n73), .I4(n74), .O(n78));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n79 (.I0(x21), .I1(x22), .I2(x23), .I3(n77), .I4(n78), .O(n79));
  LUT3 #(.INIT(8'hE8)) lut_n80 (.I0(x27), .I1(x28), .I2(x29), .O(n80));
  LUT5 #(.INIT(32'hE81717E8)) lut_n81 (.I0(x21), .I1(x22), .I2(x23), .I3(n77), .I4(n78), .O(n81));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n82 (.I0(x30), .I1(x31), .I2(x32), .I3(n80), .I4(n81), .O(n82));
  LUT3 #(.INIT(8'h96)) lut_n83 (.I0(n69), .I1(n72), .I2(n75), .O(n83));
  LUT3 #(.INIT(8'hE8)) lut_n84 (.I0(n79), .I1(n82), .I2(n83), .O(n84));
  LUT3 #(.INIT(8'hE8)) lut_n85 (.I0(x36), .I1(x37), .I2(x38), .O(n85));
  LUT5 #(.INIT(32'hE81717E8)) lut_n86 (.I0(x30), .I1(x31), .I2(x32), .I3(n80), .I4(n81), .O(n86));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n87 (.I0(x33), .I1(x34), .I2(x35), .I3(n85), .I4(n86), .O(n87));
  LUT3 #(.INIT(8'hE8)) lut_n88 (.I0(x42), .I1(x43), .I2(x44), .O(n88));
  LUT5 #(.INIT(32'hE81717E8)) lut_n89 (.I0(x33), .I1(x34), .I2(x35), .I3(n85), .I4(n86), .O(n89));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n90 (.I0(x39), .I1(x40), .I2(x41), .I3(n88), .I4(n89), .O(n90));
  LUT3 #(.INIT(8'h96)) lut_n91 (.I0(n79), .I1(n82), .I2(n83), .O(n91));
  LUT3 #(.INIT(8'hE8)) lut_n92 (.I0(n87), .I1(n90), .I2(n91), .O(n92));
  LUT3 #(.INIT(8'hE8)) lut_n93 (.I0(n76), .I1(n84), .I2(n92), .O(n93));
  LUT3 #(.INIT(8'hE8)) lut_n94 (.I0(x48), .I1(x49), .I2(x50), .O(n94));
  LUT5 #(.INIT(32'hE81717E8)) lut_n95 (.I0(x39), .I1(x40), .I2(x41), .I3(n88), .I4(n89), .O(n95));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n96 (.I0(x45), .I1(x46), .I2(x47), .I3(n94), .I4(n95), .O(n96));
  LUT3 #(.INIT(8'hE8)) lut_n97 (.I0(x54), .I1(x55), .I2(x56), .O(n97));
  LUT5 #(.INIT(32'hE81717E8)) lut_n98 (.I0(x45), .I1(x46), .I2(x47), .I3(n94), .I4(n95), .O(n98));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n99 (.I0(x51), .I1(x52), .I2(x53), .I3(n97), .I4(n98), .O(n99));
  LUT3 #(.INIT(8'h96)) lut_n100 (.I0(n87), .I1(n90), .I2(n91), .O(n100));
  LUT3 #(.INIT(8'hE8)) lut_n101 (.I0(n96), .I1(n99), .I2(n100), .O(n101));
  LUT3 #(.INIT(8'hE8)) lut_n102 (.I0(x60), .I1(x61), .I2(x62), .O(n102));
  LUT5 #(.INIT(32'hE81717E8)) lut_n103 (.I0(x51), .I1(x52), .I2(x53), .I3(n97), .I4(n98), .O(n103));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n104 (.I0(x57), .I1(x58), .I2(x59), .I3(n102), .I4(n103), .O(n104));
  LUT3 #(.INIT(8'h96)) lut_n105 (.I0(x0), .I1(x1), .I2(x2), .O(n105));
  LUT3 #(.INIT(8'h96)) lut_n106 (.I0(x6), .I1(x7), .I2(x8), .O(n106));
  LUT5 #(.INIT(32'hFF969600)) lut_n107 (.I0(x3), .I1(x4), .I2(x5), .I3(n105), .I4(n106), .O(n107));
  LUT3 #(.INIT(8'h96)) lut_n108 (.I0(x12), .I1(x13), .I2(x14), .O(n108));
  LUT5 #(.INIT(32'h96696996)) lut_n109 (.I0(x3), .I1(x4), .I2(x5), .I3(n105), .I4(n106), .O(n109));
  LUT5 #(.INIT(32'hFF969600)) lut_n110 (.I0(x9), .I1(x10), .I2(x11), .I3(n108), .I4(n109), .O(n110));
  LUT5 #(.INIT(32'hE81717E8)) lut_n111 (.I0(x57), .I1(x58), .I2(x59), .I3(n102), .I4(n103), .O(n111));
  LUT3 #(.INIT(8'hE8)) lut_n112 (.I0(n107), .I1(n110), .I2(n111), .O(n112));
  LUT3 #(.INIT(8'h96)) lut_n113 (.I0(n96), .I1(n99), .I2(n100), .O(n113));
  LUT3 #(.INIT(8'hE8)) lut_n114 (.I0(n104), .I1(n112), .I2(n113), .O(n114));
  LUT3 #(.INIT(8'h96)) lut_n115 (.I0(n76), .I1(n84), .I2(n92), .O(n115));
  LUT3 #(.INIT(8'hE8)) lut_n116 (.I0(n101), .I1(n114), .I2(n115), .O(n116));
  LUT3 #(.INIT(8'h96)) lut_n117 (.I0(x18), .I1(x19), .I2(x20), .O(n117));
  LUT5 #(.INIT(32'h96696996)) lut_n118 (.I0(x9), .I1(x10), .I2(x11), .I3(n108), .I4(n109), .O(n118));
  LUT5 #(.INIT(32'hFF969600)) lut_n119 (.I0(x15), .I1(x16), .I2(x17), .I3(n117), .I4(n118), .O(n119));
  LUT3 #(.INIT(8'h96)) lut_n120 (.I0(x24), .I1(x25), .I2(x26), .O(n120));
  LUT5 #(.INIT(32'h96696996)) lut_n121 (.I0(x15), .I1(x16), .I2(x17), .I3(n117), .I4(n118), .O(n121));
  LUT5 #(.INIT(32'hFF969600)) lut_n122 (.I0(x21), .I1(x22), .I2(x23), .I3(n120), .I4(n121), .O(n122));
  LUT3 #(.INIT(8'h96)) lut_n123 (.I0(n107), .I1(n110), .I2(n111), .O(n123));
  LUT3 #(.INIT(8'hE8)) lut_n124 (.I0(n119), .I1(n122), .I2(n123), .O(n124));
  LUT3 #(.INIT(8'h96)) lut_n125 (.I0(x27), .I1(x28), .I2(x29), .O(n125));
  LUT5 #(.INIT(32'h96696996)) lut_n126 (.I0(x21), .I1(x22), .I2(x23), .I3(n120), .I4(n121), .O(n126));
  LUT5 #(.INIT(32'hFF969600)) lut_n127 (.I0(x30), .I1(x31), .I2(x32), .I3(n125), .I4(n126), .O(n127));
  LUT3 #(.INIT(8'h96)) lut_n128 (.I0(x36), .I1(x37), .I2(x38), .O(n128));
  LUT5 #(.INIT(32'h96696996)) lut_n129 (.I0(x30), .I1(x31), .I2(x32), .I3(n125), .I4(n126), .O(n129));
  LUT5 #(.INIT(32'hFF969600)) lut_n130 (.I0(x33), .I1(x34), .I2(x35), .I3(n128), .I4(n129), .O(n130));
  LUT3 #(.INIT(8'h96)) lut_n131 (.I0(n119), .I1(n122), .I2(n123), .O(n131));
  LUT3 #(.INIT(8'hE8)) lut_n132 (.I0(n127), .I1(n130), .I2(n131), .O(n132));
  LUT3 #(.INIT(8'h96)) lut_n133 (.I0(n104), .I1(n112), .I2(n113), .O(n133));
  LUT3 #(.INIT(8'hE8)) lut_n134 (.I0(n124), .I1(n132), .I2(n133), .O(n134));
  LUT3 #(.INIT(8'h96)) lut_n135 (.I0(x42), .I1(x43), .I2(x44), .O(n135));
  LUT5 #(.INIT(32'h96696996)) lut_n136 (.I0(x33), .I1(x34), .I2(x35), .I3(n128), .I4(n129), .O(n136));
  LUT5 #(.INIT(32'hFF969600)) lut_n137 (.I0(x39), .I1(x40), .I2(x41), .I3(n135), .I4(n136), .O(n137));
  LUT3 #(.INIT(8'h96)) lut_n138 (.I0(x48), .I1(x49), .I2(x50), .O(n138));
  LUT5 #(.INIT(32'h96696996)) lut_n139 (.I0(x39), .I1(x40), .I2(x41), .I3(n135), .I4(n136), .O(n139));
  LUT5 #(.INIT(32'hFF969600)) lut_n140 (.I0(x45), .I1(x46), .I2(x47), .I3(n138), .I4(n139), .O(n140));
  LUT3 #(.INIT(8'h96)) lut_n141 (.I0(n127), .I1(n130), .I2(n131), .O(n141));
  LUT3 #(.INIT(8'hE8)) lut_n142 (.I0(n137), .I1(n140), .I2(n141), .O(n142));
  LUT3 #(.INIT(8'h96)) lut_n143 (.I0(x54), .I1(x55), .I2(x56), .O(n143));
  LUT5 #(.INIT(32'h96696996)) lut_n144 (.I0(x45), .I1(x46), .I2(x47), .I3(n138), .I4(n139), .O(n144));
  LUT5 #(.INIT(32'hFF969600)) lut_n145 (.I0(x51), .I1(x52), .I2(x53), .I3(n143), .I4(n144), .O(n145));
  LUT3 #(.INIT(8'h96)) lut_n146 (.I0(x60), .I1(x61), .I2(x62), .O(n146));
  LUT5 #(.INIT(32'h96696996)) lut_n147 (.I0(x51), .I1(x52), .I2(x53), .I3(n143), .I4(n144), .O(n147));
  LUT5 #(.INIT(32'hFF969600)) lut_n148 (.I0(x57), .I1(x58), .I2(x59), .I3(n146), .I4(n147), .O(n148));
  LUT3 #(.INIT(8'h96)) lut_n149 (.I0(n137), .I1(n140), .I2(n141), .O(n149));
  LUT3 #(.INIT(8'hE8)) lut_n150 (.I0(n145), .I1(n148), .I2(n149), .O(n150));
  LUT3 #(.INIT(8'h96)) lut_n151 (.I0(n124), .I1(n132), .I2(n133), .O(n151));
  LUT3 #(.INIT(8'hE8)) lut_n152 (.I0(n142), .I1(n150), .I2(n151), .O(n152));
  LUT3 #(.INIT(8'h96)) lut_n153 (.I0(n101), .I1(n114), .I2(n115), .O(n153));
  LUT3 #(.INIT(8'hE8)) lut_n154 (.I0(n134), .I1(n152), .I2(n153), .O(n154));
  LUT5 #(.INIT(32'h96696996)) lut_n155 (.I0(x57), .I1(x58), .I2(x59), .I3(n146), .I4(n147), .O(n155));
  LUT3 #(.INIT(8'h96)) lut_n156 (.I0(n145), .I1(n148), .I2(n149), .O(n156));
  LUT3 #(.INIT(8'h96)) lut_n157 (.I0(n142), .I1(n150), .I2(n151), .O(n157));
  LUT5 #(.INIT(32'hFFFE8000)) lut_n158 (.I0(x63), .I1(x64), .I2(n155), .I3(n156), .I4(n157), .O(n158));
  LUT5 #(.INIT(32'h80017FFE)) lut_n159 (.I0(x63), .I1(x64), .I2(n155), .I3(n156), .I4(n157), .O(n159));
  LUT3 #(.INIT(8'h96)) lut_n160 (.I0(n134), .I1(n152), .I2(n153), .O(n160));
  LUT6 #(.INIT(64'hFEE8E8E8E8E8E880)) lut_n161 (.I0(n93), .I1(n116), .I2(n154), .I3(n158), .I4(n159), .I5(n160), .O(n161));
  assign y0 = n161;
endmodule
