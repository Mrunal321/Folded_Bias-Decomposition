module top (x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, y0);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18;
  output y0;
  wire n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40;
  LUT3 #(.INIT(8'hE8)) lut_n21 (.I0(x0), .I1(x1), .I2(x2), .O(n21));
  LUT3 #(.INIT(8'hE8)) lut_n22 (.I0(x6), .I1(x7), .I2(x8), .O(n22));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n23 (.I0(x3), .I1(x4), .I2(x5), .I3(n21), .I4(n22), .O(n23));
  LUT3 #(.INIT(8'hE8)) lut_n24 (.I0(x12), .I1(x13), .I2(x14), .O(n24));
  LUT5 #(.INIT(32'hE81717E8)) lut_n25 (.I0(x3), .I1(x4), .I2(x5), .I3(n21), .I4(n22), .O(n25));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n26 (.I0(x9), .I1(x10), .I2(x11), .I3(n24), .I4(n25), .O(n26));
  LUT5 #(.INIT(32'hE81717E8)) lut_n27 (.I0(x9), .I1(x10), .I2(x11), .I3(n24), .I4(n25), .O(n27));
  LUT4 #(.INIT(16'hFFE8)) lut_n28 (.I0(x15), .I1(x16), .I2(x17), .I3(n27), .O(n28));
  LUT3 #(.INIT(8'hE8)) lut_n29 (.I0(n23), .I1(n26), .I2(n28), .O(n29));
  LUT4 #(.INIT(16'h17E8)) lut_n30 (.I0(x15), .I1(x16), .I2(x17), .I3(n27), .O(n30));
  LUT3 #(.INIT(8'h96)) lut_n31 (.I0(x0), .I1(x1), .I2(x2), .O(n31));
  LUT3 #(.INIT(8'h96)) lut_n32 (.I0(x6), .I1(x7), .I2(x8), .O(n32));
  LUT5 #(.INIT(32'hFF969600)) lut_n33 (.I0(x3), .I1(x4), .I2(x5), .I3(n31), .I4(n32), .O(n33));
  LUT3 #(.INIT(8'h96)) lut_n34 (.I0(n23), .I1(n26), .I2(n28), .O(n34));
  LUT3 #(.INIT(8'h96)) lut_n35 (.I0(x12), .I1(x13), .I2(x14), .O(n35));
  LUT5 #(.INIT(32'h96696996)) lut_n36 (.I0(x3), .I1(x4), .I2(x5), .I3(n31), .I4(n32), .O(n36));
  LUT5 #(.INIT(32'hFF969600)) lut_n37 (.I0(x9), .I1(x10), .I2(x11), .I3(n35), .I4(n36), .O(n37));
  LUT5 #(.INIT(32'h96696996)) lut_n38 (.I0(x9), .I1(x10), .I2(x11), .I3(n35), .I4(n36), .O(n38));
  LUT5 #(.INIT(32'hFF969600)) lut_n39 (.I0(x15), .I1(x16), .I2(x17), .I3(x18), .I4(n38), .O(n39));
  LUT6 #(.INIT(64'hBAAAAAA2AAA2AA20)) lut_n40 (.I0(n29), .I1(n30), .I2(n33), .I3(n34), .I4(n37), .I5(n39), .O(n40));
  assign y0 = n40;
endmodule
