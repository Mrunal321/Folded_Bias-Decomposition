module top (x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255, x256, x257, x258, x259, x260, x261, x262, x263, x264, x265, x266, x267, x268, x269, x270, x271, x272, x273, x274, x275, x276, x277, x278, x279, x280, x281, x282, x283, x284, x285, x286, x287, x288, x289, x290, x291, x292, x293, x294, x295, x296, x297, x298, x299, x300, x301, x302, x303, x304, x305, x306, x307, x308, x309, x310, x311, x312, x313, x314, x315, x316, x317, x318, x319, x320, x321, x322, x323, x324, x325, x326, x327, x328, x329, x330, x331, x332, x333, x334, x335, x336, x337, x338, x339, x340, x341, x342, x343, x344, x345, x346, x347, x348, x349, x350, x351, x352, x353, x354, x355, x356, x357, x358, x359, x360, x361, x362, x363, x364, x365, x366, x367, x368, x369, x370, x371, x372, x373, x374, x375, x376, x377, x378, x379, x380, x381, x382, x383, x384, x385, x386, x387, x388, x389, x390, x391, x392, x393, x394, x395, x396, x397, x398, x399, x400, x401, x402, x403, x404, x405, x406, x407, x408, x409, x410, x411, x412, x413, x414, x415, x416, x417, x418, x419, x420, x421, x422, x423, x424, x425, x426, x427, x428, x429, x430, x431, x432, x433, x434, x435, x436, x437, x438, x439, x440, x441, x442, x443, x444, x445, x446, x447, x448, x449, x450, x451, x452, x453, x454, x455, x456, x457, x458, x459, x460, x461, x462, x463, x464, x465, x466, x467, x468, x469, x470, x471, x472, x473, x474, x475, x476, x477, x478, x479, x480, x481, x482, x483, x484, x485, x486, x487, x488, x489, x490, x491, x492, x493, x494, x495, x496, x497, x498, x499, x500, x501, x502, x503, x504, x505, x506, x507, x508, x509, x510, x511, x512, x513, x514, x515, x516, x517, x518, x519, x520, x521, x522, x523, x524, x525, x526, x527, x528, x529, x530, x531, x532, x533, x534, x535, x536, x537, x538, x539, x540, x541, x542, x543, x544, x545, x546, x547, x548, x549, x550, x551, x552, x553, x554, x555, x556, x557, x558, x559, x560, x561, x562, x563, x564, x565, x566, x567, x568, x569, x570, x571, x572, x573, x574, x575, x576, x577, x578, x579, x580, x581, x582, x583, x584, x585, x586, x587, x588, x589, x590, x591, x592, x593, x594, x595, x596, x597, x598, x599, x600, x601, x602, x603, x604, x605, x606, x607, x608, x609, x610, x611, x612, x613, x614, x615, x616, x617, x618, x619, x620, x621, x622, x623, x624, x625, x626, x627, x628, x629, x630, x631, x632, x633, x634, x635, x636, x637, x638, x639, x640, x641, x642, x643, x644, x645, x646, x647, x648, x649, x650, x651, x652, x653, x654, x655, x656, x657, x658, x659, x660, x661, x662, x663, x664, x665, x666, x667, x668, x669, x670, x671, x672, x673, x674, x675, x676, x677, x678, x679, x680, x681, x682, x683, x684, x685, x686, x687, x688, x689, x690, x691, x692, x693, x694, x695, x696, x697, x698, x699, x700, x701, x702, x703, x704, x705, x706, x707, x708, x709, x710, x711, x712, x713, x714, x715, x716, x717, x718, x719, x720, x721, x722, x723, x724, x725, x726, x727, x728, x729, x730, x731, x732, x733, x734, x735, x736, x737, x738, x739, x740, x741, x742, x743, x744, x745, x746, x747, x748, x749, x750, x751, x752, x753, x754, x755, x756, x757, x758, x759, x760, x761, x762, x763, x764, x765, x766, x767, x768, x769, x770, x771, x772, x773, x774, x775, x776, x777, x778, x779, x780, x781, x782, x783, x784, x785, x786, x787, x788, x789, x790, x791, x792, x793, x794, x795, x796, x797, x798, x799, x800, x801, x802, x803, x804, x805, x806, x807, x808, x809, x810, x811, x812, x813, x814, x815, x816, x817, x818, x819, x820, x821, x822, x823, x824, x825, x826, x827, x828, x829, x830, x831, x832, x833, x834, x835, x836, x837, x838, x839, x840, x841, x842, x843, x844, x845, x846, x847, x848, x849, x850, x851, x852, x853, x854, x855, x856, x857, x858, x859, x860, x861, x862, x863, x864, x865, x866, x867, x868, x869, x870, x871, x872, x873, x874, x875, x876, x877, x878, x879, x880, x881, x882, x883, x884, x885, x886, x887, x888, x889, x890, x891, x892, x893, x894, x895, x896, x897, x898, x899, x900, x901, x902, x903, x904, x905, x906, x907, x908, x909, x910, x911, x912, x913, x914, x915, x916, x917, x918, x919, x920, x921, x922, x923, x924, x925, x926, x927, x928, x929, x930, x931, x932, x933, x934, x935, x936, x937, x938, x939, x940, x941, x942, x943, x944, x945, x946, x947, x948, x949, x950, x951, x952, x953, x954, x955, x956, x957, x958, x959, x960, x961, x962, x963, x964, x965, x966, x967, x968, x969, x970, x971, x972, x973, x974, x975, x976, x977, x978, x979, x980, x981, x982, x983, x984, x985, x986, x987, x988, x989, x990, x991, x992, x993, x994, x995, x996, x997, x998, x999, x1000, x1001, x1002, x1003, x1004, x1005, x1006, x1007, x1008, x1009, x1010, x1011, x1012, x1013, x1014, x1015, x1016, x1017, x1018, x1019, x1020, x1021, x1022, x1023, x1024, x1025, x1026, x1027, x1028, x1029, x1030, x1031, x1032, x1033, x1034, x1035, x1036, x1037, x1038, x1039, x1040, x1041, x1042, x1043, x1044, x1045, x1046, x1047, x1048, x1049, x1050, x1051, x1052, x1053, x1054, x1055, x1056, x1057, x1058, x1059, x1060, x1061, x1062, x1063, x1064, x1065, x1066, x1067, x1068, x1069, x1070, x1071, x1072, x1073, x1074, x1075, x1076, x1077, x1078, x1079, x1080, x1081, x1082, x1083, x1084, x1085, x1086, x1087, x1088, x1089, x1090, x1091, x1092, x1093, x1094, x1095, x1096, x1097, x1098, x1099, x1100, x1101, x1102, x1103, x1104, x1105, x1106, x1107, x1108, x1109, x1110, x1111, x1112, x1113, x1114, x1115, x1116, x1117, x1118, x1119, x1120, x1121, x1122, x1123, x1124, x1125, x1126, x1127, x1128, x1129, x1130, x1131, x1132, x1133, x1134, x1135, x1136, x1137, x1138, x1139, x1140, x1141, x1142, x1143, x1144, x1145, x1146, x1147, x1148, x1149, x1150, x1151, x1152, x1153, x1154, x1155, x1156, x1157, x1158, x1159, x1160, x1161, x1162, x1163, x1164, x1165, x1166, x1167, x1168, x1169, x1170, x1171, x1172, x1173, x1174, x1175, x1176, x1177, x1178, x1179, x1180, x1181, x1182, x1183, x1184, x1185, x1186, x1187, x1188, x1189, x1190, x1191, x1192, x1193, x1194, x1195, x1196, x1197, x1198, x1199, x1200, x1201, x1202, x1203, x1204, x1205, x1206, x1207, x1208, x1209, x1210, x1211, x1212, x1213, x1214, x1215, x1216, x1217, x1218, x1219, x1220, x1221, x1222, x1223, x1224, x1225, x1226, x1227, x1228, x1229, x1230, x1231, x1232, x1233, x1234, x1235, x1236, x1237, x1238, x1239, x1240, x1241, x1242, x1243, x1244, x1245, x1246, x1247, x1248, x1249, x1250, x1251, x1252, x1253, x1254, x1255, x1256, x1257, x1258, x1259, x1260, x1261, x1262, x1263, x1264, x1265, x1266, x1267, x1268, x1269, x1270, x1271, x1272, x1273, x1274, x1275, x1276, x1277, x1278, x1279, x1280, x1281, x1282, x1283, x1284, x1285, x1286, x1287, x1288, x1289, x1290, x1291, x1292, x1293, x1294, x1295, x1296, x1297, x1298, x1299, x1300, x1301, x1302, x1303, x1304, x1305, x1306, x1307, x1308, x1309, x1310, x1311, x1312, x1313, x1314, x1315, x1316, x1317, x1318, x1319, x1320, x1321, x1322, x1323, x1324, x1325, x1326, x1327, x1328, x1329, x1330, x1331, x1332, x1333, x1334, x1335, x1336, x1337, x1338, x1339, x1340, x1341, x1342, x1343, x1344, x1345, x1346, x1347, x1348, x1349, x1350, x1351, x1352, x1353, x1354, x1355, x1356, x1357, x1358, x1359, x1360, x1361, x1362, x1363, x1364, x1365, x1366, x1367, x1368, x1369, x1370, x1371, x1372, x1373, x1374, x1375, x1376, x1377, x1378, x1379, x1380, x1381, x1382, x1383, x1384, x1385, x1386, x1387, x1388, x1389, x1390, x1391, x1392, x1393, x1394, x1395, x1396, x1397, x1398, x1399, x1400, x1401, x1402, x1403, x1404, x1405, x1406, x1407, x1408, x1409, x1410, x1411, x1412, x1413, x1414, x1415, x1416, x1417, x1418, x1419, x1420, x1421, x1422, x1423, x1424, x1425, x1426, x1427, x1428, x1429, x1430, x1431, x1432, x1433, x1434, x1435, x1436, x1437, x1438, x1439, x1440, x1441, x1442, x1443, x1444, x1445, x1446, x1447, x1448, x1449, x1450, x1451, x1452, x1453, x1454, x1455, x1456, x1457, x1458, x1459, x1460, x1461, x1462, x1463, x1464, x1465, x1466, x1467, x1468, x1469, x1470, x1471, x1472, x1473, x1474, x1475, x1476, x1477, x1478, x1479, x1480, x1481, x1482, x1483, x1484, x1485, x1486, x1487, x1488, x1489, x1490, x1491, x1492, x1493, x1494, x1495, x1496, x1497, x1498, x1499, x1500, x1501, x1502, x1503, x1504, x1505, x1506, x1507, x1508, x1509, x1510, x1511, x1512, x1513, x1514, x1515, x1516, x1517, x1518, x1519, x1520, x1521, x1522, x1523, x1524, x1525, x1526, x1527, x1528, x1529, x1530, x1531, x1532, x1533, x1534, x1535, x1536, x1537, x1538, x1539, x1540, x1541, x1542, x1543, x1544, x1545, x1546, x1547, x1548, x1549, x1550, x1551, x1552, x1553, x1554, x1555, x1556, x1557, x1558, x1559, x1560, x1561, x1562, x1563, x1564, x1565, x1566, x1567, x1568, x1569, x1570, x1571, x1572, x1573, x1574, x1575, x1576, x1577, x1578, x1579, x1580, x1581, x1582, x1583, x1584, x1585, x1586, x1587, x1588, x1589, x1590, x1591, x1592, x1593, x1594, x1595, x1596, x1597, x1598, x1599, x1600, x1601, x1602, x1603, x1604, x1605, x1606, x1607, x1608, x1609, x1610, x1611, x1612, x1613, x1614, x1615, x1616, x1617, x1618, x1619, x1620, x1621, x1622, x1623, x1624, x1625, x1626, x1627, x1628, x1629, x1630, x1631, x1632, x1633, x1634, x1635, x1636, x1637, x1638, x1639, x1640, x1641, x1642, x1643, x1644, x1645, x1646, x1647, x1648, x1649, x1650, x1651, x1652, x1653, x1654, x1655, x1656, x1657, x1658, x1659, x1660, x1661, x1662, x1663, x1664, x1665, x1666, x1667, x1668, x1669, x1670, x1671, x1672, x1673, x1674, x1675, x1676, x1677, x1678, x1679, x1680, x1681, x1682, x1683, x1684, x1685, x1686, x1687, x1688, x1689, x1690, x1691, x1692, x1693, x1694, x1695, x1696, x1697, x1698, x1699, x1700, x1701, x1702, x1703, x1704, x1705, x1706, x1707, x1708, x1709, x1710, x1711, x1712, x1713, x1714, x1715, x1716, x1717, x1718, x1719, x1720, x1721, x1722, x1723, x1724, x1725, x1726, x1727, x1728, x1729, x1730, x1731, x1732, x1733, x1734, x1735, x1736, x1737, x1738, x1739, x1740, x1741, x1742, x1743, x1744, x1745, x1746, x1747, x1748, x1749, x1750, x1751, x1752, x1753, x1754, x1755, x1756, x1757, x1758, x1759, x1760, x1761, x1762, x1763, x1764, x1765, x1766, x1767, x1768, x1769, x1770, x1771, x1772, x1773, x1774, x1775, x1776, x1777, x1778, x1779, x1780, x1781, x1782, x1783, x1784, x1785, x1786, x1787, x1788, x1789, x1790, x1791, x1792, x1793, x1794, x1795, x1796, x1797, x1798, x1799, x1800, x1801, x1802, x1803, x1804, x1805, x1806, x1807, x1808, x1809, x1810, x1811, x1812, x1813, x1814, x1815, x1816, x1817, x1818, x1819, x1820, x1821, x1822, x1823, x1824, x1825, x1826, x1827, x1828, x1829, x1830, x1831, x1832, x1833, x1834, x1835, x1836, x1837, x1838, x1839, x1840, x1841, x1842, x1843, x1844, x1845, x1846, x1847, x1848, x1849, x1850, x1851, x1852, x1853, x1854, x1855, x1856, x1857, x1858, x1859, x1860, x1861, x1862, x1863, x1864, x1865, x1866, x1867, x1868, x1869, x1870, x1871, x1872, x1873, x1874, x1875, x1876, x1877, x1878, x1879, x1880, x1881, x1882, x1883, x1884, x1885, x1886, x1887, x1888, x1889, x1890, x1891, x1892, x1893, x1894, x1895, x1896, x1897, x1898, x1899, x1900, x1901, x1902, x1903, x1904, x1905, x1906, x1907, x1908, x1909, x1910, x1911, x1912, x1913, x1914, x1915, x1916, x1917, x1918, x1919, x1920, x1921, x1922, x1923, x1924, x1925, x1926, x1927, x1928, x1929, x1930, x1931, x1932, x1933, x1934, x1935, x1936, x1937, x1938, x1939, x1940, x1941, x1942, x1943, x1944, x1945, x1946, x1947, x1948, x1949, x1950, x1951, x1952, x1953, x1954, x1955, x1956, x1957, x1958, x1959, x1960, x1961, x1962, x1963, x1964, x1965, x1966, x1967, x1968, x1969, x1970, x1971, x1972, x1973, x1974, x1975, x1976, x1977, x1978, x1979, x1980, x1981, x1982, x1983, x1984, x1985, x1986, x1987, x1988, x1989, x1990, x1991, x1992, x1993, x1994, x1995, x1996, x1997, x1998, x1999, x2000, x2001, x2002, x2003, x2004, x2005, x2006, x2007, x2008, x2009, x2010, x2011, x2012, x2013, x2014, x2015, x2016, x2017, x2018, x2019, x2020, x2021, x2022, x2023, x2024, x2025, x2026, x2027, x2028, x2029, x2030, x2031, x2032, x2033, x2034, x2035, x2036, x2037, x2038, x2039, x2040, x2041, x2042, x2043, x2044, x2045, x2046, x2047, x2048, x2049, x2050, x2051, x2052, x2053, x2054, x2055, x2056, x2057, x2058, x2059, x2060, x2061, x2062, x2063, x2064, x2065, x2066, x2067, x2068, x2069, x2070, x2071, x2072, x2073, x2074, x2075, x2076, x2077, x2078, x2079, x2080, x2081, x2082, x2083, x2084, x2085, x2086, x2087, x2088, x2089, x2090, x2091, x2092, x2093, x2094, x2095, x2096, x2097, x2098, x2099, x2100, x2101, x2102, x2103, x2104, x2105, x2106, x2107, x2108, x2109, x2110, x2111, x2112, x2113, x2114, x2115, x2116, x2117, x2118, x2119, x2120, x2121, x2122, x2123, x2124, x2125, x2126, x2127, x2128, x2129, x2130, x2131, x2132, x2133, x2134, x2135, x2136, x2137, x2138, x2139, x2140, x2141, x2142, x2143, x2144, x2145, x2146, x2147, x2148, x2149, x2150, x2151, x2152, x2153, x2154, x2155, x2156, x2157, x2158, x2159, x2160, x2161, x2162, x2163, x2164, x2165, x2166, x2167, x2168, x2169, x2170, x2171, x2172, x2173, x2174, x2175, x2176, x2177, x2178, x2179, x2180, x2181, x2182, x2183, x2184, x2185, x2186, x2187, x2188, x2189, x2190, x2191, x2192, x2193, x2194, x2195, x2196, x2197, x2198, x2199, x2200, x2201, x2202, x2203, x2204, x2205, x2206, x2207, x2208, x2209, x2210, x2211, x2212, x2213, x2214, x2215, x2216, x2217, x2218, x2219, x2220, x2221, x2222, x2223, x2224, x2225, x2226, x2227, x2228, x2229, x2230, x2231, x2232, x2233, x2234, x2235, x2236, x2237, x2238, x2239, x2240, x2241, x2242, x2243, x2244, x2245, x2246, x2247, x2248, x2249, x2250, x2251, x2252, x2253, x2254, x2255, x2256, x2257, x2258, x2259, x2260, x2261, x2262, x2263, x2264, x2265, x2266, x2267, x2268, x2269, x2270, x2271, x2272, x2273, x2274, x2275, x2276, x2277, x2278, x2279, x2280, x2281, x2282, x2283, x2284, x2285, x2286, x2287, x2288, x2289, x2290, x2291, x2292, x2293, x2294, x2295, x2296, x2297, x2298, x2299, x2300, x2301, x2302, x2303, x2304, x2305, x2306, x2307, x2308, x2309, x2310, x2311, x2312, x2313, x2314, x2315, x2316, x2317, x2318, x2319, x2320, x2321, x2322, x2323, x2324, x2325, x2326, x2327, x2328, x2329, x2330, x2331, x2332, x2333, x2334, x2335, x2336, x2337, x2338, x2339, x2340, x2341, x2342, x2343, x2344, x2345, x2346, x2347, x2348, x2349, x2350, x2351, x2352, x2353, x2354, x2355, x2356, x2357, x2358, x2359, x2360, x2361, x2362, x2363, x2364, x2365, x2366, x2367, x2368, x2369, x2370, x2371, x2372, x2373, x2374, x2375, x2376, x2377, x2378, x2379, x2380, x2381, x2382, x2383, x2384, x2385, x2386, x2387, x2388, x2389, x2390, x2391, x2392, x2393, x2394, x2395, x2396, x2397, x2398, x2399, x2400, x2401, x2402, x2403, x2404, x2405, x2406, x2407, x2408, x2409, x2410, x2411, x2412, x2413, x2414, x2415, x2416, x2417, x2418, x2419, x2420, x2421, x2422, x2423, x2424, x2425, x2426, x2427, x2428, x2429, x2430, x2431, x2432, x2433, x2434, x2435, x2436, x2437, x2438, x2439, x2440, x2441, x2442, x2443, x2444, x2445, x2446, x2447, x2448, x2449, x2450, x2451, x2452, x2453, x2454, x2455, x2456, x2457, x2458, x2459, x2460, x2461, x2462, x2463, x2464, x2465, x2466, x2467, x2468, x2469, x2470, x2471, x2472, x2473, x2474, x2475, x2476, x2477, x2478, x2479, x2480, x2481, x2482, x2483, x2484, x2485, x2486, x2487, x2488, x2489, x2490, x2491, x2492, x2493, x2494, x2495, x2496, x2497, x2498, x2499, x2500, x2501, x2502, x2503, x2504, x2505, x2506, x2507, x2508, x2509, x2510, x2511, x2512, x2513, x2514, x2515, x2516, x2517, x2518, x2519, x2520, x2521, x2522, x2523, x2524, x2525, x2526, x2527, x2528, x2529, x2530, x2531, x2532, x2533, x2534, x2535, x2536, x2537, x2538, x2539, x2540, x2541, x2542, x2543, x2544, x2545, x2546, x2547, x2548, x2549, x2550, x2551, x2552, x2553, x2554, x2555, x2556, x2557, x2558, x2559, x2560, x2561, x2562, x2563, x2564, x2565, x2566, x2567, x2568, x2569, x2570, x2571, x2572, x2573, x2574, x2575, x2576, x2577, x2578, x2579, x2580, x2581, x2582, x2583, x2584, x2585, x2586, x2587, x2588, x2589, x2590, x2591, x2592, x2593, x2594, x2595, x2596, x2597, x2598, x2599, x2600, x2601, x2602, x2603, x2604, x2605, x2606, x2607, x2608, x2609, x2610, x2611, x2612, x2613, x2614, x2615, x2616, x2617, x2618, x2619, x2620, x2621, x2622, x2623, x2624, x2625, x2626, x2627, x2628, x2629, x2630, x2631, x2632, x2633, x2634, x2635, x2636, x2637, x2638, x2639, x2640, x2641, x2642, x2643, x2644, x2645, x2646, x2647, x2648, x2649, x2650, x2651, x2652, x2653, x2654, x2655, x2656, x2657, x2658, x2659, x2660, x2661, x2662, x2663, x2664, x2665, x2666, x2667, x2668, x2669, x2670, x2671, x2672, x2673, x2674, x2675, x2676, x2677, x2678, x2679, x2680, x2681, x2682, x2683, x2684, x2685, x2686, x2687, x2688, x2689, x2690, x2691, x2692, x2693, x2694, x2695, x2696, x2697, x2698, x2699, x2700, x2701, x2702, x2703, x2704, x2705, x2706, x2707, x2708, x2709, x2710, x2711, x2712, x2713, x2714, x2715, x2716, x2717, x2718, x2719, x2720, x2721, x2722, x2723, x2724, x2725, x2726, x2727, x2728, x2729, x2730, x2731, x2732, x2733, x2734, x2735, x2736, x2737, x2738, x2739, x2740, x2741, x2742, x2743, x2744, x2745, x2746, x2747, x2748, x2749, x2750, x2751, x2752, x2753, x2754, x2755, x2756, x2757, x2758, x2759, x2760, x2761, x2762, x2763, x2764, x2765, x2766, x2767, x2768, x2769, x2770, x2771, x2772, x2773, x2774, x2775, x2776, x2777, x2778, x2779, x2780, x2781, x2782, x2783, x2784, x2785, x2786, x2787, x2788, x2789, x2790, x2791, x2792, x2793, x2794, x2795, x2796, x2797, x2798, x2799, x2800, x2801, x2802, x2803, x2804, x2805, x2806, x2807, x2808, x2809, x2810, x2811, x2812, x2813, x2814, x2815, x2816, x2817, x2818, x2819, x2820, x2821, x2822, x2823, x2824, x2825, x2826, x2827, x2828, x2829, x2830, x2831, x2832, x2833, x2834, x2835, x2836, x2837, x2838, x2839, x2840, x2841, x2842, x2843, x2844, x2845, x2846, x2847, x2848, x2849, x2850, x2851, x2852, x2853, x2854, x2855, x2856, x2857, x2858, x2859, x2860, x2861, x2862, x2863, x2864, x2865, x2866, x2867, x2868, x2869, x2870, x2871, x2872, x2873, x2874, x2875, x2876, x2877, x2878, x2879, x2880, x2881, x2882, x2883, x2884, x2885, x2886, x2887, x2888, x2889, x2890, x2891, x2892, x2893, x2894, x2895, x2896, x2897, x2898, x2899, x2900, x2901, x2902, x2903, x2904, x2905, x2906, x2907, x2908, x2909, x2910, x2911, x2912, x2913, x2914, x2915, x2916, x2917, x2918, x2919, x2920, x2921, x2922, x2923, x2924, x2925, x2926, x2927, x2928, x2929, x2930, x2931, x2932, x2933, x2934, x2935, x2936, x2937, x2938, x2939, x2940, x2941, x2942, x2943, x2944, x2945, x2946, x2947, x2948, x2949, x2950, x2951, x2952, x2953, x2954, x2955, x2956, x2957, x2958, x2959, x2960, x2961, x2962, x2963, x2964, x2965, x2966, x2967, x2968, x2969, x2970, x2971, x2972, x2973, x2974, x2975, x2976, x2977, x2978, x2979, x2980, x2981, x2982, x2983, x2984, x2985, x2986, x2987, x2988, x2989, x2990, x2991, x2992, x2993, x2994, x2995, x2996, x2997, x2998, x2999, x3000, x3001, x3002, x3003, x3004, x3005, x3006, x3007, x3008, x3009, x3010, x3011, x3012, x3013, x3014, x3015, x3016, x3017, x3018, x3019, x3020, x3021, x3022, x3023, x3024, x3025, x3026, x3027, x3028, x3029, x3030, x3031, x3032, x3033, x3034, x3035, x3036, x3037, x3038, x3039, x3040, x3041, x3042, x3043, x3044, x3045, x3046, x3047, x3048, x3049, x3050, x3051, x3052, x3053, x3054, x3055, x3056, x3057, x3058, x3059, x3060, x3061, x3062, x3063, x3064, x3065, x3066, x3067, x3068, x3069, x3070, x3071, x3072, x3073, x3074, x3075, x3076, x3077, x3078, x3079, x3080, x3081, x3082, x3083, x3084, x3085, x3086, x3087, x3088, x3089, x3090, x3091, x3092, x3093, x3094, x3095, x3096, x3097, x3098, x3099, x3100, x3101, x3102, x3103, x3104, x3105, x3106, x3107, x3108, x3109, x3110, x3111, x3112, x3113, x3114, x3115, x3116, x3117, x3118, x3119, x3120, x3121, x3122, x3123, x3124, x3125, x3126, x3127, x3128, x3129, x3130, x3131, x3132, x3133, x3134, x3135, x3136, x3137, x3138, x3139, x3140, x3141, x3142, x3143, x3144, x3145, x3146, x3147, x3148, x3149, x3150, x3151, x3152, x3153, x3154, x3155, x3156, x3157, x3158, x3159, x3160, x3161, x3162, x3163, x3164, x3165, x3166, x3167, x3168, x3169, x3170, x3171, x3172, x3173, x3174, x3175, x3176, x3177, x3178, x3179, x3180, x3181, x3182, x3183, x3184, x3185, x3186, x3187, x3188, x3189, x3190, x3191, x3192, x3193, x3194, x3195, x3196, x3197, x3198, x3199, x3200, x3201, x3202, x3203, x3204, x3205, x3206, x3207, x3208, x3209, x3210, x3211, x3212, x3213, x3214, x3215, x3216, x3217, x3218, x3219, x3220, x3221, x3222, x3223, x3224, x3225, x3226, x3227, x3228, x3229, x3230, x3231, x3232, x3233, x3234, x3235, x3236, x3237, x3238, x3239, x3240, x3241, x3242, x3243, x3244, x3245, x3246, x3247, x3248, x3249, x3250, x3251, x3252, x3253, x3254, x3255, x3256, x3257, x3258, x3259, x3260, x3261, x3262, x3263, x3264, x3265, x3266, x3267, x3268, x3269, x3270, x3271, x3272, x3273, x3274, x3275, x3276, x3277, x3278, x3279, x3280, x3281, x3282, x3283, x3284, x3285, x3286, x3287, x3288, x3289, x3290, x3291, x3292, x3293, x3294, x3295, x3296, x3297, x3298, x3299, x3300, x3301, x3302, x3303, x3304, x3305, x3306, x3307, x3308, x3309, x3310, x3311, x3312, x3313, x3314, x3315, x3316, x3317, x3318, x3319, x3320, x3321, x3322, x3323, x3324, x3325, x3326, x3327, x3328, x3329, x3330, x3331, x3332, x3333, x3334, x3335, x3336, x3337, x3338, x3339, x3340, x3341, x3342, x3343, x3344, x3345, x3346, x3347, x3348, x3349, x3350, x3351, x3352, x3353, x3354, x3355, x3356, x3357, x3358, x3359, x3360, x3361, x3362, x3363, x3364, x3365, x3366, x3367, x3368, x3369, x3370, x3371, x3372, x3373, x3374, x3375, x3376, x3377, x3378, x3379, x3380, x3381, x3382, x3383, x3384, x3385, x3386, x3387, x3388, x3389, x3390, x3391, x3392, x3393, x3394, x3395, x3396, x3397, x3398, x3399, x3400, x3401, x3402, x3403, x3404, x3405, x3406, x3407, x3408, x3409, x3410, x3411, x3412, x3413, x3414, x3415, x3416, x3417, x3418, x3419, x3420, x3421, x3422, x3423, x3424, x3425, x3426, x3427, x3428, x3429, x3430, x3431, x3432, x3433, x3434, x3435, x3436, x3437, x3438, x3439, x3440, x3441, x3442, x3443, x3444, x3445, x3446, x3447, x3448, x3449, x3450, x3451, x3452, x3453, x3454, x3455, x3456, x3457, x3458, x3459, x3460, x3461, x3462, x3463, x3464, x3465, x3466, x3467, x3468, x3469, x3470, x3471, x3472, x3473, x3474, x3475, x3476, x3477, x3478, x3479, x3480, x3481, x3482, x3483, x3484, x3485, x3486, x3487, x3488, x3489, x3490, x3491, x3492, x3493, x3494, x3495, x3496, x3497, x3498, x3499, x3500, x3501, x3502, x3503, x3504, x3505, x3506, x3507, x3508, x3509, x3510, x3511, x3512, x3513, x3514, x3515, x3516, x3517, x3518, x3519, x3520, x3521, x3522, x3523, x3524, x3525, x3526, x3527, x3528, x3529, x3530, x3531, x3532, x3533, x3534, x3535, x3536, x3537, x3538, x3539, x3540, x3541, x3542, x3543, x3544, x3545, x3546, x3547, x3548, x3549, x3550, x3551, x3552, x3553, x3554, x3555, x3556, x3557, x3558, x3559, x3560, x3561, x3562, x3563, x3564, x3565, x3566, x3567, x3568, x3569, x3570, x3571, x3572, x3573, x3574, x3575, x3576, x3577, x3578, x3579, x3580, x3581, x3582, x3583, x3584, x3585, x3586, x3587, x3588, x3589, x3590, x3591, x3592, x3593, x3594, x3595, x3596, x3597, x3598, x3599, x3600, x3601, x3602, x3603, x3604, x3605, x3606, x3607, x3608, x3609, x3610, x3611, x3612, x3613, x3614, x3615, x3616, x3617, x3618, x3619, x3620, x3621, x3622, x3623, x3624, x3625, x3626, x3627, x3628, x3629, x3630, x3631, x3632, x3633, x3634, x3635, x3636, x3637, x3638, x3639, x3640, x3641, x3642, x3643, x3644, x3645, x3646, x3647, x3648, x3649, x3650, x3651, x3652, x3653, x3654, x3655, x3656, x3657, x3658, x3659, x3660, x3661, x3662, x3663, x3664, x3665, x3666, x3667, x3668, x3669, x3670, x3671, x3672, x3673, x3674, x3675, x3676, x3677, x3678, x3679, x3680, x3681, x3682, x3683, x3684, x3685, x3686, x3687, x3688, x3689, x3690, x3691, x3692, x3693, x3694, x3695, x3696, x3697, x3698, x3699, x3700, x3701, x3702, x3703, x3704, x3705, x3706, x3707, x3708, x3709, x3710, x3711, x3712, x3713, x3714, x3715, x3716, x3717, x3718, x3719, x3720, x3721, x3722, x3723, x3724, x3725, x3726, x3727, x3728, x3729, x3730, x3731, x3732, x3733, x3734, x3735, x3736, x3737, x3738, x3739, x3740, x3741, x3742, x3743, x3744, x3745, x3746, x3747, x3748, x3749, x3750, x3751, x3752, x3753, x3754, x3755, x3756, x3757, x3758, x3759, x3760, x3761, x3762, x3763, x3764, x3765, x3766, x3767, x3768, x3769, x3770, x3771, x3772, x3773, x3774, x3775, x3776, x3777, x3778, x3779, x3780, x3781, x3782, x3783, x3784, x3785, x3786, x3787, x3788, x3789, x3790, x3791, x3792, x3793, x3794, x3795, x3796, x3797, x3798, x3799, x3800, x3801, x3802, x3803, x3804, x3805, x3806, x3807, x3808, x3809, x3810, x3811, x3812, x3813, x3814, x3815, x3816, x3817, x3818, x3819, x3820, x3821, x3822, x3823, x3824, x3825, x3826, x3827, x3828, x3829, x3830, x3831, x3832, x3833, x3834, x3835, x3836, x3837, x3838, x3839, x3840, x3841, x3842, x3843, x3844, x3845, x3846, x3847, x3848, x3849, x3850, x3851, x3852, x3853, x3854, x3855, x3856, x3857, x3858, x3859, x3860, x3861, x3862, x3863, x3864, x3865, x3866, x3867, x3868, x3869, x3870, x3871, x3872, x3873, x3874, x3875, x3876, x3877, x3878, x3879, x3880, x3881, x3882, x3883, x3884, x3885, x3886, x3887, x3888, x3889, x3890, x3891, x3892, x3893, x3894, x3895, x3896, x3897, x3898, x3899, x3900, x3901, x3902, x3903, x3904, x3905, x3906, x3907, x3908, x3909, x3910, x3911, x3912, x3913, x3914, x3915, x3916, x3917, x3918, x3919, x3920, x3921, x3922, x3923, x3924, x3925, x3926, x3927, x3928, x3929, x3930, x3931, x3932, x3933, x3934, x3935, x3936, x3937, x3938, x3939, x3940, x3941, x3942, x3943, x3944, x3945, x3946, x3947, x3948, x3949, x3950, x3951, x3952, x3953, x3954, x3955, x3956, x3957, x3958, x3959, x3960, x3961, x3962, x3963, x3964, x3965, x3966, x3967, x3968, x3969, x3970, x3971, x3972, x3973, x3974, x3975, x3976, x3977, x3978, x3979, x3980, x3981, x3982, x3983, x3984, x3985, x3986, x3987, x3988, x3989, x3990, x3991, x3992, x3993, x3994, x3995, x3996, x3997, x3998, x3999, x4000, x4001, x4002, x4003, x4004, x4005, x4006, x4007, x4008, x4009, x4010, x4011, x4012, x4013, x4014, x4015, x4016, x4017, x4018, x4019, x4020, x4021, x4022, x4023, x4024, x4025, x4026, x4027, x4028, x4029, x4030, x4031, x4032, x4033, x4034, x4035, x4036, x4037, x4038, x4039, x4040, x4041, x4042, x4043, x4044, x4045, x4046, x4047, x4048, x4049, x4050, x4051, x4052, x4053, x4054, x4055, x4056, x4057, x4058, x4059, x4060, x4061, x4062, x4063, x4064, x4065, x4066, x4067, x4068, x4069, x4070, x4071, x4072, x4073, x4074, x4075, x4076, x4077, x4078, x4079, x4080, x4081, x4082, x4083, x4084, x4085, x4086, x4087, x4088, x4089, x4090, x4091, x4092, x4093, x4094, x4095, x4096, x4097, x4098, x4099, x4100, x4101, x4102, x4103, x4104, x4105, x4106, x4107, x4108, x4109, x4110, x4111, x4112, x4113, x4114, x4115, x4116, x4117, x4118, x4119, x4120, x4121, x4122, x4123, x4124, x4125, x4126, x4127, x4128, x4129, x4130, x4131, x4132, x4133, x4134, x4135, x4136, x4137, x4138, x4139, x4140, x4141, x4142, x4143, x4144, x4145, x4146, x4147, x4148, x4149, x4150, x4151, x4152, x4153, x4154, x4155, x4156, x4157, x4158, x4159, x4160, x4161, x4162, x4163, x4164, x4165, x4166, x4167, x4168, x4169, x4170, x4171, x4172, x4173, x4174, x4175, x4176, x4177, x4178, x4179, x4180, x4181, x4182, x4183, x4184, x4185, x4186, x4187, x4188, x4189, x4190, x4191, x4192, x4193, x4194, x4195, x4196, x4197, x4198, x4199, x4200, x4201, x4202, x4203, x4204, x4205, x4206, x4207, x4208, x4209, x4210, x4211, x4212, x4213, x4214, x4215, x4216, x4217, x4218, x4219, x4220, x4221, x4222, x4223, x4224, x4225, x4226, x4227, x4228, x4229, x4230, x4231, x4232, x4233, x4234, x4235, x4236, x4237, x4238, x4239, x4240, x4241, x4242, x4243, x4244, x4245, x4246, x4247, x4248, x4249, x4250, x4251, x4252, x4253, x4254, x4255, x4256, x4257, x4258, x4259, x4260, x4261, x4262, x4263, x4264, x4265, x4266, x4267, x4268, x4269, x4270, x4271, x4272, x4273, x4274, x4275, x4276, x4277, x4278, x4279, x4280, x4281, x4282, x4283, x4284, x4285, x4286, x4287, x4288, x4289, x4290, x4291, x4292, x4293, x4294, x4295, x4296, x4297, x4298, x4299, x4300, x4301, x4302, x4303, x4304, x4305, x4306, x4307, x4308, x4309, x4310, x4311, x4312, x4313, x4314, x4315, x4316, x4317, x4318, x4319, x4320, x4321, x4322, x4323, x4324, x4325, x4326, x4327, x4328, x4329, x4330, x4331, x4332, x4333, x4334, x4335, x4336, x4337, x4338, x4339, x4340, x4341, x4342, x4343, x4344, x4345, x4346, x4347, x4348, x4349, x4350, x4351, x4352, x4353, x4354, x4355, x4356, x4357, x4358, x4359, x4360, x4361, x4362, x4363, x4364, x4365, x4366, x4367, x4368, x4369, x4370, x4371, x4372, x4373, x4374, x4375, x4376, x4377, x4378, x4379, x4380, x4381, x4382, x4383, x4384, x4385, x4386, x4387, x4388, x4389, x4390, x4391, x4392, x4393, x4394, x4395, x4396, x4397, x4398, x4399, x4400, x4401, x4402, x4403, x4404, x4405, x4406, x4407, x4408, x4409, x4410, x4411, x4412, x4413, x4414, x4415, x4416, x4417, x4418, x4419, x4420, x4421, x4422, x4423, x4424, x4425, x4426, x4427, x4428, x4429, x4430, x4431, x4432, x4433, x4434, x4435, x4436, x4437, x4438, x4439, x4440, x4441, x4442, x4443, x4444, x4445, x4446, x4447, x4448, x4449, x4450, x4451, x4452, x4453, x4454, x4455, x4456, x4457, x4458, x4459, x4460, x4461, x4462, x4463, x4464, x4465, x4466, x4467, x4468, x4469, x4470, x4471, x4472, x4473, x4474, x4475, x4476, x4477, x4478, x4479, x4480, x4481, x4482, x4483, x4484, x4485, x4486, x4487, x4488, x4489, x4490, x4491, x4492, x4493, x4494, x4495, x4496, x4497, x4498, x4499, x4500, x4501, x4502, x4503, x4504, x4505, x4506, x4507, x4508, x4509, x4510, x4511, x4512, x4513, x4514, x4515, x4516, x4517, x4518, x4519, x4520, x4521, x4522, x4523, x4524, x4525, x4526, x4527, x4528, x4529, x4530, x4531, x4532, x4533, x4534, x4535, x4536, x4537, x4538, x4539, x4540, x4541, x4542, x4543, x4544, x4545, x4546, x4547, x4548, x4549, x4550, x4551, x4552, x4553, x4554, x4555, x4556, x4557, x4558, x4559, x4560, x4561, x4562, x4563, x4564, x4565, x4566, x4567, x4568, x4569, x4570, x4571, x4572, x4573, x4574, x4575, x4576, x4577, x4578, x4579, x4580, x4581, x4582, x4583, x4584, x4585, x4586, x4587, x4588, x4589, x4590, x4591, x4592, x4593, x4594, x4595, x4596, x4597, x4598, x4599, x4600, x4601, x4602, x4603, x4604, x4605, x4606, x4607, x4608, x4609, x4610, x4611, x4612, x4613, x4614, x4615, x4616, x4617, x4618, x4619, x4620, x4621, x4622, x4623, x4624, x4625, x4626, x4627, x4628, x4629, x4630, x4631, x4632, x4633, x4634, x4635, x4636, x4637, x4638, x4639, x4640, x4641, x4642, x4643, x4644, x4645, x4646, x4647, x4648, x4649, x4650, x4651, x4652, x4653, x4654, x4655, x4656, x4657, x4658, x4659, x4660, x4661, x4662, x4663, x4664, x4665, x4666, x4667, x4668, x4669, x4670, x4671, x4672, x4673, x4674, x4675, x4676, x4677, x4678, x4679, x4680, x4681, x4682, x4683, x4684, x4685, x4686, x4687, x4688, x4689, x4690, x4691, x4692, x4693, x4694, x4695, x4696, x4697, x4698, x4699, x4700, x4701, x4702, x4703, x4704, x4705, x4706, x4707, x4708, x4709, x4710, x4711, x4712, x4713, x4714, x4715, x4716, x4717, x4718, x4719, x4720, x4721, x4722, x4723, x4724, x4725, x4726, x4727, x4728, x4729, x4730, x4731, x4732, x4733, x4734, x4735, x4736, x4737, x4738, x4739, x4740, x4741, x4742, x4743, x4744, x4745, x4746, x4747, x4748, x4749, x4750, x4751, x4752, x4753, x4754, x4755, x4756, x4757, x4758, x4759, x4760, x4761, x4762, x4763, x4764, x4765, x4766, x4767, x4768, x4769, x4770, x4771, x4772, x4773, x4774, x4775, x4776, x4777, x4778, x4779, x4780, x4781, x4782, x4783, x4784, x4785, x4786, x4787, x4788, x4789, x4790, x4791, x4792, x4793, x4794, x4795, x4796, x4797, x4798, x4799, x4800, x4801, x4802, x4803, x4804, x4805, x4806, x4807, x4808, x4809, x4810, x4811, x4812, x4813, x4814, x4815, x4816, x4817, x4818, x4819, x4820, x4821, x4822, x4823, x4824, x4825, x4826, x4827, x4828, x4829, x4830, x4831, x4832, x4833, x4834, x4835, x4836, x4837, x4838, x4839, x4840, x4841, x4842, x4843, x4844, x4845, x4846, x4847, x4848, x4849, x4850, x4851, x4852, x4853, x4854, x4855, x4856, x4857, x4858, x4859, x4860, x4861, x4862, x4863, x4864, x4865, x4866, x4867, x4868, x4869, x4870, x4871, x4872, x4873, x4874, x4875, x4876, x4877, x4878, x4879, x4880, x4881, x4882, x4883, x4884, x4885, x4886, x4887, x4888, x4889, x4890, x4891, x4892, x4893, x4894, x4895, x4896, x4897, x4898, x4899, x4900, x4901, x4902, x4903, x4904, x4905, x4906, x4907, x4908, x4909, x4910, x4911, x4912, x4913, x4914, x4915, x4916, x4917, x4918, x4919, x4920, x4921, x4922, x4923, x4924, x4925, x4926, x4927, x4928, x4929, x4930, x4931, x4932, x4933, x4934, x4935, x4936, x4937, x4938, x4939, x4940, x4941, x4942, x4943, x4944, x4945, x4946, x4947, x4948, x4949, x4950, x4951, x4952, x4953, x4954, x4955, x4956, x4957, x4958, x4959, x4960, x4961, x4962, x4963, x4964, x4965, x4966, x4967, x4968, x4969, x4970, x4971, x4972, x4973, x4974, x4975, x4976, x4977, x4978, x4979, x4980, x4981, x4982, x4983, x4984, x4985, x4986, x4987, x4988, x4989, x4990, x4991, x4992, x4993, x4994, x4995, x4996, x4997, x4998, x4999, x5000, x5001, x5002, x5003, x5004, x5005, x5006, x5007, x5008, x5009, x5010, x5011, x5012, x5013, x5014, x5015, x5016, x5017, x5018, x5019, x5020, x5021, x5022, x5023, x5024, y0);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255, x256, x257, x258, x259, x260, x261, x262, x263, x264, x265, x266, x267, x268, x269, x270, x271, x272, x273, x274, x275, x276, x277, x278, x279, x280, x281, x282, x283, x284, x285, x286, x287, x288, x289, x290, x291, x292, x293, x294, x295, x296, x297, x298, x299, x300, x301, x302, x303, x304, x305, x306, x307, x308, x309, x310, x311, x312, x313, x314, x315, x316, x317, x318, x319, x320, x321, x322, x323, x324, x325, x326, x327, x328, x329, x330, x331, x332, x333, x334, x335, x336, x337, x338, x339, x340, x341, x342, x343, x344, x345, x346, x347, x348, x349, x350, x351, x352, x353, x354, x355, x356, x357, x358, x359, x360, x361, x362, x363, x364, x365, x366, x367, x368, x369, x370, x371, x372, x373, x374, x375, x376, x377, x378, x379, x380, x381, x382, x383, x384, x385, x386, x387, x388, x389, x390, x391, x392, x393, x394, x395, x396, x397, x398, x399, x400, x401, x402, x403, x404, x405, x406, x407, x408, x409, x410, x411, x412, x413, x414, x415, x416, x417, x418, x419, x420, x421, x422, x423, x424, x425, x426, x427, x428, x429, x430, x431, x432, x433, x434, x435, x436, x437, x438, x439, x440, x441, x442, x443, x444, x445, x446, x447, x448, x449, x450, x451, x452, x453, x454, x455, x456, x457, x458, x459, x460, x461, x462, x463, x464, x465, x466, x467, x468, x469, x470, x471, x472, x473, x474, x475, x476, x477, x478, x479, x480, x481, x482, x483, x484, x485, x486, x487, x488, x489, x490, x491, x492, x493, x494, x495, x496, x497, x498, x499, x500, x501, x502, x503, x504, x505, x506, x507, x508, x509, x510, x511, x512, x513, x514, x515, x516, x517, x518, x519, x520, x521, x522, x523, x524, x525, x526, x527, x528, x529, x530, x531, x532, x533, x534, x535, x536, x537, x538, x539, x540, x541, x542, x543, x544, x545, x546, x547, x548, x549, x550, x551, x552, x553, x554, x555, x556, x557, x558, x559, x560, x561, x562, x563, x564, x565, x566, x567, x568, x569, x570, x571, x572, x573, x574, x575, x576, x577, x578, x579, x580, x581, x582, x583, x584, x585, x586, x587, x588, x589, x590, x591, x592, x593, x594, x595, x596, x597, x598, x599, x600, x601, x602, x603, x604, x605, x606, x607, x608, x609, x610, x611, x612, x613, x614, x615, x616, x617, x618, x619, x620, x621, x622, x623, x624, x625, x626, x627, x628, x629, x630, x631, x632, x633, x634, x635, x636, x637, x638, x639, x640, x641, x642, x643, x644, x645, x646, x647, x648, x649, x650, x651, x652, x653, x654, x655, x656, x657, x658, x659, x660, x661, x662, x663, x664, x665, x666, x667, x668, x669, x670, x671, x672, x673, x674, x675, x676, x677, x678, x679, x680, x681, x682, x683, x684, x685, x686, x687, x688, x689, x690, x691, x692, x693, x694, x695, x696, x697, x698, x699, x700, x701, x702, x703, x704, x705, x706, x707, x708, x709, x710, x711, x712, x713, x714, x715, x716, x717, x718, x719, x720, x721, x722, x723, x724, x725, x726, x727, x728, x729, x730, x731, x732, x733, x734, x735, x736, x737, x738, x739, x740, x741, x742, x743, x744, x745, x746, x747, x748, x749, x750, x751, x752, x753, x754, x755, x756, x757, x758, x759, x760, x761, x762, x763, x764, x765, x766, x767, x768, x769, x770, x771, x772, x773, x774, x775, x776, x777, x778, x779, x780, x781, x782, x783, x784, x785, x786, x787, x788, x789, x790, x791, x792, x793, x794, x795, x796, x797, x798, x799, x800, x801, x802, x803, x804, x805, x806, x807, x808, x809, x810, x811, x812, x813, x814, x815, x816, x817, x818, x819, x820, x821, x822, x823, x824, x825, x826, x827, x828, x829, x830, x831, x832, x833, x834, x835, x836, x837, x838, x839, x840, x841, x842, x843, x844, x845, x846, x847, x848, x849, x850, x851, x852, x853, x854, x855, x856, x857, x858, x859, x860, x861, x862, x863, x864, x865, x866, x867, x868, x869, x870, x871, x872, x873, x874, x875, x876, x877, x878, x879, x880, x881, x882, x883, x884, x885, x886, x887, x888, x889, x890, x891, x892, x893, x894, x895, x896, x897, x898, x899, x900, x901, x902, x903, x904, x905, x906, x907, x908, x909, x910, x911, x912, x913, x914, x915, x916, x917, x918, x919, x920, x921, x922, x923, x924, x925, x926, x927, x928, x929, x930, x931, x932, x933, x934, x935, x936, x937, x938, x939, x940, x941, x942, x943, x944, x945, x946, x947, x948, x949, x950, x951, x952, x953, x954, x955, x956, x957, x958, x959, x960, x961, x962, x963, x964, x965, x966, x967, x968, x969, x970, x971, x972, x973, x974, x975, x976, x977, x978, x979, x980, x981, x982, x983, x984, x985, x986, x987, x988, x989, x990, x991, x992, x993, x994, x995, x996, x997, x998, x999, x1000, x1001, x1002, x1003, x1004, x1005, x1006, x1007, x1008, x1009, x1010, x1011, x1012, x1013, x1014, x1015, x1016, x1017, x1018, x1019, x1020, x1021, x1022, x1023, x1024, x1025, x1026, x1027, x1028, x1029, x1030, x1031, x1032, x1033, x1034, x1035, x1036, x1037, x1038, x1039, x1040, x1041, x1042, x1043, x1044, x1045, x1046, x1047, x1048, x1049, x1050, x1051, x1052, x1053, x1054, x1055, x1056, x1057, x1058, x1059, x1060, x1061, x1062, x1063, x1064, x1065, x1066, x1067, x1068, x1069, x1070, x1071, x1072, x1073, x1074, x1075, x1076, x1077, x1078, x1079, x1080, x1081, x1082, x1083, x1084, x1085, x1086, x1087, x1088, x1089, x1090, x1091, x1092, x1093, x1094, x1095, x1096, x1097, x1098, x1099, x1100, x1101, x1102, x1103, x1104, x1105, x1106, x1107, x1108, x1109, x1110, x1111, x1112, x1113, x1114, x1115, x1116, x1117, x1118, x1119, x1120, x1121, x1122, x1123, x1124, x1125, x1126, x1127, x1128, x1129, x1130, x1131, x1132, x1133, x1134, x1135, x1136, x1137, x1138, x1139, x1140, x1141, x1142, x1143, x1144, x1145, x1146, x1147, x1148, x1149, x1150, x1151, x1152, x1153, x1154, x1155, x1156, x1157, x1158, x1159, x1160, x1161, x1162, x1163, x1164, x1165, x1166, x1167, x1168, x1169, x1170, x1171, x1172, x1173, x1174, x1175, x1176, x1177, x1178, x1179, x1180, x1181, x1182, x1183, x1184, x1185, x1186, x1187, x1188, x1189, x1190, x1191, x1192, x1193, x1194, x1195, x1196, x1197, x1198, x1199, x1200, x1201, x1202, x1203, x1204, x1205, x1206, x1207, x1208, x1209, x1210, x1211, x1212, x1213, x1214, x1215, x1216, x1217, x1218, x1219, x1220, x1221, x1222, x1223, x1224, x1225, x1226, x1227, x1228, x1229, x1230, x1231, x1232, x1233, x1234, x1235, x1236, x1237, x1238, x1239, x1240, x1241, x1242, x1243, x1244, x1245, x1246, x1247, x1248, x1249, x1250, x1251, x1252, x1253, x1254, x1255, x1256, x1257, x1258, x1259, x1260, x1261, x1262, x1263, x1264, x1265, x1266, x1267, x1268, x1269, x1270, x1271, x1272, x1273, x1274, x1275, x1276, x1277, x1278, x1279, x1280, x1281, x1282, x1283, x1284, x1285, x1286, x1287, x1288, x1289, x1290, x1291, x1292, x1293, x1294, x1295, x1296, x1297, x1298, x1299, x1300, x1301, x1302, x1303, x1304, x1305, x1306, x1307, x1308, x1309, x1310, x1311, x1312, x1313, x1314, x1315, x1316, x1317, x1318, x1319, x1320, x1321, x1322, x1323, x1324, x1325, x1326, x1327, x1328, x1329, x1330, x1331, x1332, x1333, x1334, x1335, x1336, x1337, x1338, x1339, x1340, x1341, x1342, x1343, x1344, x1345, x1346, x1347, x1348, x1349, x1350, x1351, x1352, x1353, x1354, x1355, x1356, x1357, x1358, x1359, x1360, x1361, x1362, x1363, x1364, x1365, x1366, x1367, x1368, x1369, x1370, x1371, x1372, x1373, x1374, x1375, x1376, x1377, x1378, x1379, x1380, x1381, x1382, x1383, x1384, x1385, x1386, x1387, x1388, x1389, x1390, x1391, x1392, x1393, x1394, x1395, x1396, x1397, x1398, x1399, x1400, x1401, x1402, x1403, x1404, x1405, x1406, x1407, x1408, x1409, x1410, x1411, x1412, x1413, x1414, x1415, x1416, x1417, x1418, x1419, x1420, x1421, x1422, x1423, x1424, x1425, x1426, x1427, x1428, x1429, x1430, x1431, x1432, x1433, x1434, x1435, x1436, x1437, x1438, x1439, x1440, x1441, x1442, x1443, x1444, x1445, x1446, x1447, x1448, x1449, x1450, x1451, x1452, x1453, x1454, x1455, x1456, x1457, x1458, x1459, x1460, x1461, x1462, x1463, x1464, x1465, x1466, x1467, x1468, x1469, x1470, x1471, x1472, x1473, x1474, x1475, x1476, x1477, x1478, x1479, x1480, x1481, x1482, x1483, x1484, x1485, x1486, x1487, x1488, x1489, x1490, x1491, x1492, x1493, x1494, x1495, x1496, x1497, x1498, x1499, x1500, x1501, x1502, x1503, x1504, x1505, x1506, x1507, x1508, x1509, x1510, x1511, x1512, x1513, x1514, x1515, x1516, x1517, x1518, x1519, x1520, x1521, x1522, x1523, x1524, x1525, x1526, x1527, x1528, x1529, x1530, x1531, x1532, x1533, x1534, x1535, x1536, x1537, x1538, x1539, x1540, x1541, x1542, x1543, x1544, x1545, x1546, x1547, x1548, x1549, x1550, x1551, x1552, x1553, x1554, x1555, x1556, x1557, x1558, x1559, x1560, x1561, x1562, x1563, x1564, x1565, x1566, x1567, x1568, x1569, x1570, x1571, x1572, x1573, x1574, x1575, x1576, x1577, x1578, x1579, x1580, x1581, x1582, x1583, x1584, x1585, x1586, x1587, x1588, x1589, x1590, x1591, x1592, x1593, x1594, x1595, x1596, x1597, x1598, x1599, x1600, x1601, x1602, x1603, x1604, x1605, x1606, x1607, x1608, x1609, x1610, x1611, x1612, x1613, x1614, x1615, x1616, x1617, x1618, x1619, x1620, x1621, x1622, x1623, x1624, x1625, x1626, x1627, x1628, x1629, x1630, x1631, x1632, x1633, x1634, x1635, x1636, x1637, x1638, x1639, x1640, x1641, x1642, x1643, x1644, x1645, x1646, x1647, x1648, x1649, x1650, x1651, x1652, x1653, x1654, x1655, x1656, x1657, x1658, x1659, x1660, x1661, x1662, x1663, x1664, x1665, x1666, x1667, x1668, x1669, x1670, x1671, x1672, x1673, x1674, x1675, x1676, x1677, x1678, x1679, x1680, x1681, x1682, x1683, x1684, x1685, x1686, x1687, x1688, x1689, x1690, x1691, x1692, x1693, x1694, x1695, x1696, x1697, x1698, x1699, x1700, x1701, x1702, x1703, x1704, x1705, x1706, x1707, x1708, x1709, x1710, x1711, x1712, x1713, x1714, x1715, x1716, x1717, x1718, x1719, x1720, x1721, x1722, x1723, x1724, x1725, x1726, x1727, x1728, x1729, x1730, x1731, x1732, x1733, x1734, x1735, x1736, x1737, x1738, x1739, x1740, x1741, x1742, x1743, x1744, x1745, x1746, x1747, x1748, x1749, x1750, x1751, x1752, x1753, x1754, x1755, x1756, x1757, x1758, x1759, x1760, x1761, x1762, x1763, x1764, x1765, x1766, x1767, x1768, x1769, x1770, x1771, x1772, x1773, x1774, x1775, x1776, x1777, x1778, x1779, x1780, x1781, x1782, x1783, x1784, x1785, x1786, x1787, x1788, x1789, x1790, x1791, x1792, x1793, x1794, x1795, x1796, x1797, x1798, x1799, x1800, x1801, x1802, x1803, x1804, x1805, x1806, x1807, x1808, x1809, x1810, x1811, x1812, x1813, x1814, x1815, x1816, x1817, x1818, x1819, x1820, x1821, x1822, x1823, x1824, x1825, x1826, x1827, x1828, x1829, x1830, x1831, x1832, x1833, x1834, x1835, x1836, x1837, x1838, x1839, x1840, x1841, x1842, x1843, x1844, x1845, x1846, x1847, x1848, x1849, x1850, x1851, x1852, x1853, x1854, x1855, x1856, x1857, x1858, x1859, x1860, x1861, x1862, x1863, x1864, x1865, x1866, x1867, x1868, x1869, x1870, x1871, x1872, x1873, x1874, x1875, x1876, x1877, x1878, x1879, x1880, x1881, x1882, x1883, x1884, x1885, x1886, x1887, x1888, x1889, x1890, x1891, x1892, x1893, x1894, x1895, x1896, x1897, x1898, x1899, x1900, x1901, x1902, x1903, x1904, x1905, x1906, x1907, x1908, x1909, x1910, x1911, x1912, x1913, x1914, x1915, x1916, x1917, x1918, x1919, x1920, x1921, x1922, x1923, x1924, x1925, x1926, x1927, x1928, x1929, x1930, x1931, x1932, x1933, x1934, x1935, x1936, x1937, x1938, x1939, x1940, x1941, x1942, x1943, x1944, x1945, x1946, x1947, x1948, x1949, x1950, x1951, x1952, x1953, x1954, x1955, x1956, x1957, x1958, x1959, x1960, x1961, x1962, x1963, x1964, x1965, x1966, x1967, x1968, x1969, x1970, x1971, x1972, x1973, x1974, x1975, x1976, x1977, x1978, x1979, x1980, x1981, x1982, x1983, x1984, x1985, x1986, x1987, x1988, x1989, x1990, x1991, x1992, x1993, x1994, x1995, x1996, x1997, x1998, x1999, x2000, x2001, x2002, x2003, x2004, x2005, x2006, x2007, x2008, x2009, x2010, x2011, x2012, x2013, x2014, x2015, x2016, x2017, x2018, x2019, x2020, x2021, x2022, x2023, x2024, x2025, x2026, x2027, x2028, x2029, x2030, x2031, x2032, x2033, x2034, x2035, x2036, x2037, x2038, x2039, x2040, x2041, x2042, x2043, x2044, x2045, x2046, x2047, x2048, x2049, x2050, x2051, x2052, x2053, x2054, x2055, x2056, x2057, x2058, x2059, x2060, x2061, x2062, x2063, x2064, x2065, x2066, x2067, x2068, x2069, x2070, x2071, x2072, x2073, x2074, x2075, x2076, x2077, x2078, x2079, x2080, x2081, x2082, x2083, x2084, x2085, x2086, x2087, x2088, x2089, x2090, x2091, x2092, x2093, x2094, x2095, x2096, x2097, x2098, x2099, x2100, x2101, x2102, x2103, x2104, x2105, x2106, x2107, x2108, x2109, x2110, x2111, x2112, x2113, x2114, x2115, x2116, x2117, x2118, x2119, x2120, x2121, x2122, x2123, x2124, x2125, x2126, x2127, x2128, x2129, x2130, x2131, x2132, x2133, x2134, x2135, x2136, x2137, x2138, x2139, x2140, x2141, x2142, x2143, x2144, x2145, x2146, x2147, x2148, x2149, x2150, x2151, x2152, x2153, x2154, x2155, x2156, x2157, x2158, x2159, x2160, x2161, x2162, x2163, x2164, x2165, x2166, x2167, x2168, x2169, x2170, x2171, x2172, x2173, x2174, x2175, x2176, x2177, x2178, x2179, x2180, x2181, x2182, x2183, x2184, x2185, x2186, x2187, x2188, x2189, x2190, x2191, x2192, x2193, x2194, x2195, x2196, x2197, x2198, x2199, x2200, x2201, x2202, x2203, x2204, x2205, x2206, x2207, x2208, x2209, x2210, x2211, x2212, x2213, x2214, x2215, x2216, x2217, x2218, x2219, x2220, x2221, x2222, x2223, x2224, x2225, x2226, x2227, x2228, x2229, x2230, x2231, x2232, x2233, x2234, x2235, x2236, x2237, x2238, x2239, x2240, x2241, x2242, x2243, x2244, x2245, x2246, x2247, x2248, x2249, x2250, x2251, x2252, x2253, x2254, x2255, x2256, x2257, x2258, x2259, x2260, x2261, x2262, x2263, x2264, x2265, x2266, x2267, x2268, x2269, x2270, x2271, x2272, x2273, x2274, x2275, x2276, x2277, x2278, x2279, x2280, x2281, x2282, x2283, x2284, x2285, x2286, x2287, x2288, x2289, x2290, x2291, x2292, x2293, x2294, x2295, x2296, x2297, x2298, x2299, x2300, x2301, x2302, x2303, x2304, x2305, x2306, x2307, x2308, x2309, x2310, x2311, x2312, x2313, x2314, x2315, x2316, x2317, x2318, x2319, x2320, x2321, x2322, x2323, x2324, x2325, x2326, x2327, x2328, x2329, x2330, x2331, x2332, x2333, x2334, x2335, x2336, x2337, x2338, x2339, x2340, x2341, x2342, x2343, x2344, x2345, x2346, x2347, x2348, x2349, x2350, x2351, x2352, x2353, x2354, x2355, x2356, x2357, x2358, x2359, x2360, x2361, x2362, x2363, x2364, x2365, x2366, x2367, x2368, x2369, x2370, x2371, x2372, x2373, x2374, x2375, x2376, x2377, x2378, x2379, x2380, x2381, x2382, x2383, x2384, x2385, x2386, x2387, x2388, x2389, x2390, x2391, x2392, x2393, x2394, x2395, x2396, x2397, x2398, x2399, x2400, x2401, x2402, x2403, x2404, x2405, x2406, x2407, x2408, x2409, x2410, x2411, x2412, x2413, x2414, x2415, x2416, x2417, x2418, x2419, x2420, x2421, x2422, x2423, x2424, x2425, x2426, x2427, x2428, x2429, x2430, x2431, x2432, x2433, x2434, x2435, x2436, x2437, x2438, x2439, x2440, x2441, x2442, x2443, x2444, x2445, x2446, x2447, x2448, x2449, x2450, x2451, x2452, x2453, x2454, x2455, x2456, x2457, x2458, x2459, x2460, x2461, x2462, x2463, x2464, x2465, x2466, x2467, x2468, x2469, x2470, x2471, x2472, x2473, x2474, x2475, x2476, x2477, x2478, x2479, x2480, x2481, x2482, x2483, x2484, x2485, x2486, x2487, x2488, x2489, x2490, x2491, x2492, x2493, x2494, x2495, x2496, x2497, x2498, x2499, x2500, x2501, x2502, x2503, x2504, x2505, x2506, x2507, x2508, x2509, x2510, x2511, x2512, x2513, x2514, x2515, x2516, x2517, x2518, x2519, x2520, x2521, x2522, x2523, x2524, x2525, x2526, x2527, x2528, x2529, x2530, x2531, x2532, x2533, x2534, x2535, x2536, x2537, x2538, x2539, x2540, x2541, x2542, x2543, x2544, x2545, x2546, x2547, x2548, x2549, x2550, x2551, x2552, x2553, x2554, x2555, x2556, x2557, x2558, x2559, x2560, x2561, x2562, x2563, x2564, x2565, x2566, x2567, x2568, x2569, x2570, x2571, x2572, x2573, x2574, x2575, x2576, x2577, x2578, x2579, x2580, x2581, x2582, x2583, x2584, x2585, x2586, x2587, x2588, x2589, x2590, x2591, x2592, x2593, x2594, x2595, x2596, x2597, x2598, x2599, x2600, x2601, x2602, x2603, x2604, x2605, x2606, x2607, x2608, x2609, x2610, x2611, x2612, x2613, x2614, x2615, x2616, x2617, x2618, x2619, x2620, x2621, x2622, x2623, x2624, x2625, x2626, x2627, x2628, x2629, x2630, x2631, x2632, x2633, x2634, x2635, x2636, x2637, x2638, x2639, x2640, x2641, x2642, x2643, x2644, x2645, x2646, x2647, x2648, x2649, x2650, x2651, x2652, x2653, x2654, x2655, x2656, x2657, x2658, x2659, x2660, x2661, x2662, x2663, x2664, x2665, x2666, x2667, x2668, x2669, x2670, x2671, x2672, x2673, x2674, x2675, x2676, x2677, x2678, x2679, x2680, x2681, x2682, x2683, x2684, x2685, x2686, x2687, x2688, x2689, x2690, x2691, x2692, x2693, x2694, x2695, x2696, x2697, x2698, x2699, x2700, x2701, x2702, x2703, x2704, x2705, x2706, x2707, x2708, x2709, x2710, x2711, x2712, x2713, x2714, x2715, x2716, x2717, x2718, x2719, x2720, x2721, x2722, x2723, x2724, x2725, x2726, x2727, x2728, x2729, x2730, x2731, x2732, x2733, x2734, x2735, x2736, x2737, x2738, x2739, x2740, x2741, x2742, x2743, x2744, x2745, x2746, x2747, x2748, x2749, x2750, x2751, x2752, x2753, x2754, x2755, x2756, x2757, x2758, x2759, x2760, x2761, x2762, x2763, x2764, x2765, x2766, x2767, x2768, x2769, x2770, x2771, x2772, x2773, x2774, x2775, x2776, x2777, x2778, x2779, x2780, x2781, x2782, x2783, x2784, x2785, x2786, x2787, x2788, x2789, x2790, x2791, x2792, x2793, x2794, x2795, x2796, x2797, x2798, x2799, x2800, x2801, x2802, x2803, x2804, x2805, x2806, x2807, x2808, x2809, x2810, x2811, x2812, x2813, x2814, x2815, x2816, x2817, x2818, x2819, x2820, x2821, x2822, x2823, x2824, x2825, x2826, x2827, x2828, x2829, x2830, x2831, x2832, x2833, x2834, x2835, x2836, x2837, x2838, x2839, x2840, x2841, x2842, x2843, x2844, x2845, x2846, x2847, x2848, x2849, x2850, x2851, x2852, x2853, x2854, x2855, x2856, x2857, x2858, x2859, x2860, x2861, x2862, x2863, x2864, x2865, x2866, x2867, x2868, x2869, x2870, x2871, x2872, x2873, x2874, x2875, x2876, x2877, x2878, x2879, x2880, x2881, x2882, x2883, x2884, x2885, x2886, x2887, x2888, x2889, x2890, x2891, x2892, x2893, x2894, x2895, x2896, x2897, x2898, x2899, x2900, x2901, x2902, x2903, x2904, x2905, x2906, x2907, x2908, x2909, x2910, x2911, x2912, x2913, x2914, x2915, x2916, x2917, x2918, x2919, x2920, x2921, x2922, x2923, x2924, x2925, x2926, x2927, x2928, x2929, x2930, x2931, x2932, x2933, x2934, x2935, x2936, x2937, x2938, x2939, x2940, x2941, x2942, x2943, x2944, x2945, x2946, x2947, x2948, x2949, x2950, x2951, x2952, x2953, x2954, x2955, x2956, x2957, x2958, x2959, x2960, x2961, x2962, x2963, x2964, x2965, x2966, x2967, x2968, x2969, x2970, x2971, x2972, x2973, x2974, x2975, x2976, x2977, x2978, x2979, x2980, x2981, x2982, x2983, x2984, x2985, x2986, x2987, x2988, x2989, x2990, x2991, x2992, x2993, x2994, x2995, x2996, x2997, x2998, x2999, x3000, x3001, x3002, x3003, x3004, x3005, x3006, x3007, x3008, x3009, x3010, x3011, x3012, x3013, x3014, x3015, x3016, x3017, x3018, x3019, x3020, x3021, x3022, x3023, x3024, x3025, x3026, x3027, x3028, x3029, x3030, x3031, x3032, x3033, x3034, x3035, x3036, x3037, x3038, x3039, x3040, x3041, x3042, x3043, x3044, x3045, x3046, x3047, x3048, x3049, x3050, x3051, x3052, x3053, x3054, x3055, x3056, x3057, x3058, x3059, x3060, x3061, x3062, x3063, x3064, x3065, x3066, x3067, x3068, x3069, x3070, x3071, x3072, x3073, x3074, x3075, x3076, x3077, x3078, x3079, x3080, x3081, x3082, x3083, x3084, x3085, x3086, x3087, x3088, x3089, x3090, x3091, x3092, x3093, x3094, x3095, x3096, x3097, x3098, x3099, x3100, x3101, x3102, x3103, x3104, x3105, x3106, x3107, x3108, x3109, x3110, x3111, x3112, x3113, x3114, x3115, x3116, x3117, x3118, x3119, x3120, x3121, x3122, x3123, x3124, x3125, x3126, x3127, x3128, x3129, x3130, x3131, x3132, x3133, x3134, x3135, x3136, x3137, x3138, x3139, x3140, x3141, x3142, x3143, x3144, x3145, x3146, x3147, x3148, x3149, x3150, x3151, x3152, x3153, x3154, x3155, x3156, x3157, x3158, x3159, x3160, x3161, x3162, x3163, x3164, x3165, x3166, x3167, x3168, x3169, x3170, x3171, x3172, x3173, x3174, x3175, x3176, x3177, x3178, x3179, x3180, x3181, x3182, x3183, x3184, x3185, x3186, x3187, x3188, x3189, x3190, x3191, x3192, x3193, x3194, x3195, x3196, x3197, x3198, x3199, x3200, x3201, x3202, x3203, x3204, x3205, x3206, x3207, x3208, x3209, x3210, x3211, x3212, x3213, x3214, x3215, x3216, x3217, x3218, x3219, x3220, x3221, x3222, x3223, x3224, x3225, x3226, x3227, x3228, x3229, x3230, x3231, x3232, x3233, x3234, x3235, x3236, x3237, x3238, x3239, x3240, x3241, x3242, x3243, x3244, x3245, x3246, x3247, x3248, x3249, x3250, x3251, x3252, x3253, x3254, x3255, x3256, x3257, x3258, x3259, x3260, x3261, x3262, x3263, x3264, x3265, x3266, x3267, x3268, x3269, x3270, x3271, x3272, x3273, x3274, x3275, x3276, x3277, x3278, x3279, x3280, x3281, x3282, x3283, x3284, x3285, x3286, x3287, x3288, x3289, x3290, x3291, x3292, x3293, x3294, x3295, x3296, x3297, x3298, x3299, x3300, x3301, x3302, x3303, x3304, x3305, x3306, x3307, x3308, x3309, x3310, x3311, x3312, x3313, x3314, x3315, x3316, x3317, x3318, x3319, x3320, x3321, x3322, x3323, x3324, x3325, x3326, x3327, x3328, x3329, x3330, x3331, x3332, x3333, x3334, x3335, x3336, x3337, x3338, x3339, x3340, x3341, x3342, x3343, x3344, x3345, x3346, x3347, x3348, x3349, x3350, x3351, x3352, x3353, x3354, x3355, x3356, x3357, x3358, x3359, x3360, x3361, x3362, x3363, x3364, x3365, x3366, x3367, x3368, x3369, x3370, x3371, x3372, x3373, x3374, x3375, x3376, x3377, x3378, x3379, x3380, x3381, x3382, x3383, x3384, x3385, x3386, x3387, x3388, x3389, x3390, x3391, x3392, x3393, x3394, x3395, x3396, x3397, x3398, x3399, x3400, x3401, x3402, x3403, x3404, x3405, x3406, x3407, x3408, x3409, x3410, x3411, x3412, x3413, x3414, x3415, x3416, x3417, x3418, x3419, x3420, x3421, x3422, x3423, x3424, x3425, x3426, x3427, x3428, x3429, x3430, x3431, x3432, x3433, x3434, x3435, x3436, x3437, x3438, x3439, x3440, x3441, x3442, x3443, x3444, x3445, x3446, x3447, x3448, x3449, x3450, x3451, x3452, x3453, x3454, x3455, x3456, x3457, x3458, x3459, x3460, x3461, x3462, x3463, x3464, x3465, x3466, x3467, x3468, x3469, x3470, x3471, x3472, x3473, x3474, x3475, x3476, x3477, x3478, x3479, x3480, x3481, x3482, x3483, x3484, x3485, x3486, x3487, x3488, x3489, x3490, x3491, x3492, x3493, x3494, x3495, x3496, x3497, x3498, x3499, x3500, x3501, x3502, x3503, x3504, x3505, x3506, x3507, x3508, x3509, x3510, x3511, x3512, x3513, x3514, x3515, x3516, x3517, x3518, x3519, x3520, x3521, x3522, x3523, x3524, x3525, x3526, x3527, x3528, x3529, x3530, x3531, x3532, x3533, x3534, x3535, x3536, x3537, x3538, x3539, x3540, x3541, x3542, x3543, x3544, x3545, x3546, x3547, x3548, x3549, x3550, x3551, x3552, x3553, x3554, x3555, x3556, x3557, x3558, x3559, x3560, x3561, x3562, x3563, x3564, x3565, x3566, x3567, x3568, x3569, x3570, x3571, x3572, x3573, x3574, x3575, x3576, x3577, x3578, x3579, x3580, x3581, x3582, x3583, x3584, x3585, x3586, x3587, x3588, x3589, x3590, x3591, x3592, x3593, x3594, x3595, x3596, x3597, x3598, x3599, x3600, x3601, x3602, x3603, x3604, x3605, x3606, x3607, x3608, x3609, x3610, x3611, x3612, x3613, x3614, x3615, x3616, x3617, x3618, x3619, x3620, x3621, x3622, x3623, x3624, x3625, x3626, x3627, x3628, x3629, x3630, x3631, x3632, x3633, x3634, x3635, x3636, x3637, x3638, x3639, x3640, x3641, x3642, x3643, x3644, x3645, x3646, x3647, x3648, x3649, x3650, x3651, x3652, x3653, x3654, x3655, x3656, x3657, x3658, x3659, x3660, x3661, x3662, x3663, x3664, x3665, x3666, x3667, x3668, x3669, x3670, x3671, x3672, x3673, x3674, x3675, x3676, x3677, x3678, x3679, x3680, x3681, x3682, x3683, x3684, x3685, x3686, x3687, x3688, x3689, x3690, x3691, x3692, x3693, x3694, x3695, x3696, x3697, x3698, x3699, x3700, x3701, x3702, x3703, x3704, x3705, x3706, x3707, x3708, x3709, x3710, x3711, x3712, x3713, x3714, x3715, x3716, x3717, x3718, x3719, x3720, x3721, x3722, x3723, x3724, x3725, x3726, x3727, x3728, x3729, x3730, x3731, x3732, x3733, x3734, x3735, x3736, x3737, x3738, x3739, x3740, x3741, x3742, x3743, x3744, x3745, x3746, x3747, x3748, x3749, x3750, x3751, x3752, x3753, x3754, x3755, x3756, x3757, x3758, x3759, x3760, x3761, x3762, x3763, x3764, x3765, x3766, x3767, x3768, x3769, x3770, x3771, x3772, x3773, x3774, x3775, x3776, x3777, x3778, x3779, x3780, x3781, x3782, x3783, x3784, x3785, x3786, x3787, x3788, x3789, x3790, x3791, x3792, x3793, x3794, x3795, x3796, x3797, x3798, x3799, x3800, x3801, x3802, x3803, x3804, x3805, x3806, x3807, x3808, x3809, x3810, x3811, x3812, x3813, x3814, x3815, x3816, x3817, x3818, x3819, x3820, x3821, x3822, x3823, x3824, x3825, x3826, x3827, x3828, x3829, x3830, x3831, x3832, x3833, x3834, x3835, x3836, x3837, x3838, x3839, x3840, x3841, x3842, x3843, x3844, x3845, x3846, x3847, x3848, x3849, x3850, x3851, x3852, x3853, x3854, x3855, x3856, x3857, x3858, x3859, x3860, x3861, x3862, x3863, x3864, x3865, x3866, x3867, x3868, x3869, x3870, x3871, x3872, x3873, x3874, x3875, x3876, x3877, x3878, x3879, x3880, x3881, x3882, x3883, x3884, x3885, x3886, x3887, x3888, x3889, x3890, x3891, x3892, x3893, x3894, x3895, x3896, x3897, x3898, x3899, x3900, x3901, x3902, x3903, x3904, x3905, x3906, x3907, x3908, x3909, x3910, x3911, x3912, x3913, x3914, x3915, x3916, x3917, x3918, x3919, x3920, x3921, x3922, x3923, x3924, x3925, x3926, x3927, x3928, x3929, x3930, x3931, x3932, x3933, x3934, x3935, x3936, x3937, x3938, x3939, x3940, x3941, x3942, x3943, x3944, x3945, x3946, x3947, x3948, x3949, x3950, x3951, x3952, x3953, x3954, x3955, x3956, x3957, x3958, x3959, x3960, x3961, x3962, x3963, x3964, x3965, x3966, x3967, x3968, x3969, x3970, x3971, x3972, x3973, x3974, x3975, x3976, x3977, x3978, x3979, x3980, x3981, x3982, x3983, x3984, x3985, x3986, x3987, x3988, x3989, x3990, x3991, x3992, x3993, x3994, x3995, x3996, x3997, x3998, x3999, x4000, x4001, x4002, x4003, x4004, x4005, x4006, x4007, x4008, x4009, x4010, x4011, x4012, x4013, x4014, x4015, x4016, x4017, x4018, x4019, x4020, x4021, x4022, x4023, x4024, x4025, x4026, x4027, x4028, x4029, x4030, x4031, x4032, x4033, x4034, x4035, x4036, x4037, x4038, x4039, x4040, x4041, x4042, x4043, x4044, x4045, x4046, x4047, x4048, x4049, x4050, x4051, x4052, x4053, x4054, x4055, x4056, x4057, x4058, x4059, x4060, x4061, x4062, x4063, x4064, x4065, x4066, x4067, x4068, x4069, x4070, x4071, x4072, x4073, x4074, x4075, x4076, x4077, x4078, x4079, x4080, x4081, x4082, x4083, x4084, x4085, x4086, x4087, x4088, x4089, x4090, x4091, x4092, x4093, x4094, x4095, x4096, x4097, x4098, x4099, x4100, x4101, x4102, x4103, x4104, x4105, x4106, x4107, x4108, x4109, x4110, x4111, x4112, x4113, x4114, x4115, x4116, x4117, x4118, x4119, x4120, x4121, x4122, x4123, x4124, x4125, x4126, x4127, x4128, x4129, x4130, x4131, x4132, x4133, x4134, x4135, x4136, x4137, x4138, x4139, x4140, x4141, x4142, x4143, x4144, x4145, x4146, x4147, x4148, x4149, x4150, x4151, x4152, x4153, x4154, x4155, x4156, x4157, x4158, x4159, x4160, x4161, x4162, x4163, x4164, x4165, x4166, x4167, x4168, x4169, x4170, x4171, x4172, x4173, x4174, x4175, x4176, x4177, x4178, x4179, x4180, x4181, x4182, x4183, x4184, x4185, x4186, x4187, x4188, x4189, x4190, x4191, x4192, x4193, x4194, x4195, x4196, x4197, x4198, x4199, x4200, x4201, x4202, x4203, x4204, x4205, x4206, x4207, x4208, x4209, x4210, x4211, x4212, x4213, x4214, x4215, x4216, x4217, x4218, x4219, x4220, x4221, x4222, x4223, x4224, x4225, x4226, x4227, x4228, x4229, x4230, x4231, x4232, x4233, x4234, x4235, x4236, x4237, x4238, x4239, x4240, x4241, x4242, x4243, x4244, x4245, x4246, x4247, x4248, x4249, x4250, x4251, x4252, x4253, x4254, x4255, x4256, x4257, x4258, x4259, x4260, x4261, x4262, x4263, x4264, x4265, x4266, x4267, x4268, x4269, x4270, x4271, x4272, x4273, x4274, x4275, x4276, x4277, x4278, x4279, x4280, x4281, x4282, x4283, x4284, x4285, x4286, x4287, x4288, x4289, x4290, x4291, x4292, x4293, x4294, x4295, x4296, x4297, x4298, x4299, x4300, x4301, x4302, x4303, x4304, x4305, x4306, x4307, x4308, x4309, x4310, x4311, x4312, x4313, x4314, x4315, x4316, x4317, x4318, x4319, x4320, x4321, x4322, x4323, x4324, x4325, x4326, x4327, x4328, x4329, x4330, x4331, x4332, x4333, x4334, x4335, x4336, x4337, x4338, x4339, x4340, x4341, x4342, x4343, x4344, x4345, x4346, x4347, x4348, x4349, x4350, x4351, x4352, x4353, x4354, x4355, x4356, x4357, x4358, x4359, x4360, x4361, x4362, x4363, x4364, x4365, x4366, x4367, x4368, x4369, x4370, x4371, x4372, x4373, x4374, x4375, x4376, x4377, x4378, x4379, x4380, x4381, x4382, x4383, x4384, x4385, x4386, x4387, x4388, x4389, x4390, x4391, x4392, x4393, x4394, x4395, x4396, x4397, x4398, x4399, x4400, x4401, x4402, x4403, x4404, x4405, x4406, x4407, x4408, x4409, x4410, x4411, x4412, x4413, x4414, x4415, x4416, x4417, x4418, x4419, x4420, x4421, x4422, x4423, x4424, x4425, x4426, x4427, x4428, x4429, x4430, x4431, x4432, x4433, x4434, x4435, x4436, x4437, x4438, x4439, x4440, x4441, x4442, x4443, x4444, x4445, x4446, x4447, x4448, x4449, x4450, x4451, x4452, x4453, x4454, x4455, x4456, x4457, x4458, x4459, x4460, x4461, x4462, x4463, x4464, x4465, x4466, x4467, x4468, x4469, x4470, x4471, x4472, x4473, x4474, x4475, x4476, x4477, x4478, x4479, x4480, x4481, x4482, x4483, x4484, x4485, x4486, x4487, x4488, x4489, x4490, x4491, x4492, x4493, x4494, x4495, x4496, x4497, x4498, x4499, x4500, x4501, x4502, x4503, x4504, x4505, x4506, x4507, x4508, x4509, x4510, x4511, x4512, x4513, x4514, x4515, x4516, x4517, x4518, x4519, x4520, x4521, x4522, x4523, x4524, x4525, x4526, x4527, x4528, x4529, x4530, x4531, x4532, x4533, x4534, x4535, x4536, x4537, x4538, x4539, x4540, x4541, x4542, x4543, x4544, x4545, x4546, x4547, x4548, x4549, x4550, x4551, x4552, x4553, x4554, x4555, x4556, x4557, x4558, x4559, x4560, x4561, x4562, x4563, x4564, x4565, x4566, x4567, x4568, x4569, x4570, x4571, x4572, x4573, x4574, x4575, x4576, x4577, x4578, x4579, x4580, x4581, x4582, x4583, x4584, x4585, x4586, x4587, x4588, x4589, x4590, x4591, x4592, x4593, x4594, x4595, x4596, x4597, x4598, x4599, x4600, x4601, x4602, x4603, x4604, x4605, x4606, x4607, x4608, x4609, x4610, x4611, x4612, x4613, x4614, x4615, x4616, x4617, x4618, x4619, x4620, x4621, x4622, x4623, x4624, x4625, x4626, x4627, x4628, x4629, x4630, x4631, x4632, x4633, x4634, x4635, x4636, x4637, x4638, x4639, x4640, x4641, x4642, x4643, x4644, x4645, x4646, x4647, x4648, x4649, x4650, x4651, x4652, x4653, x4654, x4655, x4656, x4657, x4658, x4659, x4660, x4661, x4662, x4663, x4664, x4665, x4666, x4667, x4668, x4669, x4670, x4671, x4672, x4673, x4674, x4675, x4676, x4677, x4678, x4679, x4680, x4681, x4682, x4683, x4684, x4685, x4686, x4687, x4688, x4689, x4690, x4691, x4692, x4693, x4694, x4695, x4696, x4697, x4698, x4699, x4700, x4701, x4702, x4703, x4704, x4705, x4706, x4707, x4708, x4709, x4710, x4711, x4712, x4713, x4714, x4715, x4716, x4717, x4718, x4719, x4720, x4721, x4722, x4723, x4724, x4725, x4726, x4727, x4728, x4729, x4730, x4731, x4732, x4733, x4734, x4735, x4736, x4737, x4738, x4739, x4740, x4741, x4742, x4743, x4744, x4745, x4746, x4747, x4748, x4749, x4750, x4751, x4752, x4753, x4754, x4755, x4756, x4757, x4758, x4759, x4760, x4761, x4762, x4763, x4764, x4765, x4766, x4767, x4768, x4769, x4770, x4771, x4772, x4773, x4774, x4775, x4776, x4777, x4778, x4779, x4780, x4781, x4782, x4783, x4784, x4785, x4786, x4787, x4788, x4789, x4790, x4791, x4792, x4793, x4794, x4795, x4796, x4797, x4798, x4799, x4800, x4801, x4802, x4803, x4804, x4805, x4806, x4807, x4808, x4809, x4810, x4811, x4812, x4813, x4814, x4815, x4816, x4817, x4818, x4819, x4820, x4821, x4822, x4823, x4824, x4825, x4826, x4827, x4828, x4829, x4830, x4831, x4832, x4833, x4834, x4835, x4836, x4837, x4838, x4839, x4840, x4841, x4842, x4843, x4844, x4845, x4846, x4847, x4848, x4849, x4850, x4851, x4852, x4853, x4854, x4855, x4856, x4857, x4858, x4859, x4860, x4861, x4862, x4863, x4864, x4865, x4866, x4867, x4868, x4869, x4870, x4871, x4872, x4873, x4874, x4875, x4876, x4877, x4878, x4879, x4880, x4881, x4882, x4883, x4884, x4885, x4886, x4887, x4888, x4889, x4890, x4891, x4892, x4893, x4894, x4895, x4896, x4897, x4898, x4899, x4900, x4901, x4902, x4903, x4904, x4905, x4906, x4907, x4908, x4909, x4910, x4911, x4912, x4913, x4914, x4915, x4916, x4917, x4918, x4919, x4920, x4921, x4922, x4923, x4924, x4925, x4926, x4927, x4928, x4929, x4930, x4931, x4932, x4933, x4934, x4935, x4936, x4937, x4938, x4939, x4940, x4941, x4942, x4943, x4944, x4945, x4946, x4947, x4948, x4949, x4950, x4951, x4952, x4953, x4954, x4955, x4956, x4957, x4958, x4959, x4960, x4961, x4962, x4963, x4964, x4965, x4966, x4967, x4968, x4969, x4970, x4971, x4972, x4973, x4974, x4975, x4976, x4977, x4978, x4979, x4980, x4981, x4982, x4983, x4984, x4985, x4986, x4987, x4988, x4989, x4990, x4991, x4992, x4993, x4994, x4995, x4996, x4997, x4998, x4999, x5000, x5001, x5002, x5003, x5004, x5005, x5006, x5007, x5008, x5009, x5010, x5011, x5012, x5013, x5014, x5015, x5016, x5017, x5018, x5019, x5020, x5021, x5022, x5023, x5024;
  output y0;
  wire n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371;
  LUT3 #(.INIT(8'hE8)) lut_n5027 (.I0(x0), .I1(x1), .I2(x2), .O(n5027));
  LUT3 #(.INIT(8'hE8)) lut_n5028 (.I0(x6), .I1(x7), .I2(x8), .O(n5028));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5029 (.I0(x3), .I1(x4), .I2(x5), .I3(n5027), .I4(n5028), .O(n5029));
  LUT3 #(.INIT(8'hE8)) lut_n5030 (.I0(x12), .I1(x13), .I2(x14), .O(n5030));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5031 (.I0(x3), .I1(x4), .I2(x5), .I3(n5027), .I4(n5028), .O(n5031));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5032 (.I0(x9), .I1(x10), .I2(x11), .I3(n5030), .I4(n5031), .O(n5032));
  LUT3 #(.INIT(8'hE8)) lut_n5033 (.I0(x18), .I1(x19), .I2(x20), .O(n5033));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5034 (.I0(x9), .I1(x10), .I2(x11), .I3(n5030), .I4(n5031), .O(n5034));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5035 (.I0(x15), .I1(x16), .I2(x17), .I3(n5033), .I4(n5034), .O(n5035));
  LUT3 #(.INIT(8'hE8)) lut_n5036 (.I0(n5029), .I1(n5032), .I2(n5035), .O(n5036));
  LUT3 #(.INIT(8'hE8)) lut_n5037 (.I0(x24), .I1(x25), .I2(x26), .O(n5037));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5038 (.I0(x15), .I1(x16), .I2(x17), .I3(n5033), .I4(n5034), .O(n5038));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5039 (.I0(x21), .I1(x22), .I2(x23), .I3(n5037), .I4(n5038), .O(n5039));
  LUT3 #(.INIT(8'hE8)) lut_n5040 (.I0(x27), .I1(x28), .I2(x29), .O(n5040));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5041 (.I0(x21), .I1(x22), .I2(x23), .I3(n5037), .I4(n5038), .O(n5041));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5042 (.I0(x30), .I1(x31), .I2(x32), .I3(n5040), .I4(n5041), .O(n5042));
  LUT3 #(.INIT(8'h96)) lut_n5043 (.I0(n5029), .I1(n5032), .I2(n5035), .O(n5043));
  LUT3 #(.INIT(8'hE8)) lut_n5044 (.I0(n5039), .I1(n5042), .I2(n5043), .O(n5044));
  LUT3 #(.INIT(8'hE8)) lut_n5045 (.I0(x36), .I1(x37), .I2(x38), .O(n5045));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5046 (.I0(x30), .I1(x31), .I2(x32), .I3(n5040), .I4(n5041), .O(n5046));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5047 (.I0(x33), .I1(x34), .I2(x35), .I3(n5045), .I4(n5046), .O(n5047));
  LUT3 #(.INIT(8'hE8)) lut_n5048 (.I0(x42), .I1(x43), .I2(x44), .O(n5048));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5049 (.I0(x33), .I1(x34), .I2(x35), .I3(n5045), .I4(n5046), .O(n5049));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5050 (.I0(x39), .I1(x40), .I2(x41), .I3(n5048), .I4(n5049), .O(n5050));
  LUT3 #(.INIT(8'h96)) lut_n5051 (.I0(n5039), .I1(n5042), .I2(n5043), .O(n5051));
  LUT3 #(.INIT(8'hE8)) lut_n5052 (.I0(n5047), .I1(n5050), .I2(n5051), .O(n5052));
  LUT3 #(.INIT(8'hE8)) lut_n5053 (.I0(n5036), .I1(n5044), .I2(n5052), .O(n5053));
  LUT3 #(.INIT(8'hE8)) lut_n5054 (.I0(x48), .I1(x49), .I2(x50), .O(n5054));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5055 (.I0(x39), .I1(x40), .I2(x41), .I3(n5048), .I4(n5049), .O(n5055));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5056 (.I0(x45), .I1(x46), .I2(x47), .I3(n5054), .I4(n5055), .O(n5056));
  LUT3 #(.INIT(8'hE8)) lut_n5057 (.I0(x54), .I1(x55), .I2(x56), .O(n5057));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5058 (.I0(x45), .I1(x46), .I2(x47), .I3(n5054), .I4(n5055), .O(n5058));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5059 (.I0(x51), .I1(x52), .I2(x53), .I3(n5057), .I4(n5058), .O(n5059));
  LUT3 #(.INIT(8'h96)) lut_n5060 (.I0(n5047), .I1(n5050), .I2(n5051), .O(n5060));
  LUT3 #(.INIT(8'hE8)) lut_n5061 (.I0(n5056), .I1(n5059), .I2(n5060), .O(n5061));
  LUT3 #(.INIT(8'hE8)) lut_n5062 (.I0(x60), .I1(x61), .I2(x62), .O(n5062));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5063 (.I0(x51), .I1(x52), .I2(x53), .I3(n5057), .I4(n5058), .O(n5063));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5064 (.I0(x57), .I1(x58), .I2(x59), .I3(n5062), .I4(n5063), .O(n5064));
  LUT3 #(.INIT(8'hE8)) lut_n5065 (.I0(x66), .I1(x67), .I2(x68), .O(n5065));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5066 (.I0(x57), .I1(x58), .I2(x59), .I3(n5062), .I4(n5063), .O(n5066));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5067 (.I0(x63), .I1(x64), .I2(x65), .I3(n5065), .I4(n5066), .O(n5067));
  LUT3 #(.INIT(8'h96)) lut_n5068 (.I0(n5056), .I1(n5059), .I2(n5060), .O(n5068));
  LUT3 #(.INIT(8'hE8)) lut_n5069 (.I0(n5064), .I1(n5067), .I2(n5068), .O(n5069));
  LUT3 #(.INIT(8'h96)) lut_n5070 (.I0(n5036), .I1(n5044), .I2(n5052), .O(n5070));
  LUT3 #(.INIT(8'hE8)) lut_n5071 (.I0(n5061), .I1(n5069), .I2(n5070), .O(n5071));
  LUT3 #(.INIT(8'hE8)) lut_n5072 (.I0(x72), .I1(x73), .I2(x74), .O(n5072));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5073 (.I0(x63), .I1(x64), .I2(x65), .I3(n5065), .I4(n5066), .O(n5073));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5074 (.I0(x69), .I1(x70), .I2(x71), .I3(n5072), .I4(n5073), .O(n5074));
  LUT3 #(.INIT(8'hE8)) lut_n5075 (.I0(x78), .I1(x79), .I2(x80), .O(n5075));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5076 (.I0(x69), .I1(x70), .I2(x71), .I3(n5072), .I4(n5073), .O(n5076));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5077 (.I0(x75), .I1(x76), .I2(x77), .I3(n5075), .I4(n5076), .O(n5077));
  LUT3 #(.INIT(8'h96)) lut_n5078 (.I0(n5064), .I1(n5067), .I2(n5068), .O(n5078));
  LUT3 #(.INIT(8'hE8)) lut_n5079 (.I0(n5074), .I1(n5077), .I2(n5078), .O(n5079));
  LUT3 #(.INIT(8'hE8)) lut_n5080 (.I0(x84), .I1(x85), .I2(x86), .O(n5080));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5081 (.I0(x75), .I1(x76), .I2(x77), .I3(n5075), .I4(n5076), .O(n5081));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5082 (.I0(x81), .I1(x82), .I2(x83), .I3(n5080), .I4(n5081), .O(n5082));
  LUT3 #(.INIT(8'hE8)) lut_n5083 (.I0(x90), .I1(x91), .I2(x92), .O(n5083));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5084 (.I0(x81), .I1(x82), .I2(x83), .I3(n5080), .I4(n5081), .O(n5084));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5085 (.I0(x87), .I1(x88), .I2(x89), .I3(n5083), .I4(n5084), .O(n5085));
  LUT3 #(.INIT(8'h96)) lut_n5086 (.I0(n5074), .I1(n5077), .I2(n5078), .O(n5086));
  LUT3 #(.INIT(8'hE8)) lut_n5087 (.I0(n5082), .I1(n5085), .I2(n5086), .O(n5087));
  LUT3 #(.INIT(8'h96)) lut_n5088 (.I0(n5061), .I1(n5069), .I2(n5070), .O(n5088));
  LUT3 #(.INIT(8'hE8)) lut_n5089 (.I0(n5079), .I1(n5087), .I2(n5088), .O(n5089));
  LUT3 #(.INIT(8'hE8)) lut_n5090 (.I0(n5053), .I1(n5071), .I2(n5089), .O(n5090));
  LUT3 #(.INIT(8'hE8)) lut_n5091 (.I0(x96), .I1(x97), .I2(x98), .O(n5091));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5092 (.I0(x87), .I1(x88), .I2(x89), .I3(n5083), .I4(n5084), .O(n5092));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5093 (.I0(x93), .I1(x94), .I2(x95), .I3(n5091), .I4(n5092), .O(n5093));
  LUT3 #(.INIT(8'hE8)) lut_n5094 (.I0(x102), .I1(x103), .I2(x104), .O(n5094));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5095 (.I0(x93), .I1(x94), .I2(x95), .I3(n5091), .I4(n5092), .O(n5095));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5096 (.I0(x99), .I1(x100), .I2(x101), .I3(n5094), .I4(n5095), .O(n5096));
  LUT3 #(.INIT(8'h96)) lut_n5097 (.I0(n5082), .I1(n5085), .I2(n5086), .O(n5097));
  LUT3 #(.INIT(8'hE8)) lut_n5098 (.I0(n5093), .I1(n5096), .I2(n5097), .O(n5098));
  LUT3 #(.INIT(8'hE8)) lut_n5099 (.I0(x108), .I1(x109), .I2(x110), .O(n5099));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5100 (.I0(x99), .I1(x100), .I2(x101), .I3(n5094), .I4(n5095), .O(n5100));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5101 (.I0(x105), .I1(x106), .I2(x107), .I3(n5099), .I4(n5100), .O(n5101));
  LUT3 #(.INIT(8'hE8)) lut_n5102 (.I0(x114), .I1(x115), .I2(x116), .O(n5102));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5103 (.I0(x105), .I1(x106), .I2(x107), .I3(n5099), .I4(n5100), .O(n5103));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5104 (.I0(x111), .I1(x112), .I2(x113), .I3(n5102), .I4(n5103), .O(n5104));
  LUT3 #(.INIT(8'h96)) lut_n5105 (.I0(n5093), .I1(n5096), .I2(n5097), .O(n5105));
  LUT3 #(.INIT(8'hE8)) lut_n5106 (.I0(n5101), .I1(n5104), .I2(n5105), .O(n5106));
  LUT3 #(.INIT(8'h96)) lut_n5107 (.I0(n5079), .I1(n5087), .I2(n5088), .O(n5107));
  LUT3 #(.INIT(8'hE8)) lut_n5108 (.I0(n5098), .I1(n5106), .I2(n5107), .O(n5108));
  LUT3 #(.INIT(8'hE8)) lut_n5109 (.I0(x120), .I1(x121), .I2(x122), .O(n5109));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5110 (.I0(x111), .I1(x112), .I2(x113), .I3(n5102), .I4(n5103), .O(n5110));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5111 (.I0(x117), .I1(x118), .I2(x119), .I3(n5109), .I4(n5110), .O(n5111));
  LUT3 #(.INIT(8'hE8)) lut_n5112 (.I0(x126), .I1(x127), .I2(x128), .O(n5112));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5113 (.I0(x117), .I1(x118), .I2(x119), .I3(n5109), .I4(n5110), .O(n5113));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5114 (.I0(x123), .I1(x124), .I2(x125), .I3(n5112), .I4(n5113), .O(n5114));
  LUT3 #(.INIT(8'h96)) lut_n5115 (.I0(n5101), .I1(n5104), .I2(n5105), .O(n5115));
  LUT3 #(.INIT(8'hE8)) lut_n5116 (.I0(n5111), .I1(n5114), .I2(n5115), .O(n5116));
  LUT3 #(.INIT(8'hE8)) lut_n5117 (.I0(x132), .I1(x133), .I2(x134), .O(n5117));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5118 (.I0(x123), .I1(x124), .I2(x125), .I3(n5112), .I4(n5113), .O(n5118));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5119 (.I0(x129), .I1(x130), .I2(x131), .I3(n5117), .I4(n5118), .O(n5119));
  LUT3 #(.INIT(8'hE8)) lut_n5120 (.I0(x138), .I1(x139), .I2(x140), .O(n5120));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5121 (.I0(x129), .I1(x130), .I2(x131), .I3(n5117), .I4(n5118), .O(n5121));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5122 (.I0(x135), .I1(x136), .I2(x137), .I3(n5120), .I4(n5121), .O(n5122));
  LUT3 #(.INIT(8'h96)) lut_n5123 (.I0(n5111), .I1(n5114), .I2(n5115), .O(n5123));
  LUT3 #(.INIT(8'hE8)) lut_n5124 (.I0(n5119), .I1(n5122), .I2(n5123), .O(n5124));
  LUT3 #(.INIT(8'h96)) lut_n5125 (.I0(n5098), .I1(n5106), .I2(n5107), .O(n5125));
  LUT3 #(.INIT(8'hE8)) lut_n5126 (.I0(n5116), .I1(n5124), .I2(n5125), .O(n5126));
  LUT3 #(.INIT(8'h96)) lut_n5127 (.I0(n5053), .I1(n5071), .I2(n5089), .O(n5127));
  LUT3 #(.INIT(8'hE8)) lut_n5128 (.I0(n5108), .I1(n5126), .I2(n5127), .O(n5128));
  LUT3 #(.INIT(8'hE8)) lut_n5129 (.I0(x144), .I1(x145), .I2(x146), .O(n5129));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5130 (.I0(x135), .I1(x136), .I2(x137), .I3(n5120), .I4(n5121), .O(n5130));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5131 (.I0(x141), .I1(x142), .I2(x143), .I3(n5129), .I4(n5130), .O(n5131));
  LUT3 #(.INIT(8'hE8)) lut_n5132 (.I0(x150), .I1(x151), .I2(x152), .O(n5132));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5133 (.I0(x141), .I1(x142), .I2(x143), .I3(n5129), .I4(n5130), .O(n5133));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5134 (.I0(x147), .I1(x148), .I2(x149), .I3(n5132), .I4(n5133), .O(n5134));
  LUT3 #(.INIT(8'h96)) lut_n5135 (.I0(n5119), .I1(n5122), .I2(n5123), .O(n5135));
  LUT3 #(.INIT(8'hE8)) lut_n5136 (.I0(n5131), .I1(n5134), .I2(n5135), .O(n5136));
  LUT3 #(.INIT(8'hE8)) lut_n5137 (.I0(x156), .I1(x157), .I2(x158), .O(n5137));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5138 (.I0(x147), .I1(x148), .I2(x149), .I3(n5132), .I4(n5133), .O(n5138));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5139 (.I0(x153), .I1(x154), .I2(x155), .I3(n5137), .I4(n5138), .O(n5139));
  LUT3 #(.INIT(8'hE8)) lut_n5140 (.I0(x162), .I1(x163), .I2(x164), .O(n5140));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5141 (.I0(x153), .I1(x154), .I2(x155), .I3(n5137), .I4(n5138), .O(n5141));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5142 (.I0(x159), .I1(x160), .I2(x161), .I3(n5140), .I4(n5141), .O(n5142));
  LUT3 #(.INIT(8'h96)) lut_n5143 (.I0(n5131), .I1(n5134), .I2(n5135), .O(n5143));
  LUT3 #(.INIT(8'hE8)) lut_n5144 (.I0(n5139), .I1(n5142), .I2(n5143), .O(n5144));
  LUT3 #(.INIT(8'h96)) lut_n5145 (.I0(n5116), .I1(n5124), .I2(n5125), .O(n5145));
  LUT3 #(.INIT(8'hE8)) lut_n5146 (.I0(n5136), .I1(n5144), .I2(n5145), .O(n5146));
  LUT3 #(.INIT(8'hE8)) lut_n5147 (.I0(x168), .I1(x169), .I2(x170), .O(n5147));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5148 (.I0(x159), .I1(x160), .I2(x161), .I3(n5140), .I4(n5141), .O(n5148));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5149 (.I0(x165), .I1(x166), .I2(x167), .I3(n5147), .I4(n5148), .O(n5149));
  LUT3 #(.INIT(8'hE8)) lut_n5150 (.I0(x174), .I1(x175), .I2(x176), .O(n5150));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5151 (.I0(x165), .I1(x166), .I2(x167), .I3(n5147), .I4(n5148), .O(n5151));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5152 (.I0(x171), .I1(x172), .I2(x173), .I3(n5150), .I4(n5151), .O(n5152));
  LUT3 #(.INIT(8'h96)) lut_n5153 (.I0(n5139), .I1(n5142), .I2(n5143), .O(n5153));
  LUT3 #(.INIT(8'hE8)) lut_n5154 (.I0(n5149), .I1(n5152), .I2(n5153), .O(n5154));
  LUT3 #(.INIT(8'hE8)) lut_n5155 (.I0(x180), .I1(x181), .I2(x182), .O(n5155));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5156 (.I0(x171), .I1(x172), .I2(x173), .I3(n5150), .I4(n5151), .O(n5156));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5157 (.I0(x177), .I1(x178), .I2(x179), .I3(n5155), .I4(n5156), .O(n5157));
  LUT3 #(.INIT(8'hE8)) lut_n5158 (.I0(x186), .I1(x187), .I2(x188), .O(n5158));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5159 (.I0(x177), .I1(x178), .I2(x179), .I3(n5155), .I4(n5156), .O(n5159));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5160 (.I0(x183), .I1(x184), .I2(x185), .I3(n5158), .I4(n5159), .O(n5160));
  LUT3 #(.INIT(8'h96)) lut_n5161 (.I0(n5149), .I1(n5152), .I2(n5153), .O(n5161));
  LUT3 #(.INIT(8'hE8)) lut_n5162 (.I0(n5157), .I1(n5160), .I2(n5161), .O(n5162));
  LUT3 #(.INIT(8'h96)) lut_n5163 (.I0(n5136), .I1(n5144), .I2(n5145), .O(n5163));
  LUT3 #(.INIT(8'hE8)) lut_n5164 (.I0(n5154), .I1(n5162), .I2(n5163), .O(n5164));
  LUT3 #(.INIT(8'h96)) lut_n5165 (.I0(n5108), .I1(n5126), .I2(n5127), .O(n5165));
  LUT3 #(.INIT(8'hE8)) lut_n5166 (.I0(n5146), .I1(n5164), .I2(n5165), .O(n5166));
  LUT3 #(.INIT(8'hE8)) lut_n5167 (.I0(n5090), .I1(n5128), .I2(n5166), .O(n5167));
  LUT3 #(.INIT(8'hE8)) lut_n5168 (.I0(x192), .I1(x193), .I2(x194), .O(n5168));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5169 (.I0(x183), .I1(x184), .I2(x185), .I3(n5158), .I4(n5159), .O(n5169));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5170 (.I0(x189), .I1(x190), .I2(x191), .I3(n5168), .I4(n5169), .O(n5170));
  LUT3 #(.INIT(8'hE8)) lut_n5171 (.I0(x198), .I1(x199), .I2(x200), .O(n5171));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5172 (.I0(x189), .I1(x190), .I2(x191), .I3(n5168), .I4(n5169), .O(n5172));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5173 (.I0(x195), .I1(x196), .I2(x197), .I3(n5171), .I4(n5172), .O(n5173));
  LUT3 #(.INIT(8'h96)) lut_n5174 (.I0(n5157), .I1(n5160), .I2(n5161), .O(n5174));
  LUT3 #(.INIT(8'hE8)) lut_n5175 (.I0(n5170), .I1(n5173), .I2(n5174), .O(n5175));
  LUT3 #(.INIT(8'hE8)) lut_n5176 (.I0(x204), .I1(x205), .I2(x206), .O(n5176));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5177 (.I0(x195), .I1(x196), .I2(x197), .I3(n5171), .I4(n5172), .O(n5177));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5178 (.I0(x201), .I1(x202), .I2(x203), .I3(n5176), .I4(n5177), .O(n5178));
  LUT3 #(.INIT(8'hE8)) lut_n5179 (.I0(x210), .I1(x211), .I2(x212), .O(n5179));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5180 (.I0(x201), .I1(x202), .I2(x203), .I3(n5176), .I4(n5177), .O(n5180));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5181 (.I0(x207), .I1(x208), .I2(x209), .I3(n5179), .I4(n5180), .O(n5181));
  LUT3 #(.INIT(8'h96)) lut_n5182 (.I0(n5170), .I1(n5173), .I2(n5174), .O(n5182));
  LUT3 #(.INIT(8'hE8)) lut_n5183 (.I0(n5178), .I1(n5181), .I2(n5182), .O(n5183));
  LUT3 #(.INIT(8'h96)) lut_n5184 (.I0(n5154), .I1(n5162), .I2(n5163), .O(n5184));
  LUT3 #(.INIT(8'hE8)) lut_n5185 (.I0(n5175), .I1(n5183), .I2(n5184), .O(n5185));
  LUT3 #(.INIT(8'hE8)) lut_n5186 (.I0(x216), .I1(x217), .I2(x218), .O(n5186));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5187 (.I0(x207), .I1(x208), .I2(x209), .I3(n5179), .I4(n5180), .O(n5187));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5188 (.I0(x213), .I1(x214), .I2(x215), .I3(n5186), .I4(n5187), .O(n5188));
  LUT3 #(.INIT(8'hE8)) lut_n5189 (.I0(x222), .I1(x223), .I2(x224), .O(n5189));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5190 (.I0(x213), .I1(x214), .I2(x215), .I3(n5186), .I4(n5187), .O(n5190));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5191 (.I0(x219), .I1(x220), .I2(x221), .I3(n5189), .I4(n5190), .O(n5191));
  LUT3 #(.INIT(8'h96)) lut_n5192 (.I0(n5178), .I1(n5181), .I2(n5182), .O(n5192));
  LUT3 #(.INIT(8'hE8)) lut_n5193 (.I0(n5188), .I1(n5191), .I2(n5192), .O(n5193));
  LUT3 #(.INIT(8'hE8)) lut_n5194 (.I0(x228), .I1(x229), .I2(x230), .O(n5194));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5195 (.I0(x219), .I1(x220), .I2(x221), .I3(n5189), .I4(n5190), .O(n5195));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5196 (.I0(x225), .I1(x226), .I2(x227), .I3(n5194), .I4(n5195), .O(n5196));
  LUT3 #(.INIT(8'hE8)) lut_n5197 (.I0(x234), .I1(x235), .I2(x236), .O(n5197));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5198 (.I0(x225), .I1(x226), .I2(x227), .I3(n5194), .I4(n5195), .O(n5198));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5199 (.I0(x231), .I1(x232), .I2(x233), .I3(n5197), .I4(n5198), .O(n5199));
  LUT3 #(.INIT(8'h96)) lut_n5200 (.I0(n5188), .I1(n5191), .I2(n5192), .O(n5200));
  LUT3 #(.INIT(8'hE8)) lut_n5201 (.I0(n5196), .I1(n5199), .I2(n5200), .O(n5201));
  LUT3 #(.INIT(8'h96)) lut_n5202 (.I0(n5175), .I1(n5183), .I2(n5184), .O(n5202));
  LUT3 #(.INIT(8'hE8)) lut_n5203 (.I0(n5193), .I1(n5201), .I2(n5202), .O(n5203));
  LUT3 #(.INIT(8'h96)) lut_n5204 (.I0(n5146), .I1(n5164), .I2(n5165), .O(n5204));
  LUT3 #(.INIT(8'hE8)) lut_n5205 (.I0(n5185), .I1(n5203), .I2(n5204), .O(n5205));
  LUT3 #(.INIT(8'hE8)) lut_n5206 (.I0(x240), .I1(x241), .I2(x242), .O(n5206));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5207 (.I0(x231), .I1(x232), .I2(x233), .I3(n5197), .I4(n5198), .O(n5207));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5208 (.I0(x237), .I1(x238), .I2(x239), .I3(n5206), .I4(n5207), .O(n5208));
  LUT3 #(.INIT(8'hE8)) lut_n5209 (.I0(x246), .I1(x247), .I2(x248), .O(n5209));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5210 (.I0(x237), .I1(x238), .I2(x239), .I3(n5206), .I4(n5207), .O(n5210));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5211 (.I0(x243), .I1(x244), .I2(x245), .I3(n5209), .I4(n5210), .O(n5211));
  LUT3 #(.INIT(8'h96)) lut_n5212 (.I0(n5196), .I1(n5199), .I2(n5200), .O(n5212));
  LUT3 #(.INIT(8'hE8)) lut_n5213 (.I0(n5208), .I1(n5211), .I2(n5212), .O(n5213));
  LUT3 #(.INIT(8'hE8)) lut_n5214 (.I0(x252), .I1(x253), .I2(x254), .O(n5214));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5215 (.I0(x243), .I1(x244), .I2(x245), .I3(n5209), .I4(n5210), .O(n5215));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5216 (.I0(x249), .I1(x250), .I2(x251), .I3(n5214), .I4(n5215), .O(n5216));
  LUT3 #(.INIT(8'hE8)) lut_n5217 (.I0(x258), .I1(x259), .I2(x260), .O(n5217));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5218 (.I0(x249), .I1(x250), .I2(x251), .I3(n5214), .I4(n5215), .O(n5218));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5219 (.I0(x255), .I1(x256), .I2(x257), .I3(n5217), .I4(n5218), .O(n5219));
  LUT3 #(.INIT(8'h96)) lut_n5220 (.I0(n5208), .I1(n5211), .I2(n5212), .O(n5220));
  LUT3 #(.INIT(8'hE8)) lut_n5221 (.I0(n5216), .I1(n5219), .I2(n5220), .O(n5221));
  LUT3 #(.INIT(8'h96)) lut_n5222 (.I0(n5193), .I1(n5201), .I2(n5202), .O(n5222));
  LUT3 #(.INIT(8'hE8)) lut_n5223 (.I0(n5213), .I1(n5221), .I2(n5222), .O(n5223));
  LUT3 #(.INIT(8'hE8)) lut_n5224 (.I0(x264), .I1(x265), .I2(x266), .O(n5224));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5225 (.I0(x255), .I1(x256), .I2(x257), .I3(n5217), .I4(n5218), .O(n5225));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5226 (.I0(x261), .I1(x262), .I2(x263), .I3(n5224), .I4(n5225), .O(n5226));
  LUT3 #(.INIT(8'hE8)) lut_n5227 (.I0(x270), .I1(x271), .I2(x272), .O(n5227));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5228 (.I0(x261), .I1(x262), .I2(x263), .I3(n5224), .I4(n5225), .O(n5228));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5229 (.I0(x267), .I1(x268), .I2(x269), .I3(n5227), .I4(n5228), .O(n5229));
  LUT3 #(.INIT(8'h96)) lut_n5230 (.I0(n5216), .I1(n5219), .I2(n5220), .O(n5230));
  LUT3 #(.INIT(8'hE8)) lut_n5231 (.I0(n5226), .I1(n5229), .I2(n5230), .O(n5231));
  LUT3 #(.INIT(8'hE8)) lut_n5232 (.I0(x276), .I1(x277), .I2(x278), .O(n5232));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5233 (.I0(x267), .I1(x268), .I2(x269), .I3(n5227), .I4(n5228), .O(n5233));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5234 (.I0(x273), .I1(x274), .I2(x275), .I3(n5232), .I4(n5233), .O(n5234));
  LUT3 #(.INIT(8'hE8)) lut_n5235 (.I0(x282), .I1(x283), .I2(x284), .O(n5235));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5236 (.I0(x273), .I1(x274), .I2(x275), .I3(n5232), .I4(n5233), .O(n5236));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5237 (.I0(x279), .I1(x280), .I2(x281), .I3(n5235), .I4(n5236), .O(n5237));
  LUT3 #(.INIT(8'h96)) lut_n5238 (.I0(n5226), .I1(n5229), .I2(n5230), .O(n5238));
  LUT3 #(.INIT(8'hE8)) lut_n5239 (.I0(n5234), .I1(n5237), .I2(n5238), .O(n5239));
  LUT3 #(.INIT(8'h96)) lut_n5240 (.I0(n5213), .I1(n5221), .I2(n5222), .O(n5240));
  LUT3 #(.INIT(8'hE8)) lut_n5241 (.I0(n5231), .I1(n5239), .I2(n5240), .O(n5241));
  LUT3 #(.INIT(8'h96)) lut_n5242 (.I0(n5185), .I1(n5203), .I2(n5204), .O(n5242));
  LUT3 #(.INIT(8'hE8)) lut_n5243 (.I0(n5223), .I1(n5241), .I2(n5242), .O(n5243));
  LUT3 #(.INIT(8'h96)) lut_n5244 (.I0(n5090), .I1(n5128), .I2(n5166), .O(n5244));
  LUT3 #(.INIT(8'hE8)) lut_n5245 (.I0(n5205), .I1(n5243), .I2(n5244), .O(n5245));
  LUT3 #(.INIT(8'hE8)) lut_n5246 (.I0(x288), .I1(x289), .I2(x290), .O(n5246));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5247 (.I0(x279), .I1(x280), .I2(x281), .I3(n5235), .I4(n5236), .O(n5247));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5248 (.I0(x285), .I1(x286), .I2(x287), .I3(n5246), .I4(n5247), .O(n5248));
  LUT3 #(.INIT(8'hE8)) lut_n5249 (.I0(x294), .I1(x295), .I2(x296), .O(n5249));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5250 (.I0(x285), .I1(x286), .I2(x287), .I3(n5246), .I4(n5247), .O(n5250));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5251 (.I0(x291), .I1(x292), .I2(x293), .I3(n5249), .I4(n5250), .O(n5251));
  LUT3 #(.INIT(8'h96)) lut_n5252 (.I0(n5234), .I1(n5237), .I2(n5238), .O(n5252));
  LUT3 #(.INIT(8'hE8)) lut_n5253 (.I0(n5248), .I1(n5251), .I2(n5252), .O(n5253));
  LUT3 #(.INIT(8'hE8)) lut_n5254 (.I0(x297), .I1(x298), .I2(x299), .O(n5254));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5255 (.I0(x291), .I1(x292), .I2(x293), .I3(n5249), .I4(n5250), .O(n5255));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5256 (.I0(x300), .I1(x301), .I2(x302), .I3(n5254), .I4(n5255), .O(n5256));
  LUT3 #(.INIT(8'hE8)) lut_n5257 (.I0(x306), .I1(x307), .I2(x308), .O(n5257));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5258 (.I0(x300), .I1(x301), .I2(x302), .I3(n5254), .I4(n5255), .O(n5258));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5259 (.I0(x303), .I1(x304), .I2(x305), .I3(n5257), .I4(n5258), .O(n5259));
  LUT3 #(.INIT(8'h96)) lut_n5260 (.I0(n5248), .I1(n5251), .I2(n5252), .O(n5260));
  LUT3 #(.INIT(8'hE8)) lut_n5261 (.I0(n5256), .I1(n5259), .I2(n5260), .O(n5261));
  LUT3 #(.INIT(8'h96)) lut_n5262 (.I0(n5231), .I1(n5239), .I2(n5240), .O(n5262));
  LUT3 #(.INIT(8'hE8)) lut_n5263 (.I0(n5253), .I1(n5261), .I2(n5262), .O(n5263));
  LUT3 #(.INIT(8'hE8)) lut_n5264 (.I0(x312), .I1(x313), .I2(x314), .O(n5264));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5265 (.I0(x303), .I1(x304), .I2(x305), .I3(n5257), .I4(n5258), .O(n5265));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5266 (.I0(x309), .I1(x310), .I2(x311), .I3(n5264), .I4(n5265), .O(n5266));
  LUT3 #(.INIT(8'hE8)) lut_n5267 (.I0(x318), .I1(x319), .I2(x320), .O(n5267));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5268 (.I0(x309), .I1(x310), .I2(x311), .I3(n5264), .I4(n5265), .O(n5268));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5269 (.I0(x315), .I1(x316), .I2(x317), .I3(n5267), .I4(n5268), .O(n5269));
  LUT3 #(.INIT(8'h96)) lut_n5270 (.I0(n5256), .I1(n5259), .I2(n5260), .O(n5270));
  LUT3 #(.INIT(8'hE8)) lut_n5271 (.I0(n5266), .I1(n5269), .I2(n5270), .O(n5271));
  LUT3 #(.INIT(8'hE8)) lut_n5272 (.I0(x324), .I1(x325), .I2(x326), .O(n5272));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5273 (.I0(x315), .I1(x316), .I2(x317), .I3(n5267), .I4(n5268), .O(n5273));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5274 (.I0(x321), .I1(x322), .I2(x323), .I3(n5272), .I4(n5273), .O(n5274));
  LUT3 #(.INIT(8'hE8)) lut_n5275 (.I0(x330), .I1(x331), .I2(x332), .O(n5275));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5276 (.I0(x321), .I1(x322), .I2(x323), .I3(n5272), .I4(n5273), .O(n5276));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5277 (.I0(x327), .I1(x328), .I2(x329), .I3(n5275), .I4(n5276), .O(n5277));
  LUT3 #(.INIT(8'h96)) lut_n5278 (.I0(n5266), .I1(n5269), .I2(n5270), .O(n5278));
  LUT3 #(.INIT(8'hE8)) lut_n5279 (.I0(n5274), .I1(n5277), .I2(n5278), .O(n5279));
  LUT3 #(.INIT(8'h96)) lut_n5280 (.I0(n5253), .I1(n5261), .I2(n5262), .O(n5280));
  LUT3 #(.INIT(8'hE8)) lut_n5281 (.I0(n5271), .I1(n5279), .I2(n5280), .O(n5281));
  LUT3 #(.INIT(8'h96)) lut_n5282 (.I0(n5223), .I1(n5241), .I2(n5242), .O(n5282));
  LUT3 #(.INIT(8'hE8)) lut_n5283 (.I0(n5263), .I1(n5281), .I2(n5282), .O(n5283));
  LUT3 #(.INIT(8'hE8)) lut_n5284 (.I0(x336), .I1(x337), .I2(x338), .O(n5284));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5285 (.I0(x327), .I1(x328), .I2(x329), .I3(n5275), .I4(n5276), .O(n5285));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5286 (.I0(x333), .I1(x334), .I2(x335), .I3(n5284), .I4(n5285), .O(n5286));
  LUT3 #(.INIT(8'hE8)) lut_n5287 (.I0(x342), .I1(x343), .I2(x344), .O(n5287));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5288 (.I0(x333), .I1(x334), .I2(x335), .I3(n5284), .I4(n5285), .O(n5288));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5289 (.I0(x339), .I1(x340), .I2(x341), .I3(n5287), .I4(n5288), .O(n5289));
  LUT3 #(.INIT(8'h96)) lut_n5290 (.I0(n5274), .I1(n5277), .I2(n5278), .O(n5290));
  LUT3 #(.INIT(8'hE8)) lut_n5291 (.I0(n5286), .I1(n5289), .I2(n5290), .O(n5291));
  LUT3 #(.INIT(8'hE8)) lut_n5292 (.I0(x348), .I1(x349), .I2(x350), .O(n5292));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5293 (.I0(x339), .I1(x340), .I2(x341), .I3(n5287), .I4(n5288), .O(n5293));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5294 (.I0(x345), .I1(x346), .I2(x347), .I3(n5292), .I4(n5293), .O(n5294));
  LUT3 #(.INIT(8'hE8)) lut_n5295 (.I0(x354), .I1(x355), .I2(x356), .O(n5295));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5296 (.I0(x345), .I1(x346), .I2(x347), .I3(n5292), .I4(n5293), .O(n5296));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5297 (.I0(x351), .I1(x352), .I2(x353), .I3(n5295), .I4(n5296), .O(n5297));
  LUT3 #(.INIT(8'h96)) lut_n5298 (.I0(n5286), .I1(n5289), .I2(n5290), .O(n5298));
  LUT3 #(.INIT(8'hE8)) lut_n5299 (.I0(n5294), .I1(n5297), .I2(n5298), .O(n5299));
  LUT3 #(.INIT(8'h96)) lut_n5300 (.I0(n5271), .I1(n5279), .I2(n5280), .O(n5300));
  LUT3 #(.INIT(8'hE8)) lut_n5301 (.I0(n5291), .I1(n5299), .I2(n5300), .O(n5301));
  LUT3 #(.INIT(8'hE8)) lut_n5302 (.I0(x360), .I1(x361), .I2(x362), .O(n5302));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5303 (.I0(x351), .I1(x352), .I2(x353), .I3(n5295), .I4(n5296), .O(n5303));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5304 (.I0(x357), .I1(x358), .I2(x359), .I3(n5302), .I4(n5303), .O(n5304));
  LUT3 #(.INIT(8'hE8)) lut_n5305 (.I0(x366), .I1(x367), .I2(x368), .O(n5305));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5306 (.I0(x357), .I1(x358), .I2(x359), .I3(n5302), .I4(n5303), .O(n5306));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5307 (.I0(x363), .I1(x364), .I2(x365), .I3(n5305), .I4(n5306), .O(n5307));
  LUT3 #(.INIT(8'h96)) lut_n5308 (.I0(n5294), .I1(n5297), .I2(n5298), .O(n5308));
  LUT3 #(.INIT(8'hE8)) lut_n5309 (.I0(n5304), .I1(n5307), .I2(n5308), .O(n5309));
  LUT3 #(.INIT(8'hE8)) lut_n5310 (.I0(x372), .I1(x373), .I2(x374), .O(n5310));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5311 (.I0(x363), .I1(x364), .I2(x365), .I3(n5305), .I4(n5306), .O(n5311));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5312 (.I0(x369), .I1(x370), .I2(x371), .I3(n5310), .I4(n5311), .O(n5312));
  LUT3 #(.INIT(8'hE8)) lut_n5313 (.I0(x378), .I1(x379), .I2(x380), .O(n5313));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5314 (.I0(x369), .I1(x370), .I2(x371), .I3(n5310), .I4(n5311), .O(n5314));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5315 (.I0(x375), .I1(x376), .I2(x377), .I3(n5313), .I4(n5314), .O(n5315));
  LUT3 #(.INIT(8'h96)) lut_n5316 (.I0(n5304), .I1(n5307), .I2(n5308), .O(n5316));
  LUT3 #(.INIT(8'hE8)) lut_n5317 (.I0(n5312), .I1(n5315), .I2(n5316), .O(n5317));
  LUT3 #(.INIT(8'h96)) lut_n5318 (.I0(n5291), .I1(n5299), .I2(n5300), .O(n5318));
  LUT3 #(.INIT(8'hE8)) lut_n5319 (.I0(n5309), .I1(n5317), .I2(n5318), .O(n5319));
  LUT3 #(.INIT(8'h96)) lut_n5320 (.I0(n5263), .I1(n5281), .I2(n5282), .O(n5320));
  LUT3 #(.INIT(8'hE8)) lut_n5321 (.I0(n5301), .I1(n5319), .I2(n5320), .O(n5321));
  LUT3 #(.INIT(8'h96)) lut_n5322 (.I0(n5205), .I1(n5243), .I2(n5244), .O(n5322));
  LUT3 #(.INIT(8'hE8)) lut_n5323 (.I0(n5283), .I1(n5321), .I2(n5322), .O(n5323));
  LUT3 #(.INIT(8'hE8)) lut_n5324 (.I0(n5167), .I1(n5245), .I2(n5323), .O(n5324));
  LUT3 #(.INIT(8'hE8)) lut_n5325 (.I0(x384), .I1(x385), .I2(x386), .O(n5325));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5326 (.I0(x375), .I1(x376), .I2(x377), .I3(n5313), .I4(n5314), .O(n5326));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5327 (.I0(x381), .I1(x382), .I2(x383), .I3(n5325), .I4(n5326), .O(n5327));
  LUT3 #(.INIT(8'hE8)) lut_n5328 (.I0(x390), .I1(x391), .I2(x392), .O(n5328));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5329 (.I0(x381), .I1(x382), .I2(x383), .I3(n5325), .I4(n5326), .O(n5329));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5330 (.I0(x387), .I1(x388), .I2(x389), .I3(n5328), .I4(n5329), .O(n5330));
  LUT3 #(.INIT(8'h96)) lut_n5331 (.I0(n5312), .I1(n5315), .I2(n5316), .O(n5331));
  LUT3 #(.INIT(8'hE8)) lut_n5332 (.I0(n5327), .I1(n5330), .I2(n5331), .O(n5332));
  LUT3 #(.INIT(8'hE8)) lut_n5333 (.I0(x396), .I1(x397), .I2(x398), .O(n5333));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5334 (.I0(x387), .I1(x388), .I2(x389), .I3(n5328), .I4(n5329), .O(n5334));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5335 (.I0(x393), .I1(x394), .I2(x395), .I3(n5333), .I4(n5334), .O(n5335));
  LUT3 #(.INIT(8'hE8)) lut_n5336 (.I0(x402), .I1(x403), .I2(x404), .O(n5336));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5337 (.I0(x393), .I1(x394), .I2(x395), .I3(n5333), .I4(n5334), .O(n5337));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5338 (.I0(x399), .I1(x400), .I2(x401), .I3(n5336), .I4(n5337), .O(n5338));
  LUT3 #(.INIT(8'h96)) lut_n5339 (.I0(n5327), .I1(n5330), .I2(n5331), .O(n5339));
  LUT3 #(.INIT(8'hE8)) lut_n5340 (.I0(n5335), .I1(n5338), .I2(n5339), .O(n5340));
  LUT3 #(.INIT(8'h96)) lut_n5341 (.I0(n5309), .I1(n5317), .I2(n5318), .O(n5341));
  LUT3 #(.INIT(8'hE8)) lut_n5342 (.I0(n5332), .I1(n5340), .I2(n5341), .O(n5342));
  LUT3 #(.INIT(8'hE8)) lut_n5343 (.I0(x408), .I1(x409), .I2(x410), .O(n5343));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5344 (.I0(x399), .I1(x400), .I2(x401), .I3(n5336), .I4(n5337), .O(n5344));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5345 (.I0(x405), .I1(x406), .I2(x407), .I3(n5343), .I4(n5344), .O(n5345));
  LUT3 #(.INIT(8'hE8)) lut_n5346 (.I0(x414), .I1(x415), .I2(x416), .O(n5346));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5347 (.I0(x405), .I1(x406), .I2(x407), .I3(n5343), .I4(n5344), .O(n5347));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5348 (.I0(x411), .I1(x412), .I2(x413), .I3(n5346), .I4(n5347), .O(n5348));
  LUT3 #(.INIT(8'h96)) lut_n5349 (.I0(n5335), .I1(n5338), .I2(n5339), .O(n5349));
  LUT3 #(.INIT(8'hE8)) lut_n5350 (.I0(n5345), .I1(n5348), .I2(n5349), .O(n5350));
  LUT3 #(.INIT(8'hE8)) lut_n5351 (.I0(x420), .I1(x421), .I2(x422), .O(n5351));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5352 (.I0(x411), .I1(x412), .I2(x413), .I3(n5346), .I4(n5347), .O(n5352));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5353 (.I0(x417), .I1(x418), .I2(x419), .I3(n5351), .I4(n5352), .O(n5353));
  LUT3 #(.INIT(8'hE8)) lut_n5354 (.I0(x426), .I1(x427), .I2(x428), .O(n5354));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5355 (.I0(x417), .I1(x418), .I2(x419), .I3(n5351), .I4(n5352), .O(n5355));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5356 (.I0(x423), .I1(x424), .I2(x425), .I3(n5354), .I4(n5355), .O(n5356));
  LUT3 #(.INIT(8'h96)) lut_n5357 (.I0(n5345), .I1(n5348), .I2(n5349), .O(n5357));
  LUT3 #(.INIT(8'hE8)) lut_n5358 (.I0(n5353), .I1(n5356), .I2(n5357), .O(n5358));
  LUT3 #(.INIT(8'h96)) lut_n5359 (.I0(n5332), .I1(n5340), .I2(n5341), .O(n5359));
  LUT3 #(.INIT(8'hE8)) lut_n5360 (.I0(n5350), .I1(n5358), .I2(n5359), .O(n5360));
  LUT3 #(.INIT(8'h96)) lut_n5361 (.I0(n5301), .I1(n5319), .I2(n5320), .O(n5361));
  LUT3 #(.INIT(8'hE8)) lut_n5362 (.I0(n5342), .I1(n5360), .I2(n5361), .O(n5362));
  LUT3 #(.INIT(8'hE8)) lut_n5363 (.I0(x432), .I1(x433), .I2(x434), .O(n5363));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5364 (.I0(x423), .I1(x424), .I2(x425), .I3(n5354), .I4(n5355), .O(n5364));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5365 (.I0(x429), .I1(x430), .I2(x431), .I3(n5363), .I4(n5364), .O(n5365));
  LUT3 #(.INIT(8'hE8)) lut_n5366 (.I0(x438), .I1(x439), .I2(x440), .O(n5366));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5367 (.I0(x429), .I1(x430), .I2(x431), .I3(n5363), .I4(n5364), .O(n5367));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5368 (.I0(x435), .I1(x436), .I2(x437), .I3(n5366), .I4(n5367), .O(n5368));
  LUT3 #(.INIT(8'h96)) lut_n5369 (.I0(n5353), .I1(n5356), .I2(n5357), .O(n5369));
  LUT3 #(.INIT(8'hE8)) lut_n5370 (.I0(n5365), .I1(n5368), .I2(n5369), .O(n5370));
  LUT3 #(.INIT(8'hE8)) lut_n5371 (.I0(x444), .I1(x445), .I2(x446), .O(n5371));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5372 (.I0(x435), .I1(x436), .I2(x437), .I3(n5366), .I4(n5367), .O(n5372));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5373 (.I0(x441), .I1(x442), .I2(x443), .I3(n5371), .I4(n5372), .O(n5373));
  LUT3 #(.INIT(8'hE8)) lut_n5374 (.I0(x450), .I1(x451), .I2(x452), .O(n5374));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5375 (.I0(x441), .I1(x442), .I2(x443), .I3(n5371), .I4(n5372), .O(n5375));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5376 (.I0(x447), .I1(x448), .I2(x449), .I3(n5374), .I4(n5375), .O(n5376));
  LUT3 #(.INIT(8'h96)) lut_n5377 (.I0(n5365), .I1(n5368), .I2(n5369), .O(n5377));
  LUT3 #(.INIT(8'hE8)) lut_n5378 (.I0(n5373), .I1(n5376), .I2(n5377), .O(n5378));
  LUT3 #(.INIT(8'h96)) lut_n5379 (.I0(n5350), .I1(n5358), .I2(n5359), .O(n5379));
  LUT3 #(.INIT(8'hE8)) lut_n5380 (.I0(n5370), .I1(n5378), .I2(n5379), .O(n5380));
  LUT3 #(.INIT(8'hE8)) lut_n5381 (.I0(x456), .I1(x457), .I2(x458), .O(n5381));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5382 (.I0(x447), .I1(x448), .I2(x449), .I3(n5374), .I4(n5375), .O(n5382));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5383 (.I0(x453), .I1(x454), .I2(x455), .I3(n5381), .I4(n5382), .O(n5383));
  LUT3 #(.INIT(8'hE8)) lut_n5384 (.I0(x462), .I1(x463), .I2(x464), .O(n5384));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5385 (.I0(x453), .I1(x454), .I2(x455), .I3(n5381), .I4(n5382), .O(n5385));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5386 (.I0(x459), .I1(x460), .I2(x461), .I3(n5384), .I4(n5385), .O(n5386));
  LUT3 #(.INIT(8'h96)) lut_n5387 (.I0(n5373), .I1(n5376), .I2(n5377), .O(n5387));
  LUT3 #(.INIT(8'hE8)) lut_n5388 (.I0(n5383), .I1(n5386), .I2(n5387), .O(n5388));
  LUT3 #(.INIT(8'hE8)) lut_n5389 (.I0(x468), .I1(x469), .I2(x470), .O(n5389));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5390 (.I0(x459), .I1(x460), .I2(x461), .I3(n5384), .I4(n5385), .O(n5390));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5391 (.I0(x465), .I1(x466), .I2(x467), .I3(n5389), .I4(n5390), .O(n5391));
  LUT3 #(.INIT(8'hE8)) lut_n5392 (.I0(x474), .I1(x475), .I2(x476), .O(n5392));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5393 (.I0(x465), .I1(x466), .I2(x467), .I3(n5389), .I4(n5390), .O(n5393));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5394 (.I0(x471), .I1(x472), .I2(x473), .I3(n5392), .I4(n5393), .O(n5394));
  LUT3 #(.INIT(8'h96)) lut_n5395 (.I0(n5383), .I1(n5386), .I2(n5387), .O(n5395));
  LUT3 #(.INIT(8'hE8)) lut_n5396 (.I0(n5391), .I1(n5394), .I2(n5395), .O(n5396));
  LUT3 #(.INIT(8'h96)) lut_n5397 (.I0(n5370), .I1(n5378), .I2(n5379), .O(n5397));
  LUT3 #(.INIT(8'hE8)) lut_n5398 (.I0(n5388), .I1(n5396), .I2(n5397), .O(n5398));
  LUT3 #(.INIT(8'h96)) lut_n5399 (.I0(n5342), .I1(n5360), .I2(n5361), .O(n5399));
  LUT3 #(.INIT(8'hE8)) lut_n5400 (.I0(n5380), .I1(n5398), .I2(n5399), .O(n5400));
  LUT3 #(.INIT(8'h96)) lut_n5401 (.I0(n5283), .I1(n5321), .I2(n5322), .O(n5401));
  LUT3 #(.INIT(8'hE8)) lut_n5402 (.I0(n5362), .I1(n5400), .I2(n5401), .O(n5402));
  LUT3 #(.INIT(8'hE8)) lut_n5403 (.I0(x480), .I1(x481), .I2(x482), .O(n5403));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5404 (.I0(x471), .I1(x472), .I2(x473), .I3(n5392), .I4(n5393), .O(n5404));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5405 (.I0(x477), .I1(x478), .I2(x479), .I3(n5403), .I4(n5404), .O(n5405));
  LUT3 #(.INIT(8'hE8)) lut_n5406 (.I0(x486), .I1(x487), .I2(x488), .O(n5406));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5407 (.I0(x477), .I1(x478), .I2(x479), .I3(n5403), .I4(n5404), .O(n5407));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5408 (.I0(x483), .I1(x484), .I2(x485), .I3(n5406), .I4(n5407), .O(n5408));
  LUT3 #(.INIT(8'h96)) lut_n5409 (.I0(n5391), .I1(n5394), .I2(n5395), .O(n5409));
  LUT3 #(.INIT(8'hE8)) lut_n5410 (.I0(n5405), .I1(n5408), .I2(n5409), .O(n5410));
  LUT3 #(.INIT(8'hE8)) lut_n5411 (.I0(x492), .I1(x493), .I2(x494), .O(n5411));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5412 (.I0(x483), .I1(x484), .I2(x485), .I3(n5406), .I4(n5407), .O(n5412));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5413 (.I0(x489), .I1(x490), .I2(x491), .I3(n5411), .I4(n5412), .O(n5413));
  LUT3 #(.INIT(8'hE8)) lut_n5414 (.I0(x498), .I1(x499), .I2(x500), .O(n5414));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5415 (.I0(x489), .I1(x490), .I2(x491), .I3(n5411), .I4(n5412), .O(n5415));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5416 (.I0(x495), .I1(x496), .I2(x497), .I3(n5414), .I4(n5415), .O(n5416));
  LUT3 #(.INIT(8'h96)) lut_n5417 (.I0(n5405), .I1(n5408), .I2(n5409), .O(n5417));
  LUT3 #(.INIT(8'hE8)) lut_n5418 (.I0(n5413), .I1(n5416), .I2(n5417), .O(n5418));
  LUT3 #(.INIT(8'h96)) lut_n5419 (.I0(n5388), .I1(n5396), .I2(n5397), .O(n5419));
  LUT3 #(.INIT(8'hE8)) lut_n5420 (.I0(n5410), .I1(n5418), .I2(n5419), .O(n5420));
  LUT3 #(.INIT(8'hE8)) lut_n5421 (.I0(x504), .I1(x505), .I2(x506), .O(n5421));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5422 (.I0(x495), .I1(x496), .I2(x497), .I3(n5414), .I4(n5415), .O(n5422));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5423 (.I0(x501), .I1(x502), .I2(x503), .I3(n5421), .I4(n5422), .O(n5423));
  LUT3 #(.INIT(8'hE8)) lut_n5424 (.I0(x510), .I1(x511), .I2(x512), .O(n5424));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5425 (.I0(x501), .I1(x502), .I2(x503), .I3(n5421), .I4(n5422), .O(n5425));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5426 (.I0(x507), .I1(x508), .I2(x509), .I3(n5424), .I4(n5425), .O(n5426));
  LUT3 #(.INIT(8'h96)) lut_n5427 (.I0(n5413), .I1(n5416), .I2(n5417), .O(n5427));
  LUT3 #(.INIT(8'hE8)) lut_n5428 (.I0(n5423), .I1(n5426), .I2(n5427), .O(n5428));
  LUT3 #(.INIT(8'hE8)) lut_n5429 (.I0(x516), .I1(x517), .I2(x518), .O(n5429));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5430 (.I0(x507), .I1(x508), .I2(x509), .I3(n5424), .I4(n5425), .O(n5430));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5431 (.I0(x513), .I1(x514), .I2(x515), .I3(n5429), .I4(n5430), .O(n5431));
  LUT3 #(.INIT(8'hE8)) lut_n5432 (.I0(x522), .I1(x523), .I2(x524), .O(n5432));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5433 (.I0(x513), .I1(x514), .I2(x515), .I3(n5429), .I4(n5430), .O(n5433));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5434 (.I0(x519), .I1(x520), .I2(x521), .I3(n5432), .I4(n5433), .O(n5434));
  LUT3 #(.INIT(8'h96)) lut_n5435 (.I0(n5423), .I1(n5426), .I2(n5427), .O(n5435));
  LUT3 #(.INIT(8'hE8)) lut_n5436 (.I0(n5431), .I1(n5434), .I2(n5435), .O(n5436));
  LUT3 #(.INIT(8'h96)) lut_n5437 (.I0(n5410), .I1(n5418), .I2(n5419), .O(n5437));
  LUT3 #(.INIT(8'hE8)) lut_n5438 (.I0(n5428), .I1(n5436), .I2(n5437), .O(n5438));
  LUT3 #(.INIT(8'h96)) lut_n5439 (.I0(n5380), .I1(n5398), .I2(n5399), .O(n5439));
  LUT3 #(.INIT(8'hE8)) lut_n5440 (.I0(n5420), .I1(n5438), .I2(n5439), .O(n5440));
  LUT3 #(.INIT(8'hE8)) lut_n5441 (.I0(x528), .I1(x529), .I2(x530), .O(n5441));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5442 (.I0(x519), .I1(x520), .I2(x521), .I3(n5432), .I4(n5433), .O(n5442));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5443 (.I0(x525), .I1(x526), .I2(x527), .I3(n5441), .I4(n5442), .O(n5443));
  LUT3 #(.INIT(8'hE8)) lut_n5444 (.I0(x534), .I1(x535), .I2(x536), .O(n5444));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5445 (.I0(x525), .I1(x526), .I2(x527), .I3(n5441), .I4(n5442), .O(n5445));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5446 (.I0(x531), .I1(x532), .I2(x533), .I3(n5444), .I4(n5445), .O(n5446));
  LUT3 #(.INIT(8'h96)) lut_n5447 (.I0(n5431), .I1(n5434), .I2(n5435), .O(n5447));
  LUT3 #(.INIT(8'hE8)) lut_n5448 (.I0(n5443), .I1(n5446), .I2(n5447), .O(n5448));
  LUT3 #(.INIT(8'hE8)) lut_n5449 (.I0(x540), .I1(x541), .I2(x542), .O(n5449));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5450 (.I0(x531), .I1(x532), .I2(x533), .I3(n5444), .I4(n5445), .O(n5450));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5451 (.I0(x537), .I1(x538), .I2(x539), .I3(n5449), .I4(n5450), .O(n5451));
  LUT3 #(.INIT(8'hE8)) lut_n5452 (.I0(x546), .I1(x547), .I2(x548), .O(n5452));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5453 (.I0(x537), .I1(x538), .I2(x539), .I3(n5449), .I4(n5450), .O(n5453));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5454 (.I0(x543), .I1(x544), .I2(x545), .I3(n5452), .I4(n5453), .O(n5454));
  LUT3 #(.INIT(8'h96)) lut_n5455 (.I0(n5443), .I1(n5446), .I2(n5447), .O(n5455));
  LUT3 #(.INIT(8'hE8)) lut_n5456 (.I0(n5451), .I1(n5454), .I2(n5455), .O(n5456));
  LUT3 #(.INIT(8'h96)) lut_n5457 (.I0(n5428), .I1(n5436), .I2(n5437), .O(n5457));
  LUT3 #(.INIT(8'hE8)) lut_n5458 (.I0(n5448), .I1(n5456), .I2(n5457), .O(n5458));
  LUT3 #(.INIT(8'hE8)) lut_n5459 (.I0(x552), .I1(x553), .I2(x554), .O(n5459));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5460 (.I0(x543), .I1(x544), .I2(x545), .I3(n5452), .I4(n5453), .O(n5460));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5461 (.I0(x549), .I1(x550), .I2(x551), .I3(n5459), .I4(n5460), .O(n5461));
  LUT3 #(.INIT(8'hE8)) lut_n5462 (.I0(x558), .I1(x559), .I2(x560), .O(n5462));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5463 (.I0(x549), .I1(x550), .I2(x551), .I3(n5459), .I4(n5460), .O(n5463));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5464 (.I0(x555), .I1(x556), .I2(x557), .I3(n5462), .I4(n5463), .O(n5464));
  LUT3 #(.INIT(8'h96)) lut_n5465 (.I0(n5451), .I1(n5454), .I2(n5455), .O(n5465));
  LUT3 #(.INIT(8'hE8)) lut_n5466 (.I0(n5461), .I1(n5464), .I2(n5465), .O(n5466));
  LUT3 #(.INIT(8'hE8)) lut_n5467 (.I0(x564), .I1(x565), .I2(x566), .O(n5467));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5468 (.I0(x555), .I1(x556), .I2(x557), .I3(n5462), .I4(n5463), .O(n5468));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5469 (.I0(x561), .I1(x562), .I2(x563), .I3(n5467), .I4(n5468), .O(n5469));
  LUT3 #(.INIT(8'hE8)) lut_n5470 (.I0(x570), .I1(x571), .I2(x572), .O(n5470));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5471 (.I0(x561), .I1(x562), .I2(x563), .I3(n5467), .I4(n5468), .O(n5471));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5472 (.I0(x567), .I1(x568), .I2(x569), .I3(n5470), .I4(n5471), .O(n5472));
  LUT3 #(.INIT(8'h96)) lut_n5473 (.I0(n5461), .I1(n5464), .I2(n5465), .O(n5473));
  LUT3 #(.INIT(8'hE8)) lut_n5474 (.I0(n5469), .I1(n5472), .I2(n5473), .O(n5474));
  LUT3 #(.INIT(8'h96)) lut_n5475 (.I0(n5448), .I1(n5456), .I2(n5457), .O(n5475));
  LUT3 #(.INIT(8'hE8)) lut_n5476 (.I0(n5466), .I1(n5474), .I2(n5475), .O(n5476));
  LUT3 #(.INIT(8'h96)) lut_n5477 (.I0(n5420), .I1(n5438), .I2(n5439), .O(n5477));
  LUT3 #(.INIT(8'hE8)) lut_n5478 (.I0(n5458), .I1(n5476), .I2(n5477), .O(n5478));
  LUT3 #(.INIT(8'h96)) lut_n5479 (.I0(n5362), .I1(n5400), .I2(n5401), .O(n5479));
  LUT3 #(.INIT(8'hE8)) lut_n5480 (.I0(n5440), .I1(n5478), .I2(n5479), .O(n5480));
  LUT3 #(.INIT(8'h96)) lut_n5481 (.I0(n5167), .I1(n5245), .I2(n5323), .O(n5481));
  LUT3 #(.INIT(8'hE8)) lut_n5482 (.I0(n5402), .I1(n5480), .I2(n5481), .O(n5482));
  LUT3 #(.INIT(8'hE8)) lut_n5483 (.I0(x576), .I1(x577), .I2(x578), .O(n5483));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5484 (.I0(x567), .I1(x568), .I2(x569), .I3(n5470), .I4(n5471), .O(n5484));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5485 (.I0(x573), .I1(x574), .I2(x575), .I3(n5483), .I4(n5484), .O(n5485));
  LUT3 #(.INIT(8'hE8)) lut_n5486 (.I0(x582), .I1(x583), .I2(x584), .O(n5486));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5487 (.I0(x573), .I1(x574), .I2(x575), .I3(n5483), .I4(n5484), .O(n5487));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5488 (.I0(x579), .I1(x580), .I2(x581), .I3(n5486), .I4(n5487), .O(n5488));
  LUT3 #(.INIT(8'h96)) lut_n5489 (.I0(n5469), .I1(n5472), .I2(n5473), .O(n5489));
  LUT3 #(.INIT(8'hE8)) lut_n5490 (.I0(n5485), .I1(n5488), .I2(n5489), .O(n5490));
  LUT3 #(.INIT(8'hE8)) lut_n5491 (.I0(x588), .I1(x589), .I2(x590), .O(n5491));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5492 (.I0(x579), .I1(x580), .I2(x581), .I3(n5486), .I4(n5487), .O(n5492));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5493 (.I0(x585), .I1(x586), .I2(x587), .I3(n5491), .I4(n5492), .O(n5493));
  LUT3 #(.INIT(8'hE8)) lut_n5494 (.I0(x594), .I1(x595), .I2(x596), .O(n5494));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5495 (.I0(x585), .I1(x586), .I2(x587), .I3(n5491), .I4(n5492), .O(n5495));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5496 (.I0(x591), .I1(x592), .I2(x593), .I3(n5494), .I4(n5495), .O(n5496));
  LUT3 #(.INIT(8'h96)) lut_n5497 (.I0(n5485), .I1(n5488), .I2(n5489), .O(n5497));
  LUT3 #(.INIT(8'hE8)) lut_n5498 (.I0(n5493), .I1(n5496), .I2(n5497), .O(n5498));
  LUT3 #(.INIT(8'h96)) lut_n5499 (.I0(n5466), .I1(n5474), .I2(n5475), .O(n5499));
  LUT3 #(.INIT(8'hE8)) lut_n5500 (.I0(n5490), .I1(n5498), .I2(n5499), .O(n5500));
  LUT3 #(.INIT(8'hE8)) lut_n5501 (.I0(x600), .I1(x601), .I2(x602), .O(n5501));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5502 (.I0(x591), .I1(x592), .I2(x593), .I3(n5494), .I4(n5495), .O(n5502));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5503 (.I0(x597), .I1(x598), .I2(x599), .I3(n5501), .I4(n5502), .O(n5503));
  LUT3 #(.INIT(8'hE8)) lut_n5504 (.I0(x606), .I1(x607), .I2(x608), .O(n5504));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5505 (.I0(x597), .I1(x598), .I2(x599), .I3(n5501), .I4(n5502), .O(n5505));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5506 (.I0(x603), .I1(x604), .I2(x605), .I3(n5504), .I4(n5505), .O(n5506));
  LUT3 #(.INIT(8'h96)) lut_n5507 (.I0(n5493), .I1(n5496), .I2(n5497), .O(n5507));
  LUT3 #(.INIT(8'hE8)) lut_n5508 (.I0(n5503), .I1(n5506), .I2(n5507), .O(n5508));
  LUT3 #(.INIT(8'hE8)) lut_n5509 (.I0(x612), .I1(x613), .I2(x614), .O(n5509));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5510 (.I0(x603), .I1(x604), .I2(x605), .I3(n5504), .I4(n5505), .O(n5510));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5511 (.I0(x609), .I1(x610), .I2(x611), .I3(n5509), .I4(n5510), .O(n5511));
  LUT3 #(.INIT(8'hE8)) lut_n5512 (.I0(x618), .I1(x619), .I2(x620), .O(n5512));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5513 (.I0(x609), .I1(x610), .I2(x611), .I3(n5509), .I4(n5510), .O(n5513));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5514 (.I0(x615), .I1(x616), .I2(x617), .I3(n5512), .I4(n5513), .O(n5514));
  LUT3 #(.INIT(8'h96)) lut_n5515 (.I0(n5503), .I1(n5506), .I2(n5507), .O(n5515));
  LUT3 #(.INIT(8'hE8)) lut_n5516 (.I0(n5511), .I1(n5514), .I2(n5515), .O(n5516));
  LUT3 #(.INIT(8'h96)) lut_n5517 (.I0(n5490), .I1(n5498), .I2(n5499), .O(n5517));
  LUT3 #(.INIT(8'hE8)) lut_n5518 (.I0(n5508), .I1(n5516), .I2(n5517), .O(n5518));
  LUT3 #(.INIT(8'h96)) lut_n5519 (.I0(n5458), .I1(n5476), .I2(n5477), .O(n5519));
  LUT3 #(.INIT(8'hE8)) lut_n5520 (.I0(n5500), .I1(n5518), .I2(n5519), .O(n5520));
  LUT3 #(.INIT(8'hE8)) lut_n5521 (.I0(x624), .I1(x625), .I2(x626), .O(n5521));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5522 (.I0(x615), .I1(x616), .I2(x617), .I3(n5512), .I4(n5513), .O(n5522));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5523 (.I0(x621), .I1(x622), .I2(x623), .I3(n5521), .I4(n5522), .O(n5523));
  LUT3 #(.INIT(8'hE8)) lut_n5524 (.I0(x630), .I1(x631), .I2(x632), .O(n5524));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5525 (.I0(x621), .I1(x622), .I2(x623), .I3(n5521), .I4(n5522), .O(n5525));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5526 (.I0(x627), .I1(x628), .I2(x629), .I3(n5524), .I4(n5525), .O(n5526));
  LUT3 #(.INIT(8'h96)) lut_n5527 (.I0(n5511), .I1(n5514), .I2(n5515), .O(n5527));
  LUT3 #(.INIT(8'hE8)) lut_n5528 (.I0(n5523), .I1(n5526), .I2(n5527), .O(n5528));
  LUT3 #(.INIT(8'hE8)) lut_n5529 (.I0(x636), .I1(x637), .I2(x638), .O(n5529));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5530 (.I0(x627), .I1(x628), .I2(x629), .I3(n5524), .I4(n5525), .O(n5530));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5531 (.I0(x633), .I1(x634), .I2(x635), .I3(n5529), .I4(n5530), .O(n5531));
  LUT3 #(.INIT(8'hE8)) lut_n5532 (.I0(x642), .I1(x643), .I2(x644), .O(n5532));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5533 (.I0(x633), .I1(x634), .I2(x635), .I3(n5529), .I4(n5530), .O(n5533));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5534 (.I0(x639), .I1(x640), .I2(x641), .I3(n5532), .I4(n5533), .O(n5534));
  LUT3 #(.INIT(8'h96)) lut_n5535 (.I0(n5523), .I1(n5526), .I2(n5527), .O(n5535));
  LUT3 #(.INIT(8'hE8)) lut_n5536 (.I0(n5531), .I1(n5534), .I2(n5535), .O(n5536));
  LUT3 #(.INIT(8'h96)) lut_n5537 (.I0(n5508), .I1(n5516), .I2(n5517), .O(n5537));
  LUT3 #(.INIT(8'hE8)) lut_n5538 (.I0(n5528), .I1(n5536), .I2(n5537), .O(n5538));
  LUT3 #(.INIT(8'hE8)) lut_n5539 (.I0(x648), .I1(x649), .I2(x650), .O(n5539));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5540 (.I0(x639), .I1(x640), .I2(x641), .I3(n5532), .I4(n5533), .O(n5540));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5541 (.I0(x645), .I1(x646), .I2(x647), .I3(n5539), .I4(n5540), .O(n5541));
  LUT3 #(.INIT(8'hE8)) lut_n5542 (.I0(x654), .I1(x655), .I2(x656), .O(n5542));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5543 (.I0(x645), .I1(x646), .I2(x647), .I3(n5539), .I4(n5540), .O(n5543));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5544 (.I0(x651), .I1(x652), .I2(x653), .I3(n5542), .I4(n5543), .O(n5544));
  LUT3 #(.INIT(8'h96)) lut_n5545 (.I0(n5531), .I1(n5534), .I2(n5535), .O(n5545));
  LUT3 #(.INIT(8'hE8)) lut_n5546 (.I0(n5541), .I1(n5544), .I2(n5545), .O(n5546));
  LUT3 #(.INIT(8'hE8)) lut_n5547 (.I0(x660), .I1(x661), .I2(x662), .O(n5547));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5548 (.I0(x651), .I1(x652), .I2(x653), .I3(n5542), .I4(n5543), .O(n5548));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5549 (.I0(x657), .I1(x658), .I2(x659), .I3(n5547), .I4(n5548), .O(n5549));
  LUT3 #(.INIT(8'hE8)) lut_n5550 (.I0(x666), .I1(x667), .I2(x668), .O(n5550));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5551 (.I0(x657), .I1(x658), .I2(x659), .I3(n5547), .I4(n5548), .O(n5551));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5552 (.I0(x663), .I1(x664), .I2(x665), .I3(n5550), .I4(n5551), .O(n5552));
  LUT3 #(.INIT(8'h96)) lut_n5553 (.I0(n5541), .I1(n5544), .I2(n5545), .O(n5553));
  LUT3 #(.INIT(8'hE8)) lut_n5554 (.I0(n5549), .I1(n5552), .I2(n5553), .O(n5554));
  LUT3 #(.INIT(8'h96)) lut_n5555 (.I0(n5528), .I1(n5536), .I2(n5537), .O(n5555));
  LUT3 #(.INIT(8'hE8)) lut_n5556 (.I0(n5546), .I1(n5554), .I2(n5555), .O(n5556));
  LUT3 #(.INIT(8'h96)) lut_n5557 (.I0(n5500), .I1(n5518), .I2(n5519), .O(n5557));
  LUT3 #(.INIT(8'hE8)) lut_n5558 (.I0(n5538), .I1(n5556), .I2(n5557), .O(n5558));
  LUT3 #(.INIT(8'h96)) lut_n5559 (.I0(n5440), .I1(n5478), .I2(n5479), .O(n5559));
  LUT3 #(.INIT(8'hE8)) lut_n5560 (.I0(n5520), .I1(n5558), .I2(n5559), .O(n5560));
  LUT3 #(.INIT(8'hE8)) lut_n5561 (.I0(x672), .I1(x673), .I2(x674), .O(n5561));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5562 (.I0(x663), .I1(x664), .I2(x665), .I3(n5550), .I4(n5551), .O(n5562));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5563 (.I0(x669), .I1(x670), .I2(x671), .I3(n5561), .I4(n5562), .O(n5563));
  LUT3 #(.INIT(8'hE8)) lut_n5564 (.I0(x678), .I1(x679), .I2(x680), .O(n5564));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5565 (.I0(x669), .I1(x670), .I2(x671), .I3(n5561), .I4(n5562), .O(n5565));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5566 (.I0(x675), .I1(x676), .I2(x677), .I3(n5564), .I4(n5565), .O(n5566));
  LUT3 #(.INIT(8'h96)) lut_n5567 (.I0(n5549), .I1(n5552), .I2(n5553), .O(n5567));
  LUT3 #(.INIT(8'hE8)) lut_n5568 (.I0(n5563), .I1(n5566), .I2(n5567), .O(n5568));
  LUT3 #(.INIT(8'hE8)) lut_n5569 (.I0(x684), .I1(x685), .I2(x686), .O(n5569));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5570 (.I0(x675), .I1(x676), .I2(x677), .I3(n5564), .I4(n5565), .O(n5570));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5571 (.I0(x681), .I1(x682), .I2(x683), .I3(n5569), .I4(n5570), .O(n5571));
  LUT3 #(.INIT(8'hE8)) lut_n5572 (.I0(x690), .I1(x691), .I2(x692), .O(n5572));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5573 (.I0(x681), .I1(x682), .I2(x683), .I3(n5569), .I4(n5570), .O(n5573));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5574 (.I0(x687), .I1(x688), .I2(x689), .I3(n5572), .I4(n5573), .O(n5574));
  LUT3 #(.INIT(8'h96)) lut_n5575 (.I0(n5563), .I1(n5566), .I2(n5567), .O(n5575));
  LUT3 #(.INIT(8'hE8)) lut_n5576 (.I0(n5571), .I1(n5574), .I2(n5575), .O(n5576));
  LUT3 #(.INIT(8'h96)) lut_n5577 (.I0(n5546), .I1(n5554), .I2(n5555), .O(n5577));
  LUT3 #(.INIT(8'hE8)) lut_n5578 (.I0(n5568), .I1(n5576), .I2(n5577), .O(n5578));
  LUT3 #(.INIT(8'hE8)) lut_n5579 (.I0(x696), .I1(x697), .I2(x698), .O(n5579));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5580 (.I0(x687), .I1(x688), .I2(x689), .I3(n5572), .I4(n5573), .O(n5580));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5581 (.I0(x693), .I1(x694), .I2(x695), .I3(n5579), .I4(n5580), .O(n5581));
  LUT3 #(.INIT(8'hE8)) lut_n5582 (.I0(x702), .I1(x703), .I2(x704), .O(n5582));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5583 (.I0(x693), .I1(x694), .I2(x695), .I3(n5579), .I4(n5580), .O(n5583));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5584 (.I0(x699), .I1(x700), .I2(x701), .I3(n5582), .I4(n5583), .O(n5584));
  LUT3 #(.INIT(8'h96)) lut_n5585 (.I0(n5571), .I1(n5574), .I2(n5575), .O(n5585));
  LUT3 #(.INIT(8'hE8)) lut_n5586 (.I0(n5581), .I1(n5584), .I2(n5585), .O(n5586));
  LUT3 #(.INIT(8'hE8)) lut_n5587 (.I0(x708), .I1(x709), .I2(x710), .O(n5587));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5588 (.I0(x699), .I1(x700), .I2(x701), .I3(n5582), .I4(n5583), .O(n5588));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5589 (.I0(x705), .I1(x706), .I2(x707), .I3(n5587), .I4(n5588), .O(n5589));
  LUT3 #(.INIT(8'hE8)) lut_n5590 (.I0(x714), .I1(x715), .I2(x716), .O(n5590));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5591 (.I0(x705), .I1(x706), .I2(x707), .I3(n5587), .I4(n5588), .O(n5591));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5592 (.I0(x711), .I1(x712), .I2(x713), .I3(n5590), .I4(n5591), .O(n5592));
  LUT3 #(.INIT(8'h96)) lut_n5593 (.I0(n5581), .I1(n5584), .I2(n5585), .O(n5593));
  LUT3 #(.INIT(8'hE8)) lut_n5594 (.I0(n5589), .I1(n5592), .I2(n5593), .O(n5594));
  LUT3 #(.INIT(8'h96)) lut_n5595 (.I0(n5568), .I1(n5576), .I2(n5577), .O(n5595));
  LUT3 #(.INIT(8'hE8)) lut_n5596 (.I0(n5586), .I1(n5594), .I2(n5595), .O(n5596));
  LUT3 #(.INIT(8'h96)) lut_n5597 (.I0(n5538), .I1(n5556), .I2(n5557), .O(n5597));
  LUT3 #(.INIT(8'hE8)) lut_n5598 (.I0(n5578), .I1(n5596), .I2(n5597), .O(n5598));
  LUT3 #(.INIT(8'hE8)) lut_n5599 (.I0(x720), .I1(x721), .I2(x722), .O(n5599));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5600 (.I0(x711), .I1(x712), .I2(x713), .I3(n5590), .I4(n5591), .O(n5600));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5601 (.I0(x717), .I1(x718), .I2(x719), .I3(n5599), .I4(n5600), .O(n5601));
  LUT3 #(.INIT(8'hE8)) lut_n5602 (.I0(x726), .I1(x727), .I2(x728), .O(n5602));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5603 (.I0(x717), .I1(x718), .I2(x719), .I3(n5599), .I4(n5600), .O(n5603));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5604 (.I0(x723), .I1(x724), .I2(x725), .I3(n5602), .I4(n5603), .O(n5604));
  LUT3 #(.INIT(8'h96)) lut_n5605 (.I0(n5589), .I1(n5592), .I2(n5593), .O(n5605));
  LUT3 #(.INIT(8'hE8)) lut_n5606 (.I0(n5601), .I1(n5604), .I2(n5605), .O(n5606));
  LUT3 #(.INIT(8'hE8)) lut_n5607 (.I0(x732), .I1(x733), .I2(x734), .O(n5607));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5608 (.I0(x723), .I1(x724), .I2(x725), .I3(n5602), .I4(n5603), .O(n5608));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5609 (.I0(x729), .I1(x730), .I2(x731), .I3(n5607), .I4(n5608), .O(n5609));
  LUT3 #(.INIT(8'hE8)) lut_n5610 (.I0(x738), .I1(x739), .I2(x740), .O(n5610));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5611 (.I0(x729), .I1(x730), .I2(x731), .I3(n5607), .I4(n5608), .O(n5611));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5612 (.I0(x735), .I1(x736), .I2(x737), .I3(n5610), .I4(n5611), .O(n5612));
  LUT3 #(.INIT(8'h96)) lut_n5613 (.I0(n5601), .I1(n5604), .I2(n5605), .O(n5613));
  LUT3 #(.INIT(8'hE8)) lut_n5614 (.I0(n5609), .I1(n5612), .I2(n5613), .O(n5614));
  LUT3 #(.INIT(8'h96)) lut_n5615 (.I0(n5586), .I1(n5594), .I2(n5595), .O(n5615));
  LUT3 #(.INIT(8'hE8)) lut_n5616 (.I0(n5606), .I1(n5614), .I2(n5615), .O(n5616));
  LUT3 #(.INIT(8'hE8)) lut_n5617 (.I0(x744), .I1(x745), .I2(x746), .O(n5617));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5618 (.I0(x735), .I1(x736), .I2(x737), .I3(n5610), .I4(n5611), .O(n5618));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5619 (.I0(x741), .I1(x742), .I2(x743), .I3(n5617), .I4(n5618), .O(n5619));
  LUT3 #(.INIT(8'hE8)) lut_n5620 (.I0(x750), .I1(x751), .I2(x752), .O(n5620));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5621 (.I0(x741), .I1(x742), .I2(x743), .I3(n5617), .I4(n5618), .O(n5621));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5622 (.I0(x747), .I1(x748), .I2(x749), .I3(n5620), .I4(n5621), .O(n5622));
  LUT3 #(.INIT(8'h96)) lut_n5623 (.I0(n5609), .I1(n5612), .I2(n5613), .O(n5623));
  LUT3 #(.INIT(8'hE8)) lut_n5624 (.I0(n5619), .I1(n5622), .I2(n5623), .O(n5624));
  LUT3 #(.INIT(8'hE8)) lut_n5625 (.I0(x756), .I1(x757), .I2(x758), .O(n5625));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5626 (.I0(x747), .I1(x748), .I2(x749), .I3(n5620), .I4(n5621), .O(n5626));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5627 (.I0(x753), .I1(x754), .I2(x755), .I3(n5625), .I4(n5626), .O(n5627));
  LUT3 #(.INIT(8'hE8)) lut_n5628 (.I0(x762), .I1(x763), .I2(x764), .O(n5628));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5629 (.I0(x753), .I1(x754), .I2(x755), .I3(n5625), .I4(n5626), .O(n5629));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5630 (.I0(x759), .I1(x760), .I2(x761), .I3(n5628), .I4(n5629), .O(n5630));
  LUT3 #(.INIT(8'h96)) lut_n5631 (.I0(n5619), .I1(n5622), .I2(n5623), .O(n5631));
  LUT3 #(.INIT(8'hE8)) lut_n5632 (.I0(n5627), .I1(n5630), .I2(n5631), .O(n5632));
  LUT3 #(.INIT(8'h96)) lut_n5633 (.I0(n5606), .I1(n5614), .I2(n5615), .O(n5633));
  LUT3 #(.INIT(8'hE8)) lut_n5634 (.I0(n5624), .I1(n5632), .I2(n5633), .O(n5634));
  LUT3 #(.INIT(8'h96)) lut_n5635 (.I0(n5578), .I1(n5596), .I2(n5597), .O(n5635));
  LUT3 #(.INIT(8'hE8)) lut_n5636 (.I0(n5616), .I1(n5634), .I2(n5635), .O(n5636));
  LUT3 #(.INIT(8'h96)) lut_n5637 (.I0(n5520), .I1(n5558), .I2(n5559), .O(n5637));
  LUT3 #(.INIT(8'hE8)) lut_n5638 (.I0(n5598), .I1(n5636), .I2(n5637), .O(n5638));
  LUT3 #(.INIT(8'h96)) lut_n5639 (.I0(n5402), .I1(n5480), .I2(n5481), .O(n5639));
  LUT3 #(.INIT(8'hE8)) lut_n5640 (.I0(n5560), .I1(n5638), .I2(n5639), .O(n5640));
  LUT3 #(.INIT(8'hE8)) lut_n5641 (.I0(n5324), .I1(n5482), .I2(n5640), .O(n5641));
  LUT3 #(.INIT(8'hE8)) lut_n5642 (.I0(x768), .I1(x769), .I2(x770), .O(n5642));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5643 (.I0(x759), .I1(x760), .I2(x761), .I3(n5628), .I4(n5629), .O(n5643));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5644 (.I0(x765), .I1(x766), .I2(x767), .I3(n5642), .I4(n5643), .O(n5644));
  LUT3 #(.INIT(8'hE8)) lut_n5645 (.I0(x774), .I1(x775), .I2(x776), .O(n5645));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5646 (.I0(x765), .I1(x766), .I2(x767), .I3(n5642), .I4(n5643), .O(n5646));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5647 (.I0(x771), .I1(x772), .I2(x773), .I3(n5645), .I4(n5646), .O(n5647));
  LUT3 #(.INIT(8'h96)) lut_n5648 (.I0(n5627), .I1(n5630), .I2(n5631), .O(n5648));
  LUT3 #(.INIT(8'hE8)) lut_n5649 (.I0(n5644), .I1(n5647), .I2(n5648), .O(n5649));
  LUT3 #(.INIT(8'hE8)) lut_n5650 (.I0(x780), .I1(x781), .I2(x782), .O(n5650));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5651 (.I0(x771), .I1(x772), .I2(x773), .I3(n5645), .I4(n5646), .O(n5651));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5652 (.I0(x777), .I1(x778), .I2(x779), .I3(n5650), .I4(n5651), .O(n5652));
  LUT3 #(.INIT(8'hE8)) lut_n5653 (.I0(x786), .I1(x787), .I2(x788), .O(n5653));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5654 (.I0(x777), .I1(x778), .I2(x779), .I3(n5650), .I4(n5651), .O(n5654));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5655 (.I0(x783), .I1(x784), .I2(x785), .I3(n5653), .I4(n5654), .O(n5655));
  LUT3 #(.INIT(8'h96)) lut_n5656 (.I0(n5644), .I1(n5647), .I2(n5648), .O(n5656));
  LUT3 #(.INIT(8'hE8)) lut_n5657 (.I0(n5652), .I1(n5655), .I2(n5656), .O(n5657));
  LUT3 #(.INIT(8'h96)) lut_n5658 (.I0(n5624), .I1(n5632), .I2(n5633), .O(n5658));
  LUT3 #(.INIT(8'hE8)) lut_n5659 (.I0(n5649), .I1(n5657), .I2(n5658), .O(n5659));
  LUT3 #(.INIT(8'hE8)) lut_n5660 (.I0(x792), .I1(x793), .I2(x794), .O(n5660));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5661 (.I0(x783), .I1(x784), .I2(x785), .I3(n5653), .I4(n5654), .O(n5661));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5662 (.I0(x789), .I1(x790), .I2(x791), .I3(n5660), .I4(n5661), .O(n5662));
  LUT3 #(.INIT(8'hE8)) lut_n5663 (.I0(x798), .I1(x799), .I2(x800), .O(n5663));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5664 (.I0(x789), .I1(x790), .I2(x791), .I3(n5660), .I4(n5661), .O(n5664));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5665 (.I0(x795), .I1(x796), .I2(x797), .I3(n5663), .I4(n5664), .O(n5665));
  LUT3 #(.INIT(8'h96)) lut_n5666 (.I0(n5652), .I1(n5655), .I2(n5656), .O(n5666));
  LUT3 #(.INIT(8'hE8)) lut_n5667 (.I0(n5662), .I1(n5665), .I2(n5666), .O(n5667));
  LUT3 #(.INIT(8'hE8)) lut_n5668 (.I0(x804), .I1(x805), .I2(x806), .O(n5668));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5669 (.I0(x795), .I1(x796), .I2(x797), .I3(n5663), .I4(n5664), .O(n5669));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5670 (.I0(x801), .I1(x802), .I2(x803), .I3(n5668), .I4(n5669), .O(n5670));
  LUT3 #(.INIT(8'hE8)) lut_n5671 (.I0(x810), .I1(x811), .I2(x812), .O(n5671));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5672 (.I0(x801), .I1(x802), .I2(x803), .I3(n5668), .I4(n5669), .O(n5672));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5673 (.I0(x807), .I1(x808), .I2(x809), .I3(n5671), .I4(n5672), .O(n5673));
  LUT3 #(.INIT(8'h96)) lut_n5674 (.I0(n5662), .I1(n5665), .I2(n5666), .O(n5674));
  LUT3 #(.INIT(8'hE8)) lut_n5675 (.I0(n5670), .I1(n5673), .I2(n5674), .O(n5675));
  LUT3 #(.INIT(8'h96)) lut_n5676 (.I0(n5649), .I1(n5657), .I2(n5658), .O(n5676));
  LUT3 #(.INIT(8'hE8)) lut_n5677 (.I0(n5667), .I1(n5675), .I2(n5676), .O(n5677));
  LUT3 #(.INIT(8'h96)) lut_n5678 (.I0(n5616), .I1(n5634), .I2(n5635), .O(n5678));
  LUT3 #(.INIT(8'hE8)) lut_n5679 (.I0(n5659), .I1(n5677), .I2(n5678), .O(n5679));
  LUT3 #(.INIT(8'hE8)) lut_n5680 (.I0(x816), .I1(x817), .I2(x818), .O(n5680));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5681 (.I0(x807), .I1(x808), .I2(x809), .I3(n5671), .I4(n5672), .O(n5681));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5682 (.I0(x813), .I1(x814), .I2(x815), .I3(n5680), .I4(n5681), .O(n5682));
  LUT3 #(.INIT(8'hE8)) lut_n5683 (.I0(x822), .I1(x823), .I2(x824), .O(n5683));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5684 (.I0(x813), .I1(x814), .I2(x815), .I3(n5680), .I4(n5681), .O(n5684));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5685 (.I0(x819), .I1(x820), .I2(x821), .I3(n5683), .I4(n5684), .O(n5685));
  LUT3 #(.INIT(8'h96)) lut_n5686 (.I0(n5670), .I1(n5673), .I2(n5674), .O(n5686));
  LUT3 #(.INIT(8'hE8)) lut_n5687 (.I0(n5682), .I1(n5685), .I2(n5686), .O(n5687));
  LUT3 #(.INIT(8'hE8)) lut_n5688 (.I0(x828), .I1(x829), .I2(x830), .O(n5688));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5689 (.I0(x819), .I1(x820), .I2(x821), .I3(n5683), .I4(n5684), .O(n5689));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5690 (.I0(x825), .I1(x826), .I2(x827), .I3(n5688), .I4(n5689), .O(n5690));
  LUT3 #(.INIT(8'hE8)) lut_n5691 (.I0(x834), .I1(x835), .I2(x836), .O(n5691));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5692 (.I0(x825), .I1(x826), .I2(x827), .I3(n5688), .I4(n5689), .O(n5692));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5693 (.I0(x831), .I1(x832), .I2(x833), .I3(n5691), .I4(n5692), .O(n5693));
  LUT3 #(.INIT(8'h96)) lut_n5694 (.I0(n5682), .I1(n5685), .I2(n5686), .O(n5694));
  LUT3 #(.INIT(8'hE8)) lut_n5695 (.I0(n5690), .I1(n5693), .I2(n5694), .O(n5695));
  LUT3 #(.INIT(8'h96)) lut_n5696 (.I0(n5667), .I1(n5675), .I2(n5676), .O(n5696));
  LUT3 #(.INIT(8'hE8)) lut_n5697 (.I0(n5687), .I1(n5695), .I2(n5696), .O(n5697));
  LUT3 #(.INIT(8'hE8)) lut_n5698 (.I0(x840), .I1(x841), .I2(x842), .O(n5698));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5699 (.I0(x831), .I1(x832), .I2(x833), .I3(n5691), .I4(n5692), .O(n5699));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5700 (.I0(x837), .I1(x838), .I2(x839), .I3(n5698), .I4(n5699), .O(n5700));
  LUT3 #(.INIT(8'hE8)) lut_n5701 (.I0(x846), .I1(x847), .I2(x848), .O(n5701));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5702 (.I0(x837), .I1(x838), .I2(x839), .I3(n5698), .I4(n5699), .O(n5702));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5703 (.I0(x843), .I1(x844), .I2(x845), .I3(n5701), .I4(n5702), .O(n5703));
  LUT3 #(.INIT(8'h96)) lut_n5704 (.I0(n5690), .I1(n5693), .I2(n5694), .O(n5704));
  LUT3 #(.INIT(8'hE8)) lut_n5705 (.I0(n5700), .I1(n5703), .I2(n5704), .O(n5705));
  LUT3 #(.INIT(8'hE8)) lut_n5706 (.I0(x852), .I1(x853), .I2(x854), .O(n5706));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5707 (.I0(x843), .I1(x844), .I2(x845), .I3(n5701), .I4(n5702), .O(n5707));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5708 (.I0(x849), .I1(x850), .I2(x851), .I3(n5706), .I4(n5707), .O(n5708));
  LUT3 #(.INIT(8'hE8)) lut_n5709 (.I0(x858), .I1(x859), .I2(x860), .O(n5709));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5710 (.I0(x849), .I1(x850), .I2(x851), .I3(n5706), .I4(n5707), .O(n5710));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5711 (.I0(x855), .I1(x856), .I2(x857), .I3(n5709), .I4(n5710), .O(n5711));
  LUT3 #(.INIT(8'h96)) lut_n5712 (.I0(n5700), .I1(n5703), .I2(n5704), .O(n5712));
  LUT3 #(.INIT(8'hE8)) lut_n5713 (.I0(n5708), .I1(n5711), .I2(n5712), .O(n5713));
  LUT3 #(.INIT(8'h96)) lut_n5714 (.I0(n5687), .I1(n5695), .I2(n5696), .O(n5714));
  LUT3 #(.INIT(8'hE8)) lut_n5715 (.I0(n5705), .I1(n5713), .I2(n5714), .O(n5715));
  LUT3 #(.INIT(8'h96)) lut_n5716 (.I0(n5659), .I1(n5677), .I2(n5678), .O(n5716));
  LUT3 #(.INIT(8'hE8)) lut_n5717 (.I0(n5697), .I1(n5715), .I2(n5716), .O(n5717));
  LUT3 #(.INIT(8'h96)) lut_n5718 (.I0(n5598), .I1(n5636), .I2(n5637), .O(n5718));
  LUT3 #(.INIT(8'hE8)) lut_n5719 (.I0(n5679), .I1(n5717), .I2(n5718), .O(n5719));
  LUT3 #(.INIT(8'hE8)) lut_n5720 (.I0(x864), .I1(x865), .I2(x866), .O(n5720));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5721 (.I0(x855), .I1(x856), .I2(x857), .I3(n5709), .I4(n5710), .O(n5721));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5722 (.I0(x861), .I1(x862), .I2(x863), .I3(n5720), .I4(n5721), .O(n5722));
  LUT3 #(.INIT(8'hE8)) lut_n5723 (.I0(x870), .I1(x871), .I2(x872), .O(n5723));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5724 (.I0(x861), .I1(x862), .I2(x863), .I3(n5720), .I4(n5721), .O(n5724));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5725 (.I0(x867), .I1(x868), .I2(x869), .I3(n5723), .I4(n5724), .O(n5725));
  LUT3 #(.INIT(8'h96)) lut_n5726 (.I0(n5708), .I1(n5711), .I2(n5712), .O(n5726));
  LUT3 #(.INIT(8'hE8)) lut_n5727 (.I0(n5722), .I1(n5725), .I2(n5726), .O(n5727));
  LUT3 #(.INIT(8'hE8)) lut_n5728 (.I0(x876), .I1(x877), .I2(x878), .O(n5728));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5729 (.I0(x867), .I1(x868), .I2(x869), .I3(n5723), .I4(n5724), .O(n5729));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5730 (.I0(x873), .I1(x874), .I2(x875), .I3(n5728), .I4(n5729), .O(n5730));
  LUT3 #(.INIT(8'hE8)) lut_n5731 (.I0(x882), .I1(x883), .I2(x884), .O(n5731));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5732 (.I0(x873), .I1(x874), .I2(x875), .I3(n5728), .I4(n5729), .O(n5732));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5733 (.I0(x879), .I1(x880), .I2(x881), .I3(n5731), .I4(n5732), .O(n5733));
  LUT3 #(.INIT(8'h96)) lut_n5734 (.I0(n5722), .I1(n5725), .I2(n5726), .O(n5734));
  LUT3 #(.INIT(8'hE8)) lut_n5735 (.I0(n5730), .I1(n5733), .I2(n5734), .O(n5735));
  LUT3 #(.INIT(8'h96)) lut_n5736 (.I0(n5705), .I1(n5713), .I2(n5714), .O(n5736));
  LUT3 #(.INIT(8'hE8)) lut_n5737 (.I0(n5727), .I1(n5735), .I2(n5736), .O(n5737));
  LUT3 #(.INIT(8'hE8)) lut_n5738 (.I0(x888), .I1(x889), .I2(x890), .O(n5738));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5739 (.I0(x879), .I1(x880), .I2(x881), .I3(n5731), .I4(n5732), .O(n5739));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5740 (.I0(x885), .I1(x886), .I2(x887), .I3(n5738), .I4(n5739), .O(n5740));
  LUT3 #(.INIT(8'hE8)) lut_n5741 (.I0(x894), .I1(x895), .I2(x896), .O(n5741));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5742 (.I0(x885), .I1(x886), .I2(x887), .I3(n5738), .I4(n5739), .O(n5742));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5743 (.I0(x891), .I1(x892), .I2(x893), .I3(n5741), .I4(n5742), .O(n5743));
  LUT3 #(.INIT(8'h96)) lut_n5744 (.I0(n5730), .I1(n5733), .I2(n5734), .O(n5744));
  LUT3 #(.INIT(8'hE8)) lut_n5745 (.I0(n5740), .I1(n5743), .I2(n5744), .O(n5745));
  LUT3 #(.INIT(8'hE8)) lut_n5746 (.I0(x900), .I1(x901), .I2(x902), .O(n5746));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5747 (.I0(x891), .I1(x892), .I2(x893), .I3(n5741), .I4(n5742), .O(n5747));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5748 (.I0(x897), .I1(x898), .I2(x899), .I3(n5746), .I4(n5747), .O(n5748));
  LUT3 #(.INIT(8'hE8)) lut_n5749 (.I0(x906), .I1(x907), .I2(x908), .O(n5749));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5750 (.I0(x897), .I1(x898), .I2(x899), .I3(n5746), .I4(n5747), .O(n5750));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5751 (.I0(x903), .I1(x904), .I2(x905), .I3(n5749), .I4(n5750), .O(n5751));
  LUT3 #(.INIT(8'h96)) lut_n5752 (.I0(n5740), .I1(n5743), .I2(n5744), .O(n5752));
  LUT3 #(.INIT(8'hE8)) lut_n5753 (.I0(n5748), .I1(n5751), .I2(n5752), .O(n5753));
  LUT3 #(.INIT(8'h96)) lut_n5754 (.I0(n5727), .I1(n5735), .I2(n5736), .O(n5754));
  LUT3 #(.INIT(8'hE8)) lut_n5755 (.I0(n5745), .I1(n5753), .I2(n5754), .O(n5755));
  LUT3 #(.INIT(8'h96)) lut_n5756 (.I0(n5697), .I1(n5715), .I2(n5716), .O(n5756));
  LUT3 #(.INIT(8'hE8)) lut_n5757 (.I0(n5737), .I1(n5755), .I2(n5756), .O(n5757));
  LUT3 #(.INIT(8'hE8)) lut_n5758 (.I0(x912), .I1(x913), .I2(x914), .O(n5758));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5759 (.I0(x903), .I1(x904), .I2(x905), .I3(n5749), .I4(n5750), .O(n5759));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5760 (.I0(x909), .I1(x910), .I2(x911), .I3(n5758), .I4(n5759), .O(n5760));
  LUT3 #(.INIT(8'hE8)) lut_n5761 (.I0(x918), .I1(x919), .I2(x920), .O(n5761));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5762 (.I0(x909), .I1(x910), .I2(x911), .I3(n5758), .I4(n5759), .O(n5762));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5763 (.I0(x915), .I1(x916), .I2(x917), .I3(n5761), .I4(n5762), .O(n5763));
  LUT3 #(.INIT(8'h96)) lut_n5764 (.I0(n5748), .I1(n5751), .I2(n5752), .O(n5764));
  LUT3 #(.INIT(8'hE8)) lut_n5765 (.I0(n5760), .I1(n5763), .I2(n5764), .O(n5765));
  LUT3 #(.INIT(8'hE8)) lut_n5766 (.I0(x924), .I1(x925), .I2(x926), .O(n5766));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5767 (.I0(x915), .I1(x916), .I2(x917), .I3(n5761), .I4(n5762), .O(n5767));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5768 (.I0(x921), .I1(x922), .I2(x923), .I3(n5766), .I4(n5767), .O(n5768));
  LUT3 #(.INIT(8'hE8)) lut_n5769 (.I0(x930), .I1(x931), .I2(x932), .O(n5769));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5770 (.I0(x921), .I1(x922), .I2(x923), .I3(n5766), .I4(n5767), .O(n5770));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5771 (.I0(x927), .I1(x928), .I2(x929), .I3(n5769), .I4(n5770), .O(n5771));
  LUT3 #(.INIT(8'h96)) lut_n5772 (.I0(n5760), .I1(n5763), .I2(n5764), .O(n5772));
  LUT3 #(.INIT(8'hE8)) lut_n5773 (.I0(n5768), .I1(n5771), .I2(n5772), .O(n5773));
  LUT3 #(.INIT(8'h96)) lut_n5774 (.I0(n5745), .I1(n5753), .I2(n5754), .O(n5774));
  LUT3 #(.INIT(8'hE8)) lut_n5775 (.I0(n5765), .I1(n5773), .I2(n5774), .O(n5775));
  LUT3 #(.INIT(8'hE8)) lut_n5776 (.I0(x936), .I1(x937), .I2(x938), .O(n5776));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5777 (.I0(x927), .I1(x928), .I2(x929), .I3(n5769), .I4(n5770), .O(n5777));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5778 (.I0(x933), .I1(x934), .I2(x935), .I3(n5776), .I4(n5777), .O(n5778));
  LUT3 #(.INIT(8'hE8)) lut_n5779 (.I0(x942), .I1(x943), .I2(x944), .O(n5779));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5780 (.I0(x933), .I1(x934), .I2(x935), .I3(n5776), .I4(n5777), .O(n5780));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5781 (.I0(x939), .I1(x940), .I2(x941), .I3(n5779), .I4(n5780), .O(n5781));
  LUT3 #(.INIT(8'h96)) lut_n5782 (.I0(n5768), .I1(n5771), .I2(n5772), .O(n5782));
  LUT3 #(.INIT(8'hE8)) lut_n5783 (.I0(n5778), .I1(n5781), .I2(n5782), .O(n5783));
  LUT3 #(.INIT(8'hE8)) lut_n5784 (.I0(x948), .I1(x949), .I2(x950), .O(n5784));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5785 (.I0(x939), .I1(x940), .I2(x941), .I3(n5779), .I4(n5780), .O(n5785));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5786 (.I0(x945), .I1(x946), .I2(x947), .I3(n5784), .I4(n5785), .O(n5786));
  LUT3 #(.INIT(8'hE8)) lut_n5787 (.I0(x954), .I1(x955), .I2(x956), .O(n5787));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5788 (.I0(x945), .I1(x946), .I2(x947), .I3(n5784), .I4(n5785), .O(n5788));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5789 (.I0(x951), .I1(x952), .I2(x953), .I3(n5787), .I4(n5788), .O(n5789));
  LUT3 #(.INIT(8'h96)) lut_n5790 (.I0(n5778), .I1(n5781), .I2(n5782), .O(n5790));
  LUT3 #(.INIT(8'hE8)) lut_n5791 (.I0(n5786), .I1(n5789), .I2(n5790), .O(n5791));
  LUT3 #(.INIT(8'h96)) lut_n5792 (.I0(n5765), .I1(n5773), .I2(n5774), .O(n5792));
  LUT3 #(.INIT(8'hE8)) lut_n5793 (.I0(n5783), .I1(n5791), .I2(n5792), .O(n5793));
  LUT3 #(.INIT(8'h96)) lut_n5794 (.I0(n5737), .I1(n5755), .I2(n5756), .O(n5794));
  LUT3 #(.INIT(8'hE8)) lut_n5795 (.I0(n5775), .I1(n5793), .I2(n5794), .O(n5795));
  LUT3 #(.INIT(8'h96)) lut_n5796 (.I0(n5679), .I1(n5717), .I2(n5718), .O(n5796));
  LUT3 #(.INIT(8'hE8)) lut_n5797 (.I0(n5757), .I1(n5795), .I2(n5796), .O(n5797));
  LUT3 #(.INIT(8'h96)) lut_n5798 (.I0(n5560), .I1(n5638), .I2(n5639), .O(n5798));
  LUT3 #(.INIT(8'hE8)) lut_n5799 (.I0(n5719), .I1(n5797), .I2(n5798), .O(n5799));
  LUT3 #(.INIT(8'hE8)) lut_n5800 (.I0(x960), .I1(x961), .I2(x962), .O(n5800));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5801 (.I0(x951), .I1(x952), .I2(x953), .I3(n5787), .I4(n5788), .O(n5801));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5802 (.I0(x957), .I1(x958), .I2(x959), .I3(n5800), .I4(n5801), .O(n5802));
  LUT3 #(.INIT(8'hE8)) lut_n5803 (.I0(x966), .I1(x967), .I2(x968), .O(n5803));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5804 (.I0(x957), .I1(x958), .I2(x959), .I3(n5800), .I4(n5801), .O(n5804));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5805 (.I0(x963), .I1(x964), .I2(x965), .I3(n5803), .I4(n5804), .O(n5805));
  LUT3 #(.INIT(8'h96)) lut_n5806 (.I0(n5786), .I1(n5789), .I2(n5790), .O(n5806));
  LUT3 #(.INIT(8'hE8)) lut_n5807 (.I0(n5802), .I1(n5805), .I2(n5806), .O(n5807));
  LUT3 #(.INIT(8'hE8)) lut_n5808 (.I0(x972), .I1(x973), .I2(x974), .O(n5808));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5809 (.I0(x963), .I1(x964), .I2(x965), .I3(n5803), .I4(n5804), .O(n5809));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5810 (.I0(x969), .I1(x970), .I2(x971), .I3(n5808), .I4(n5809), .O(n5810));
  LUT3 #(.INIT(8'hE8)) lut_n5811 (.I0(x978), .I1(x979), .I2(x980), .O(n5811));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5812 (.I0(x969), .I1(x970), .I2(x971), .I3(n5808), .I4(n5809), .O(n5812));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5813 (.I0(x975), .I1(x976), .I2(x977), .I3(n5811), .I4(n5812), .O(n5813));
  LUT3 #(.INIT(8'h96)) lut_n5814 (.I0(n5802), .I1(n5805), .I2(n5806), .O(n5814));
  LUT3 #(.INIT(8'hE8)) lut_n5815 (.I0(n5810), .I1(n5813), .I2(n5814), .O(n5815));
  LUT3 #(.INIT(8'h96)) lut_n5816 (.I0(n5783), .I1(n5791), .I2(n5792), .O(n5816));
  LUT3 #(.INIT(8'hE8)) lut_n5817 (.I0(n5807), .I1(n5815), .I2(n5816), .O(n5817));
  LUT3 #(.INIT(8'hE8)) lut_n5818 (.I0(x984), .I1(x985), .I2(x986), .O(n5818));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5819 (.I0(x975), .I1(x976), .I2(x977), .I3(n5811), .I4(n5812), .O(n5819));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5820 (.I0(x981), .I1(x982), .I2(x983), .I3(n5818), .I4(n5819), .O(n5820));
  LUT3 #(.INIT(8'hE8)) lut_n5821 (.I0(x990), .I1(x991), .I2(x992), .O(n5821));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5822 (.I0(x981), .I1(x982), .I2(x983), .I3(n5818), .I4(n5819), .O(n5822));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5823 (.I0(x987), .I1(x988), .I2(x989), .I3(n5821), .I4(n5822), .O(n5823));
  LUT3 #(.INIT(8'h96)) lut_n5824 (.I0(n5810), .I1(n5813), .I2(n5814), .O(n5824));
  LUT3 #(.INIT(8'hE8)) lut_n5825 (.I0(n5820), .I1(n5823), .I2(n5824), .O(n5825));
  LUT3 #(.INIT(8'hE8)) lut_n5826 (.I0(x996), .I1(x997), .I2(x998), .O(n5826));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5827 (.I0(x987), .I1(x988), .I2(x989), .I3(n5821), .I4(n5822), .O(n5827));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5828 (.I0(x993), .I1(x994), .I2(x995), .I3(n5826), .I4(n5827), .O(n5828));
  LUT3 #(.INIT(8'hE8)) lut_n5829 (.I0(x1002), .I1(x1003), .I2(x1004), .O(n5829));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5830 (.I0(x993), .I1(x994), .I2(x995), .I3(n5826), .I4(n5827), .O(n5830));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5831 (.I0(x999), .I1(x1000), .I2(x1001), .I3(n5829), .I4(n5830), .O(n5831));
  LUT3 #(.INIT(8'h96)) lut_n5832 (.I0(n5820), .I1(n5823), .I2(n5824), .O(n5832));
  LUT3 #(.INIT(8'hE8)) lut_n5833 (.I0(n5828), .I1(n5831), .I2(n5832), .O(n5833));
  LUT3 #(.INIT(8'h96)) lut_n5834 (.I0(n5807), .I1(n5815), .I2(n5816), .O(n5834));
  LUT3 #(.INIT(8'hE8)) lut_n5835 (.I0(n5825), .I1(n5833), .I2(n5834), .O(n5835));
  LUT3 #(.INIT(8'h96)) lut_n5836 (.I0(n5775), .I1(n5793), .I2(n5794), .O(n5836));
  LUT3 #(.INIT(8'hE8)) lut_n5837 (.I0(n5817), .I1(n5835), .I2(n5836), .O(n5837));
  LUT3 #(.INIT(8'hE8)) lut_n5838 (.I0(x1008), .I1(x1009), .I2(x1010), .O(n5838));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5839 (.I0(x999), .I1(x1000), .I2(x1001), .I3(n5829), .I4(n5830), .O(n5839));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5840 (.I0(x1005), .I1(x1006), .I2(x1007), .I3(n5838), .I4(n5839), .O(n5840));
  LUT3 #(.INIT(8'hE8)) lut_n5841 (.I0(x1014), .I1(x1015), .I2(x1016), .O(n5841));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5842 (.I0(x1005), .I1(x1006), .I2(x1007), .I3(n5838), .I4(n5839), .O(n5842));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5843 (.I0(x1011), .I1(x1012), .I2(x1013), .I3(n5841), .I4(n5842), .O(n5843));
  LUT3 #(.INIT(8'h96)) lut_n5844 (.I0(n5828), .I1(n5831), .I2(n5832), .O(n5844));
  LUT3 #(.INIT(8'hE8)) lut_n5845 (.I0(n5840), .I1(n5843), .I2(n5844), .O(n5845));
  LUT3 #(.INIT(8'hE8)) lut_n5846 (.I0(x1020), .I1(x1021), .I2(x1022), .O(n5846));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5847 (.I0(x1011), .I1(x1012), .I2(x1013), .I3(n5841), .I4(n5842), .O(n5847));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5848 (.I0(x1017), .I1(x1018), .I2(x1019), .I3(n5846), .I4(n5847), .O(n5848));
  LUT3 #(.INIT(8'hE8)) lut_n5849 (.I0(x1026), .I1(x1027), .I2(x1028), .O(n5849));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5850 (.I0(x1017), .I1(x1018), .I2(x1019), .I3(n5846), .I4(n5847), .O(n5850));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5851 (.I0(x1023), .I1(x1024), .I2(x1025), .I3(n5849), .I4(n5850), .O(n5851));
  LUT3 #(.INIT(8'h96)) lut_n5852 (.I0(n5840), .I1(n5843), .I2(n5844), .O(n5852));
  LUT3 #(.INIT(8'hE8)) lut_n5853 (.I0(n5848), .I1(n5851), .I2(n5852), .O(n5853));
  LUT3 #(.INIT(8'h96)) lut_n5854 (.I0(n5825), .I1(n5833), .I2(n5834), .O(n5854));
  LUT3 #(.INIT(8'hE8)) lut_n5855 (.I0(n5845), .I1(n5853), .I2(n5854), .O(n5855));
  LUT3 #(.INIT(8'hE8)) lut_n5856 (.I0(x1032), .I1(x1033), .I2(x1034), .O(n5856));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5857 (.I0(x1023), .I1(x1024), .I2(x1025), .I3(n5849), .I4(n5850), .O(n5857));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5858 (.I0(x1029), .I1(x1030), .I2(x1031), .I3(n5856), .I4(n5857), .O(n5858));
  LUT3 #(.INIT(8'hE8)) lut_n5859 (.I0(x1038), .I1(x1039), .I2(x1040), .O(n5859));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5860 (.I0(x1029), .I1(x1030), .I2(x1031), .I3(n5856), .I4(n5857), .O(n5860));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5861 (.I0(x1035), .I1(x1036), .I2(x1037), .I3(n5859), .I4(n5860), .O(n5861));
  LUT3 #(.INIT(8'h96)) lut_n5862 (.I0(n5848), .I1(n5851), .I2(n5852), .O(n5862));
  LUT3 #(.INIT(8'hE8)) lut_n5863 (.I0(n5858), .I1(n5861), .I2(n5862), .O(n5863));
  LUT3 #(.INIT(8'hE8)) lut_n5864 (.I0(x1044), .I1(x1045), .I2(x1046), .O(n5864));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5865 (.I0(x1035), .I1(x1036), .I2(x1037), .I3(n5859), .I4(n5860), .O(n5865));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5866 (.I0(x1041), .I1(x1042), .I2(x1043), .I3(n5864), .I4(n5865), .O(n5866));
  LUT3 #(.INIT(8'hE8)) lut_n5867 (.I0(x1050), .I1(x1051), .I2(x1052), .O(n5867));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5868 (.I0(x1041), .I1(x1042), .I2(x1043), .I3(n5864), .I4(n5865), .O(n5868));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5869 (.I0(x1047), .I1(x1048), .I2(x1049), .I3(n5867), .I4(n5868), .O(n5869));
  LUT3 #(.INIT(8'h96)) lut_n5870 (.I0(n5858), .I1(n5861), .I2(n5862), .O(n5870));
  LUT3 #(.INIT(8'hE8)) lut_n5871 (.I0(n5866), .I1(n5869), .I2(n5870), .O(n5871));
  LUT3 #(.INIT(8'h96)) lut_n5872 (.I0(n5845), .I1(n5853), .I2(n5854), .O(n5872));
  LUT3 #(.INIT(8'hE8)) lut_n5873 (.I0(n5863), .I1(n5871), .I2(n5872), .O(n5873));
  LUT3 #(.INIT(8'h96)) lut_n5874 (.I0(n5817), .I1(n5835), .I2(n5836), .O(n5874));
  LUT3 #(.INIT(8'hE8)) lut_n5875 (.I0(n5855), .I1(n5873), .I2(n5874), .O(n5875));
  LUT3 #(.INIT(8'h96)) lut_n5876 (.I0(n5757), .I1(n5795), .I2(n5796), .O(n5876));
  LUT3 #(.INIT(8'hE8)) lut_n5877 (.I0(n5837), .I1(n5875), .I2(n5876), .O(n5877));
  LUT3 #(.INIT(8'hE8)) lut_n5878 (.I0(x1056), .I1(x1057), .I2(x1058), .O(n5878));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5879 (.I0(x1047), .I1(x1048), .I2(x1049), .I3(n5867), .I4(n5868), .O(n5879));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5880 (.I0(x1053), .I1(x1054), .I2(x1055), .I3(n5878), .I4(n5879), .O(n5880));
  LUT3 #(.INIT(8'hE8)) lut_n5881 (.I0(x1062), .I1(x1063), .I2(x1064), .O(n5881));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5882 (.I0(x1053), .I1(x1054), .I2(x1055), .I3(n5878), .I4(n5879), .O(n5882));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5883 (.I0(x1059), .I1(x1060), .I2(x1061), .I3(n5881), .I4(n5882), .O(n5883));
  LUT3 #(.INIT(8'h96)) lut_n5884 (.I0(n5866), .I1(n5869), .I2(n5870), .O(n5884));
  LUT3 #(.INIT(8'hE8)) lut_n5885 (.I0(n5880), .I1(n5883), .I2(n5884), .O(n5885));
  LUT3 #(.INIT(8'hE8)) lut_n5886 (.I0(x1068), .I1(x1069), .I2(x1070), .O(n5886));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5887 (.I0(x1059), .I1(x1060), .I2(x1061), .I3(n5881), .I4(n5882), .O(n5887));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5888 (.I0(x1065), .I1(x1066), .I2(x1067), .I3(n5886), .I4(n5887), .O(n5888));
  LUT3 #(.INIT(8'hE8)) lut_n5889 (.I0(x1074), .I1(x1075), .I2(x1076), .O(n5889));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5890 (.I0(x1065), .I1(x1066), .I2(x1067), .I3(n5886), .I4(n5887), .O(n5890));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5891 (.I0(x1071), .I1(x1072), .I2(x1073), .I3(n5889), .I4(n5890), .O(n5891));
  LUT3 #(.INIT(8'h96)) lut_n5892 (.I0(n5880), .I1(n5883), .I2(n5884), .O(n5892));
  LUT3 #(.INIT(8'hE8)) lut_n5893 (.I0(n5888), .I1(n5891), .I2(n5892), .O(n5893));
  LUT3 #(.INIT(8'h96)) lut_n5894 (.I0(n5863), .I1(n5871), .I2(n5872), .O(n5894));
  LUT3 #(.INIT(8'hE8)) lut_n5895 (.I0(n5885), .I1(n5893), .I2(n5894), .O(n5895));
  LUT3 #(.INIT(8'hE8)) lut_n5896 (.I0(x1080), .I1(x1081), .I2(x1082), .O(n5896));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5897 (.I0(x1071), .I1(x1072), .I2(x1073), .I3(n5889), .I4(n5890), .O(n5897));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5898 (.I0(x1077), .I1(x1078), .I2(x1079), .I3(n5896), .I4(n5897), .O(n5898));
  LUT3 #(.INIT(8'hE8)) lut_n5899 (.I0(x1086), .I1(x1087), .I2(x1088), .O(n5899));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5900 (.I0(x1077), .I1(x1078), .I2(x1079), .I3(n5896), .I4(n5897), .O(n5900));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5901 (.I0(x1083), .I1(x1084), .I2(x1085), .I3(n5899), .I4(n5900), .O(n5901));
  LUT3 #(.INIT(8'h96)) lut_n5902 (.I0(n5888), .I1(n5891), .I2(n5892), .O(n5902));
  LUT3 #(.INIT(8'hE8)) lut_n5903 (.I0(n5898), .I1(n5901), .I2(n5902), .O(n5903));
  LUT3 #(.INIT(8'hE8)) lut_n5904 (.I0(x1092), .I1(x1093), .I2(x1094), .O(n5904));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5905 (.I0(x1083), .I1(x1084), .I2(x1085), .I3(n5899), .I4(n5900), .O(n5905));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5906 (.I0(x1089), .I1(x1090), .I2(x1091), .I3(n5904), .I4(n5905), .O(n5906));
  LUT3 #(.INIT(8'hE8)) lut_n5907 (.I0(x1098), .I1(x1099), .I2(x1100), .O(n5907));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5908 (.I0(x1089), .I1(x1090), .I2(x1091), .I3(n5904), .I4(n5905), .O(n5908));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5909 (.I0(x1095), .I1(x1096), .I2(x1097), .I3(n5907), .I4(n5908), .O(n5909));
  LUT3 #(.INIT(8'h96)) lut_n5910 (.I0(n5898), .I1(n5901), .I2(n5902), .O(n5910));
  LUT3 #(.INIT(8'hE8)) lut_n5911 (.I0(n5906), .I1(n5909), .I2(n5910), .O(n5911));
  LUT3 #(.INIT(8'h96)) lut_n5912 (.I0(n5885), .I1(n5893), .I2(n5894), .O(n5912));
  LUT3 #(.INIT(8'hE8)) lut_n5913 (.I0(n5903), .I1(n5911), .I2(n5912), .O(n5913));
  LUT3 #(.INIT(8'h96)) lut_n5914 (.I0(n5855), .I1(n5873), .I2(n5874), .O(n5914));
  LUT3 #(.INIT(8'hE8)) lut_n5915 (.I0(n5895), .I1(n5913), .I2(n5914), .O(n5915));
  LUT3 #(.INIT(8'hE8)) lut_n5916 (.I0(x1104), .I1(x1105), .I2(x1106), .O(n5916));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5917 (.I0(x1095), .I1(x1096), .I2(x1097), .I3(n5907), .I4(n5908), .O(n5917));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5918 (.I0(x1101), .I1(x1102), .I2(x1103), .I3(n5916), .I4(n5917), .O(n5918));
  LUT3 #(.INIT(8'hE8)) lut_n5919 (.I0(x1110), .I1(x1111), .I2(x1112), .O(n5919));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5920 (.I0(x1101), .I1(x1102), .I2(x1103), .I3(n5916), .I4(n5917), .O(n5920));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5921 (.I0(x1107), .I1(x1108), .I2(x1109), .I3(n5919), .I4(n5920), .O(n5921));
  LUT3 #(.INIT(8'h96)) lut_n5922 (.I0(n5906), .I1(n5909), .I2(n5910), .O(n5922));
  LUT3 #(.INIT(8'hE8)) lut_n5923 (.I0(n5918), .I1(n5921), .I2(n5922), .O(n5923));
  LUT3 #(.INIT(8'hE8)) lut_n5924 (.I0(x1116), .I1(x1117), .I2(x1118), .O(n5924));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5925 (.I0(x1107), .I1(x1108), .I2(x1109), .I3(n5919), .I4(n5920), .O(n5925));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5926 (.I0(x1113), .I1(x1114), .I2(x1115), .I3(n5924), .I4(n5925), .O(n5926));
  LUT3 #(.INIT(8'hE8)) lut_n5927 (.I0(x1122), .I1(x1123), .I2(x1124), .O(n5927));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5928 (.I0(x1113), .I1(x1114), .I2(x1115), .I3(n5924), .I4(n5925), .O(n5928));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5929 (.I0(x1119), .I1(x1120), .I2(x1121), .I3(n5927), .I4(n5928), .O(n5929));
  LUT3 #(.INIT(8'h96)) lut_n5930 (.I0(n5918), .I1(n5921), .I2(n5922), .O(n5930));
  LUT3 #(.INIT(8'hE8)) lut_n5931 (.I0(n5926), .I1(n5929), .I2(n5930), .O(n5931));
  LUT3 #(.INIT(8'h96)) lut_n5932 (.I0(n5903), .I1(n5911), .I2(n5912), .O(n5932));
  LUT3 #(.INIT(8'hE8)) lut_n5933 (.I0(n5923), .I1(n5931), .I2(n5932), .O(n5933));
  LUT3 #(.INIT(8'hE8)) lut_n5934 (.I0(x1128), .I1(x1129), .I2(x1130), .O(n5934));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5935 (.I0(x1119), .I1(x1120), .I2(x1121), .I3(n5927), .I4(n5928), .O(n5935));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5936 (.I0(x1125), .I1(x1126), .I2(x1127), .I3(n5934), .I4(n5935), .O(n5936));
  LUT3 #(.INIT(8'hE8)) lut_n5937 (.I0(x1134), .I1(x1135), .I2(x1136), .O(n5937));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5938 (.I0(x1125), .I1(x1126), .I2(x1127), .I3(n5934), .I4(n5935), .O(n5938));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5939 (.I0(x1131), .I1(x1132), .I2(x1133), .I3(n5937), .I4(n5938), .O(n5939));
  LUT3 #(.INIT(8'h96)) lut_n5940 (.I0(n5926), .I1(n5929), .I2(n5930), .O(n5940));
  LUT3 #(.INIT(8'hE8)) lut_n5941 (.I0(n5936), .I1(n5939), .I2(n5940), .O(n5941));
  LUT3 #(.INIT(8'hE8)) lut_n5942 (.I0(x1140), .I1(x1141), .I2(x1142), .O(n5942));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5943 (.I0(x1131), .I1(x1132), .I2(x1133), .I3(n5937), .I4(n5938), .O(n5943));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5944 (.I0(x1137), .I1(x1138), .I2(x1139), .I3(n5942), .I4(n5943), .O(n5944));
  LUT3 #(.INIT(8'hE8)) lut_n5945 (.I0(x1146), .I1(x1147), .I2(x1148), .O(n5945));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5946 (.I0(x1137), .I1(x1138), .I2(x1139), .I3(n5942), .I4(n5943), .O(n5946));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5947 (.I0(x1143), .I1(x1144), .I2(x1145), .I3(n5945), .I4(n5946), .O(n5947));
  LUT3 #(.INIT(8'h96)) lut_n5948 (.I0(n5936), .I1(n5939), .I2(n5940), .O(n5948));
  LUT3 #(.INIT(8'hE8)) lut_n5949 (.I0(n5944), .I1(n5947), .I2(n5948), .O(n5949));
  LUT3 #(.INIT(8'h96)) lut_n5950 (.I0(n5923), .I1(n5931), .I2(n5932), .O(n5950));
  LUT3 #(.INIT(8'hE8)) lut_n5951 (.I0(n5941), .I1(n5949), .I2(n5950), .O(n5951));
  LUT3 #(.INIT(8'h96)) lut_n5952 (.I0(n5895), .I1(n5913), .I2(n5914), .O(n5952));
  LUT3 #(.INIT(8'hE8)) lut_n5953 (.I0(n5933), .I1(n5951), .I2(n5952), .O(n5953));
  LUT3 #(.INIT(8'h96)) lut_n5954 (.I0(n5837), .I1(n5875), .I2(n5876), .O(n5954));
  LUT3 #(.INIT(8'hE8)) lut_n5955 (.I0(n5915), .I1(n5953), .I2(n5954), .O(n5955));
  LUT3 #(.INIT(8'h96)) lut_n5956 (.I0(n5719), .I1(n5797), .I2(n5798), .O(n5956));
  LUT3 #(.INIT(8'hE8)) lut_n5957 (.I0(n5877), .I1(n5955), .I2(n5956), .O(n5957));
  LUT3 #(.INIT(8'h96)) lut_n5958 (.I0(n5324), .I1(n5482), .I2(n5640), .O(n5958));
  LUT3 #(.INIT(8'hE8)) lut_n5959 (.I0(n5799), .I1(n5957), .I2(n5958), .O(n5959));
  LUT3 #(.INIT(8'hE8)) lut_n5960 (.I0(x1152), .I1(x1153), .I2(x1154), .O(n5960));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5961 (.I0(x1143), .I1(x1144), .I2(x1145), .I3(n5945), .I4(n5946), .O(n5961));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5962 (.I0(x1149), .I1(x1150), .I2(x1151), .I3(n5960), .I4(n5961), .O(n5962));
  LUT3 #(.INIT(8'hE8)) lut_n5963 (.I0(x1158), .I1(x1159), .I2(x1160), .O(n5963));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5964 (.I0(x1149), .I1(x1150), .I2(x1151), .I3(n5960), .I4(n5961), .O(n5964));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5965 (.I0(x1155), .I1(x1156), .I2(x1157), .I3(n5963), .I4(n5964), .O(n5965));
  LUT3 #(.INIT(8'h96)) lut_n5966 (.I0(n5944), .I1(n5947), .I2(n5948), .O(n5966));
  LUT3 #(.INIT(8'hE8)) lut_n5967 (.I0(n5962), .I1(n5965), .I2(n5966), .O(n5967));
  LUT3 #(.INIT(8'hE8)) lut_n5968 (.I0(x1164), .I1(x1165), .I2(x1166), .O(n5968));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5969 (.I0(x1155), .I1(x1156), .I2(x1157), .I3(n5963), .I4(n5964), .O(n5969));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5970 (.I0(x1161), .I1(x1162), .I2(x1163), .I3(n5968), .I4(n5969), .O(n5970));
  LUT3 #(.INIT(8'hE8)) lut_n5971 (.I0(x1170), .I1(x1171), .I2(x1172), .O(n5971));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5972 (.I0(x1161), .I1(x1162), .I2(x1163), .I3(n5968), .I4(n5969), .O(n5972));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5973 (.I0(x1167), .I1(x1168), .I2(x1169), .I3(n5971), .I4(n5972), .O(n5973));
  LUT3 #(.INIT(8'h96)) lut_n5974 (.I0(n5962), .I1(n5965), .I2(n5966), .O(n5974));
  LUT3 #(.INIT(8'hE8)) lut_n5975 (.I0(n5970), .I1(n5973), .I2(n5974), .O(n5975));
  LUT3 #(.INIT(8'h96)) lut_n5976 (.I0(n5941), .I1(n5949), .I2(n5950), .O(n5976));
  LUT3 #(.INIT(8'hE8)) lut_n5977 (.I0(n5967), .I1(n5975), .I2(n5976), .O(n5977));
  LUT3 #(.INIT(8'hE8)) lut_n5978 (.I0(x1176), .I1(x1177), .I2(x1178), .O(n5978));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5979 (.I0(x1167), .I1(x1168), .I2(x1169), .I3(n5971), .I4(n5972), .O(n5979));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5980 (.I0(x1173), .I1(x1174), .I2(x1175), .I3(n5978), .I4(n5979), .O(n5980));
  LUT3 #(.INIT(8'hE8)) lut_n5981 (.I0(x1182), .I1(x1183), .I2(x1184), .O(n5981));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5982 (.I0(x1173), .I1(x1174), .I2(x1175), .I3(n5978), .I4(n5979), .O(n5982));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5983 (.I0(x1179), .I1(x1180), .I2(x1181), .I3(n5981), .I4(n5982), .O(n5983));
  LUT3 #(.INIT(8'h96)) lut_n5984 (.I0(n5970), .I1(n5973), .I2(n5974), .O(n5984));
  LUT3 #(.INIT(8'hE8)) lut_n5985 (.I0(n5980), .I1(n5983), .I2(n5984), .O(n5985));
  LUT3 #(.INIT(8'hE8)) lut_n5986 (.I0(x1188), .I1(x1189), .I2(x1190), .O(n5986));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5987 (.I0(x1179), .I1(x1180), .I2(x1181), .I3(n5981), .I4(n5982), .O(n5987));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5988 (.I0(x1185), .I1(x1186), .I2(x1187), .I3(n5986), .I4(n5987), .O(n5988));
  LUT3 #(.INIT(8'hE8)) lut_n5989 (.I0(x1194), .I1(x1195), .I2(x1196), .O(n5989));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5990 (.I0(x1185), .I1(x1186), .I2(x1187), .I3(n5986), .I4(n5987), .O(n5990));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n5991 (.I0(x1191), .I1(x1192), .I2(x1193), .I3(n5989), .I4(n5990), .O(n5991));
  LUT3 #(.INIT(8'h96)) lut_n5992 (.I0(n5980), .I1(n5983), .I2(n5984), .O(n5992));
  LUT3 #(.INIT(8'hE8)) lut_n5993 (.I0(n5988), .I1(n5991), .I2(n5992), .O(n5993));
  LUT3 #(.INIT(8'h96)) lut_n5994 (.I0(n5967), .I1(n5975), .I2(n5976), .O(n5994));
  LUT3 #(.INIT(8'hE8)) lut_n5995 (.I0(n5985), .I1(n5993), .I2(n5994), .O(n5995));
  LUT3 #(.INIT(8'h96)) lut_n5996 (.I0(n5933), .I1(n5951), .I2(n5952), .O(n5996));
  LUT3 #(.INIT(8'hE8)) lut_n5997 (.I0(n5977), .I1(n5995), .I2(n5996), .O(n5997));
  LUT3 #(.INIT(8'hE8)) lut_n5998 (.I0(x1200), .I1(x1201), .I2(x1202), .O(n5998));
  LUT5 #(.INIT(32'hE81717E8)) lut_n5999 (.I0(x1191), .I1(x1192), .I2(x1193), .I3(n5989), .I4(n5990), .O(n5999));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6000 (.I0(x1197), .I1(x1198), .I2(x1199), .I3(n5998), .I4(n5999), .O(n6000));
  LUT3 #(.INIT(8'hE8)) lut_n6001 (.I0(x1206), .I1(x1207), .I2(x1208), .O(n6001));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6002 (.I0(x1197), .I1(x1198), .I2(x1199), .I3(n5998), .I4(n5999), .O(n6002));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6003 (.I0(x1203), .I1(x1204), .I2(x1205), .I3(n6001), .I4(n6002), .O(n6003));
  LUT3 #(.INIT(8'h96)) lut_n6004 (.I0(n5988), .I1(n5991), .I2(n5992), .O(n6004));
  LUT3 #(.INIT(8'hE8)) lut_n6005 (.I0(n6000), .I1(n6003), .I2(n6004), .O(n6005));
  LUT3 #(.INIT(8'hE8)) lut_n6006 (.I0(x1212), .I1(x1213), .I2(x1214), .O(n6006));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6007 (.I0(x1203), .I1(x1204), .I2(x1205), .I3(n6001), .I4(n6002), .O(n6007));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6008 (.I0(x1209), .I1(x1210), .I2(x1211), .I3(n6006), .I4(n6007), .O(n6008));
  LUT3 #(.INIT(8'hE8)) lut_n6009 (.I0(x1218), .I1(x1219), .I2(x1220), .O(n6009));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6010 (.I0(x1209), .I1(x1210), .I2(x1211), .I3(n6006), .I4(n6007), .O(n6010));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6011 (.I0(x1215), .I1(x1216), .I2(x1217), .I3(n6009), .I4(n6010), .O(n6011));
  LUT3 #(.INIT(8'h96)) lut_n6012 (.I0(n6000), .I1(n6003), .I2(n6004), .O(n6012));
  LUT3 #(.INIT(8'hE8)) lut_n6013 (.I0(n6008), .I1(n6011), .I2(n6012), .O(n6013));
  LUT3 #(.INIT(8'h96)) lut_n6014 (.I0(n5985), .I1(n5993), .I2(n5994), .O(n6014));
  LUT3 #(.INIT(8'hE8)) lut_n6015 (.I0(n6005), .I1(n6013), .I2(n6014), .O(n6015));
  LUT3 #(.INIT(8'hE8)) lut_n6016 (.I0(x1224), .I1(x1225), .I2(x1226), .O(n6016));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6017 (.I0(x1215), .I1(x1216), .I2(x1217), .I3(n6009), .I4(n6010), .O(n6017));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6018 (.I0(x1221), .I1(x1222), .I2(x1223), .I3(n6016), .I4(n6017), .O(n6018));
  LUT3 #(.INIT(8'hE8)) lut_n6019 (.I0(x1230), .I1(x1231), .I2(x1232), .O(n6019));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6020 (.I0(x1221), .I1(x1222), .I2(x1223), .I3(n6016), .I4(n6017), .O(n6020));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6021 (.I0(x1227), .I1(x1228), .I2(x1229), .I3(n6019), .I4(n6020), .O(n6021));
  LUT3 #(.INIT(8'h96)) lut_n6022 (.I0(n6008), .I1(n6011), .I2(n6012), .O(n6022));
  LUT3 #(.INIT(8'hE8)) lut_n6023 (.I0(n6018), .I1(n6021), .I2(n6022), .O(n6023));
  LUT3 #(.INIT(8'hE8)) lut_n6024 (.I0(x1236), .I1(x1237), .I2(x1238), .O(n6024));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6025 (.I0(x1227), .I1(x1228), .I2(x1229), .I3(n6019), .I4(n6020), .O(n6025));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6026 (.I0(x1233), .I1(x1234), .I2(x1235), .I3(n6024), .I4(n6025), .O(n6026));
  LUT3 #(.INIT(8'hE8)) lut_n6027 (.I0(x1242), .I1(x1243), .I2(x1244), .O(n6027));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6028 (.I0(x1233), .I1(x1234), .I2(x1235), .I3(n6024), .I4(n6025), .O(n6028));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6029 (.I0(x1239), .I1(x1240), .I2(x1241), .I3(n6027), .I4(n6028), .O(n6029));
  LUT3 #(.INIT(8'h96)) lut_n6030 (.I0(n6018), .I1(n6021), .I2(n6022), .O(n6030));
  LUT3 #(.INIT(8'hE8)) lut_n6031 (.I0(n6026), .I1(n6029), .I2(n6030), .O(n6031));
  LUT3 #(.INIT(8'h96)) lut_n6032 (.I0(n6005), .I1(n6013), .I2(n6014), .O(n6032));
  LUT3 #(.INIT(8'hE8)) lut_n6033 (.I0(n6023), .I1(n6031), .I2(n6032), .O(n6033));
  LUT3 #(.INIT(8'h96)) lut_n6034 (.I0(n5977), .I1(n5995), .I2(n5996), .O(n6034));
  LUT3 #(.INIT(8'hE8)) lut_n6035 (.I0(n6015), .I1(n6033), .I2(n6034), .O(n6035));
  LUT3 #(.INIT(8'h96)) lut_n6036 (.I0(n5915), .I1(n5953), .I2(n5954), .O(n6036));
  LUT3 #(.INIT(8'hE8)) lut_n6037 (.I0(n5997), .I1(n6035), .I2(n6036), .O(n6037));
  LUT3 #(.INIT(8'hE8)) lut_n6038 (.I0(x1248), .I1(x1249), .I2(x1250), .O(n6038));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6039 (.I0(x1239), .I1(x1240), .I2(x1241), .I3(n6027), .I4(n6028), .O(n6039));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6040 (.I0(x1245), .I1(x1246), .I2(x1247), .I3(n6038), .I4(n6039), .O(n6040));
  LUT3 #(.INIT(8'hE8)) lut_n6041 (.I0(x1254), .I1(x1255), .I2(x1256), .O(n6041));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6042 (.I0(x1245), .I1(x1246), .I2(x1247), .I3(n6038), .I4(n6039), .O(n6042));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6043 (.I0(x1251), .I1(x1252), .I2(x1253), .I3(n6041), .I4(n6042), .O(n6043));
  LUT3 #(.INIT(8'h96)) lut_n6044 (.I0(n6026), .I1(n6029), .I2(n6030), .O(n6044));
  LUT3 #(.INIT(8'hE8)) lut_n6045 (.I0(n6040), .I1(n6043), .I2(n6044), .O(n6045));
  LUT3 #(.INIT(8'hE8)) lut_n6046 (.I0(x1260), .I1(x1261), .I2(x1262), .O(n6046));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6047 (.I0(x1251), .I1(x1252), .I2(x1253), .I3(n6041), .I4(n6042), .O(n6047));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6048 (.I0(x1257), .I1(x1258), .I2(x1259), .I3(n6046), .I4(n6047), .O(n6048));
  LUT3 #(.INIT(8'hE8)) lut_n6049 (.I0(x1266), .I1(x1267), .I2(x1268), .O(n6049));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6050 (.I0(x1257), .I1(x1258), .I2(x1259), .I3(n6046), .I4(n6047), .O(n6050));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6051 (.I0(x1263), .I1(x1264), .I2(x1265), .I3(n6049), .I4(n6050), .O(n6051));
  LUT3 #(.INIT(8'h96)) lut_n6052 (.I0(n6040), .I1(n6043), .I2(n6044), .O(n6052));
  LUT3 #(.INIT(8'hE8)) lut_n6053 (.I0(n6048), .I1(n6051), .I2(n6052), .O(n6053));
  LUT3 #(.INIT(8'h96)) lut_n6054 (.I0(n6023), .I1(n6031), .I2(n6032), .O(n6054));
  LUT3 #(.INIT(8'hE8)) lut_n6055 (.I0(n6045), .I1(n6053), .I2(n6054), .O(n6055));
  LUT3 #(.INIT(8'hE8)) lut_n6056 (.I0(x1272), .I1(x1273), .I2(x1274), .O(n6056));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6057 (.I0(x1263), .I1(x1264), .I2(x1265), .I3(n6049), .I4(n6050), .O(n6057));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6058 (.I0(x1269), .I1(x1270), .I2(x1271), .I3(n6056), .I4(n6057), .O(n6058));
  LUT3 #(.INIT(8'hE8)) lut_n6059 (.I0(x1278), .I1(x1279), .I2(x1280), .O(n6059));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6060 (.I0(x1269), .I1(x1270), .I2(x1271), .I3(n6056), .I4(n6057), .O(n6060));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6061 (.I0(x1275), .I1(x1276), .I2(x1277), .I3(n6059), .I4(n6060), .O(n6061));
  LUT3 #(.INIT(8'h96)) lut_n6062 (.I0(n6048), .I1(n6051), .I2(n6052), .O(n6062));
  LUT3 #(.INIT(8'hE8)) lut_n6063 (.I0(n6058), .I1(n6061), .I2(n6062), .O(n6063));
  LUT3 #(.INIT(8'hE8)) lut_n6064 (.I0(x1284), .I1(x1285), .I2(x1286), .O(n6064));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6065 (.I0(x1275), .I1(x1276), .I2(x1277), .I3(n6059), .I4(n6060), .O(n6065));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6066 (.I0(x1281), .I1(x1282), .I2(x1283), .I3(n6064), .I4(n6065), .O(n6066));
  LUT3 #(.INIT(8'hE8)) lut_n6067 (.I0(x1290), .I1(x1291), .I2(x1292), .O(n6067));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6068 (.I0(x1281), .I1(x1282), .I2(x1283), .I3(n6064), .I4(n6065), .O(n6068));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6069 (.I0(x1287), .I1(x1288), .I2(x1289), .I3(n6067), .I4(n6068), .O(n6069));
  LUT3 #(.INIT(8'h96)) lut_n6070 (.I0(n6058), .I1(n6061), .I2(n6062), .O(n6070));
  LUT3 #(.INIT(8'hE8)) lut_n6071 (.I0(n6066), .I1(n6069), .I2(n6070), .O(n6071));
  LUT3 #(.INIT(8'h96)) lut_n6072 (.I0(n6045), .I1(n6053), .I2(n6054), .O(n6072));
  LUT3 #(.INIT(8'hE8)) lut_n6073 (.I0(n6063), .I1(n6071), .I2(n6072), .O(n6073));
  LUT3 #(.INIT(8'h96)) lut_n6074 (.I0(n6015), .I1(n6033), .I2(n6034), .O(n6074));
  LUT3 #(.INIT(8'hE8)) lut_n6075 (.I0(n6055), .I1(n6073), .I2(n6074), .O(n6075));
  LUT3 #(.INIT(8'hE8)) lut_n6076 (.I0(x1296), .I1(x1297), .I2(x1298), .O(n6076));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6077 (.I0(x1287), .I1(x1288), .I2(x1289), .I3(n6067), .I4(n6068), .O(n6077));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6078 (.I0(x1293), .I1(x1294), .I2(x1295), .I3(n6076), .I4(n6077), .O(n6078));
  LUT3 #(.INIT(8'hE8)) lut_n6079 (.I0(x1302), .I1(x1303), .I2(x1304), .O(n6079));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6080 (.I0(x1293), .I1(x1294), .I2(x1295), .I3(n6076), .I4(n6077), .O(n6080));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6081 (.I0(x1299), .I1(x1300), .I2(x1301), .I3(n6079), .I4(n6080), .O(n6081));
  LUT3 #(.INIT(8'h96)) lut_n6082 (.I0(n6066), .I1(n6069), .I2(n6070), .O(n6082));
  LUT3 #(.INIT(8'hE8)) lut_n6083 (.I0(n6078), .I1(n6081), .I2(n6082), .O(n6083));
  LUT3 #(.INIT(8'hE8)) lut_n6084 (.I0(x1308), .I1(x1309), .I2(x1310), .O(n6084));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6085 (.I0(x1299), .I1(x1300), .I2(x1301), .I3(n6079), .I4(n6080), .O(n6085));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6086 (.I0(x1305), .I1(x1306), .I2(x1307), .I3(n6084), .I4(n6085), .O(n6086));
  LUT3 #(.INIT(8'hE8)) lut_n6087 (.I0(x1314), .I1(x1315), .I2(x1316), .O(n6087));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6088 (.I0(x1305), .I1(x1306), .I2(x1307), .I3(n6084), .I4(n6085), .O(n6088));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6089 (.I0(x1311), .I1(x1312), .I2(x1313), .I3(n6087), .I4(n6088), .O(n6089));
  LUT3 #(.INIT(8'h96)) lut_n6090 (.I0(n6078), .I1(n6081), .I2(n6082), .O(n6090));
  LUT3 #(.INIT(8'hE8)) lut_n6091 (.I0(n6086), .I1(n6089), .I2(n6090), .O(n6091));
  LUT3 #(.INIT(8'h96)) lut_n6092 (.I0(n6063), .I1(n6071), .I2(n6072), .O(n6092));
  LUT3 #(.INIT(8'hE8)) lut_n6093 (.I0(n6083), .I1(n6091), .I2(n6092), .O(n6093));
  LUT3 #(.INIT(8'hE8)) lut_n6094 (.I0(x1320), .I1(x1321), .I2(x1322), .O(n6094));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6095 (.I0(x1311), .I1(x1312), .I2(x1313), .I3(n6087), .I4(n6088), .O(n6095));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6096 (.I0(x1317), .I1(x1318), .I2(x1319), .I3(n6094), .I4(n6095), .O(n6096));
  LUT3 #(.INIT(8'hE8)) lut_n6097 (.I0(x1326), .I1(x1327), .I2(x1328), .O(n6097));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6098 (.I0(x1317), .I1(x1318), .I2(x1319), .I3(n6094), .I4(n6095), .O(n6098));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6099 (.I0(x1323), .I1(x1324), .I2(x1325), .I3(n6097), .I4(n6098), .O(n6099));
  LUT3 #(.INIT(8'h96)) lut_n6100 (.I0(n6086), .I1(n6089), .I2(n6090), .O(n6100));
  LUT3 #(.INIT(8'hE8)) lut_n6101 (.I0(n6096), .I1(n6099), .I2(n6100), .O(n6101));
  LUT3 #(.INIT(8'hE8)) lut_n6102 (.I0(x1332), .I1(x1333), .I2(x1334), .O(n6102));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6103 (.I0(x1323), .I1(x1324), .I2(x1325), .I3(n6097), .I4(n6098), .O(n6103));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6104 (.I0(x1329), .I1(x1330), .I2(x1331), .I3(n6102), .I4(n6103), .O(n6104));
  LUT3 #(.INIT(8'hE8)) lut_n6105 (.I0(x1338), .I1(x1339), .I2(x1340), .O(n6105));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6106 (.I0(x1329), .I1(x1330), .I2(x1331), .I3(n6102), .I4(n6103), .O(n6106));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6107 (.I0(x1335), .I1(x1336), .I2(x1337), .I3(n6105), .I4(n6106), .O(n6107));
  LUT3 #(.INIT(8'h96)) lut_n6108 (.I0(n6096), .I1(n6099), .I2(n6100), .O(n6108));
  LUT3 #(.INIT(8'hE8)) lut_n6109 (.I0(n6104), .I1(n6107), .I2(n6108), .O(n6109));
  LUT3 #(.INIT(8'h96)) lut_n6110 (.I0(n6083), .I1(n6091), .I2(n6092), .O(n6110));
  LUT3 #(.INIT(8'hE8)) lut_n6111 (.I0(n6101), .I1(n6109), .I2(n6110), .O(n6111));
  LUT3 #(.INIT(8'h96)) lut_n6112 (.I0(n6055), .I1(n6073), .I2(n6074), .O(n6112));
  LUT3 #(.INIT(8'hE8)) lut_n6113 (.I0(n6093), .I1(n6111), .I2(n6112), .O(n6113));
  LUT3 #(.INIT(8'h96)) lut_n6114 (.I0(n5997), .I1(n6035), .I2(n6036), .O(n6114));
  LUT3 #(.INIT(8'hE8)) lut_n6115 (.I0(n6075), .I1(n6113), .I2(n6114), .O(n6115));
  LUT3 #(.INIT(8'h96)) lut_n6116 (.I0(n5877), .I1(n5955), .I2(n5956), .O(n6116));
  LUT3 #(.INIT(8'hE8)) lut_n6117 (.I0(n6037), .I1(n6115), .I2(n6116), .O(n6117));
  LUT3 #(.INIT(8'hE8)) lut_n6118 (.I0(x1344), .I1(x1345), .I2(x1346), .O(n6118));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6119 (.I0(x1335), .I1(x1336), .I2(x1337), .I3(n6105), .I4(n6106), .O(n6119));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6120 (.I0(x1341), .I1(x1342), .I2(x1343), .I3(n6118), .I4(n6119), .O(n6120));
  LUT3 #(.INIT(8'hE8)) lut_n6121 (.I0(x1350), .I1(x1351), .I2(x1352), .O(n6121));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6122 (.I0(x1341), .I1(x1342), .I2(x1343), .I3(n6118), .I4(n6119), .O(n6122));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6123 (.I0(x1347), .I1(x1348), .I2(x1349), .I3(n6121), .I4(n6122), .O(n6123));
  LUT3 #(.INIT(8'h96)) lut_n6124 (.I0(n6104), .I1(n6107), .I2(n6108), .O(n6124));
  LUT3 #(.INIT(8'hE8)) lut_n6125 (.I0(n6120), .I1(n6123), .I2(n6124), .O(n6125));
  LUT3 #(.INIT(8'hE8)) lut_n6126 (.I0(x1356), .I1(x1357), .I2(x1358), .O(n6126));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6127 (.I0(x1347), .I1(x1348), .I2(x1349), .I3(n6121), .I4(n6122), .O(n6127));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6128 (.I0(x1353), .I1(x1354), .I2(x1355), .I3(n6126), .I4(n6127), .O(n6128));
  LUT3 #(.INIT(8'hE8)) lut_n6129 (.I0(x1362), .I1(x1363), .I2(x1364), .O(n6129));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6130 (.I0(x1353), .I1(x1354), .I2(x1355), .I3(n6126), .I4(n6127), .O(n6130));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6131 (.I0(x1359), .I1(x1360), .I2(x1361), .I3(n6129), .I4(n6130), .O(n6131));
  LUT3 #(.INIT(8'h96)) lut_n6132 (.I0(n6120), .I1(n6123), .I2(n6124), .O(n6132));
  LUT3 #(.INIT(8'hE8)) lut_n6133 (.I0(n6128), .I1(n6131), .I2(n6132), .O(n6133));
  LUT3 #(.INIT(8'h96)) lut_n6134 (.I0(n6101), .I1(n6109), .I2(n6110), .O(n6134));
  LUT3 #(.INIT(8'hE8)) lut_n6135 (.I0(n6125), .I1(n6133), .I2(n6134), .O(n6135));
  LUT3 #(.INIT(8'hE8)) lut_n6136 (.I0(x1368), .I1(x1369), .I2(x1370), .O(n6136));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6137 (.I0(x1359), .I1(x1360), .I2(x1361), .I3(n6129), .I4(n6130), .O(n6137));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6138 (.I0(x1365), .I1(x1366), .I2(x1367), .I3(n6136), .I4(n6137), .O(n6138));
  LUT3 #(.INIT(8'hE8)) lut_n6139 (.I0(x1374), .I1(x1375), .I2(x1376), .O(n6139));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6140 (.I0(x1365), .I1(x1366), .I2(x1367), .I3(n6136), .I4(n6137), .O(n6140));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6141 (.I0(x1371), .I1(x1372), .I2(x1373), .I3(n6139), .I4(n6140), .O(n6141));
  LUT3 #(.INIT(8'h96)) lut_n6142 (.I0(n6128), .I1(n6131), .I2(n6132), .O(n6142));
  LUT3 #(.INIT(8'hE8)) lut_n6143 (.I0(n6138), .I1(n6141), .I2(n6142), .O(n6143));
  LUT3 #(.INIT(8'hE8)) lut_n6144 (.I0(x1380), .I1(x1381), .I2(x1382), .O(n6144));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6145 (.I0(x1371), .I1(x1372), .I2(x1373), .I3(n6139), .I4(n6140), .O(n6145));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6146 (.I0(x1377), .I1(x1378), .I2(x1379), .I3(n6144), .I4(n6145), .O(n6146));
  LUT3 #(.INIT(8'hE8)) lut_n6147 (.I0(x1386), .I1(x1387), .I2(x1388), .O(n6147));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6148 (.I0(x1377), .I1(x1378), .I2(x1379), .I3(n6144), .I4(n6145), .O(n6148));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6149 (.I0(x1383), .I1(x1384), .I2(x1385), .I3(n6147), .I4(n6148), .O(n6149));
  LUT3 #(.INIT(8'h96)) lut_n6150 (.I0(n6138), .I1(n6141), .I2(n6142), .O(n6150));
  LUT3 #(.INIT(8'hE8)) lut_n6151 (.I0(n6146), .I1(n6149), .I2(n6150), .O(n6151));
  LUT3 #(.INIT(8'h96)) lut_n6152 (.I0(n6125), .I1(n6133), .I2(n6134), .O(n6152));
  LUT3 #(.INIT(8'hE8)) lut_n6153 (.I0(n6143), .I1(n6151), .I2(n6152), .O(n6153));
  LUT3 #(.INIT(8'h96)) lut_n6154 (.I0(n6093), .I1(n6111), .I2(n6112), .O(n6154));
  LUT3 #(.INIT(8'hE8)) lut_n6155 (.I0(n6135), .I1(n6153), .I2(n6154), .O(n6155));
  LUT3 #(.INIT(8'hE8)) lut_n6156 (.I0(x1392), .I1(x1393), .I2(x1394), .O(n6156));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6157 (.I0(x1383), .I1(x1384), .I2(x1385), .I3(n6147), .I4(n6148), .O(n6157));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6158 (.I0(x1389), .I1(x1390), .I2(x1391), .I3(n6156), .I4(n6157), .O(n6158));
  LUT3 #(.INIT(8'hE8)) lut_n6159 (.I0(x1398), .I1(x1399), .I2(x1400), .O(n6159));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6160 (.I0(x1389), .I1(x1390), .I2(x1391), .I3(n6156), .I4(n6157), .O(n6160));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6161 (.I0(x1395), .I1(x1396), .I2(x1397), .I3(n6159), .I4(n6160), .O(n6161));
  LUT3 #(.INIT(8'h96)) lut_n6162 (.I0(n6146), .I1(n6149), .I2(n6150), .O(n6162));
  LUT3 #(.INIT(8'hE8)) lut_n6163 (.I0(n6158), .I1(n6161), .I2(n6162), .O(n6163));
  LUT3 #(.INIT(8'hE8)) lut_n6164 (.I0(x1404), .I1(x1405), .I2(x1406), .O(n6164));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6165 (.I0(x1395), .I1(x1396), .I2(x1397), .I3(n6159), .I4(n6160), .O(n6165));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6166 (.I0(x1401), .I1(x1402), .I2(x1403), .I3(n6164), .I4(n6165), .O(n6166));
  LUT3 #(.INIT(8'hE8)) lut_n6167 (.I0(x1410), .I1(x1411), .I2(x1412), .O(n6167));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6168 (.I0(x1401), .I1(x1402), .I2(x1403), .I3(n6164), .I4(n6165), .O(n6168));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6169 (.I0(x1407), .I1(x1408), .I2(x1409), .I3(n6167), .I4(n6168), .O(n6169));
  LUT3 #(.INIT(8'h96)) lut_n6170 (.I0(n6158), .I1(n6161), .I2(n6162), .O(n6170));
  LUT3 #(.INIT(8'hE8)) lut_n6171 (.I0(n6166), .I1(n6169), .I2(n6170), .O(n6171));
  LUT3 #(.INIT(8'h96)) lut_n6172 (.I0(n6143), .I1(n6151), .I2(n6152), .O(n6172));
  LUT3 #(.INIT(8'hE8)) lut_n6173 (.I0(n6163), .I1(n6171), .I2(n6172), .O(n6173));
  LUT3 #(.INIT(8'hE8)) lut_n6174 (.I0(x1416), .I1(x1417), .I2(x1418), .O(n6174));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6175 (.I0(x1407), .I1(x1408), .I2(x1409), .I3(n6167), .I4(n6168), .O(n6175));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6176 (.I0(x1413), .I1(x1414), .I2(x1415), .I3(n6174), .I4(n6175), .O(n6176));
  LUT3 #(.INIT(8'hE8)) lut_n6177 (.I0(x1422), .I1(x1423), .I2(x1424), .O(n6177));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6178 (.I0(x1413), .I1(x1414), .I2(x1415), .I3(n6174), .I4(n6175), .O(n6178));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6179 (.I0(x1419), .I1(x1420), .I2(x1421), .I3(n6177), .I4(n6178), .O(n6179));
  LUT3 #(.INIT(8'h96)) lut_n6180 (.I0(n6166), .I1(n6169), .I2(n6170), .O(n6180));
  LUT3 #(.INIT(8'hE8)) lut_n6181 (.I0(n6176), .I1(n6179), .I2(n6180), .O(n6181));
  LUT3 #(.INIT(8'hE8)) lut_n6182 (.I0(x1428), .I1(x1429), .I2(x1430), .O(n6182));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6183 (.I0(x1419), .I1(x1420), .I2(x1421), .I3(n6177), .I4(n6178), .O(n6183));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6184 (.I0(x1425), .I1(x1426), .I2(x1427), .I3(n6182), .I4(n6183), .O(n6184));
  LUT3 #(.INIT(8'hE8)) lut_n6185 (.I0(x1434), .I1(x1435), .I2(x1436), .O(n6185));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6186 (.I0(x1425), .I1(x1426), .I2(x1427), .I3(n6182), .I4(n6183), .O(n6186));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6187 (.I0(x1431), .I1(x1432), .I2(x1433), .I3(n6185), .I4(n6186), .O(n6187));
  LUT3 #(.INIT(8'h96)) lut_n6188 (.I0(n6176), .I1(n6179), .I2(n6180), .O(n6188));
  LUT3 #(.INIT(8'hE8)) lut_n6189 (.I0(n6184), .I1(n6187), .I2(n6188), .O(n6189));
  LUT3 #(.INIT(8'h96)) lut_n6190 (.I0(n6163), .I1(n6171), .I2(n6172), .O(n6190));
  LUT3 #(.INIT(8'hE8)) lut_n6191 (.I0(n6181), .I1(n6189), .I2(n6190), .O(n6191));
  LUT3 #(.INIT(8'h96)) lut_n6192 (.I0(n6135), .I1(n6153), .I2(n6154), .O(n6192));
  LUT3 #(.INIT(8'hE8)) lut_n6193 (.I0(n6173), .I1(n6191), .I2(n6192), .O(n6193));
  LUT3 #(.INIT(8'h96)) lut_n6194 (.I0(n6075), .I1(n6113), .I2(n6114), .O(n6194));
  LUT3 #(.INIT(8'hE8)) lut_n6195 (.I0(n6155), .I1(n6193), .I2(n6194), .O(n6195));
  LUT3 #(.INIT(8'hE8)) lut_n6196 (.I0(x1440), .I1(x1441), .I2(x1442), .O(n6196));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6197 (.I0(x1431), .I1(x1432), .I2(x1433), .I3(n6185), .I4(n6186), .O(n6197));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6198 (.I0(x1437), .I1(x1438), .I2(x1439), .I3(n6196), .I4(n6197), .O(n6198));
  LUT3 #(.INIT(8'hE8)) lut_n6199 (.I0(x1446), .I1(x1447), .I2(x1448), .O(n6199));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6200 (.I0(x1437), .I1(x1438), .I2(x1439), .I3(n6196), .I4(n6197), .O(n6200));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6201 (.I0(x1443), .I1(x1444), .I2(x1445), .I3(n6199), .I4(n6200), .O(n6201));
  LUT3 #(.INIT(8'h96)) lut_n6202 (.I0(n6184), .I1(n6187), .I2(n6188), .O(n6202));
  LUT3 #(.INIT(8'hE8)) lut_n6203 (.I0(n6198), .I1(n6201), .I2(n6202), .O(n6203));
  LUT3 #(.INIT(8'hE8)) lut_n6204 (.I0(x1452), .I1(x1453), .I2(x1454), .O(n6204));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6205 (.I0(x1443), .I1(x1444), .I2(x1445), .I3(n6199), .I4(n6200), .O(n6205));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6206 (.I0(x1449), .I1(x1450), .I2(x1451), .I3(n6204), .I4(n6205), .O(n6206));
  LUT3 #(.INIT(8'hE8)) lut_n6207 (.I0(x1458), .I1(x1459), .I2(x1460), .O(n6207));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6208 (.I0(x1449), .I1(x1450), .I2(x1451), .I3(n6204), .I4(n6205), .O(n6208));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6209 (.I0(x1455), .I1(x1456), .I2(x1457), .I3(n6207), .I4(n6208), .O(n6209));
  LUT3 #(.INIT(8'h96)) lut_n6210 (.I0(n6198), .I1(n6201), .I2(n6202), .O(n6210));
  LUT3 #(.INIT(8'hE8)) lut_n6211 (.I0(n6206), .I1(n6209), .I2(n6210), .O(n6211));
  LUT3 #(.INIT(8'h96)) lut_n6212 (.I0(n6181), .I1(n6189), .I2(n6190), .O(n6212));
  LUT3 #(.INIT(8'hE8)) lut_n6213 (.I0(n6203), .I1(n6211), .I2(n6212), .O(n6213));
  LUT3 #(.INIT(8'hE8)) lut_n6214 (.I0(x1464), .I1(x1465), .I2(x1466), .O(n6214));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6215 (.I0(x1455), .I1(x1456), .I2(x1457), .I3(n6207), .I4(n6208), .O(n6215));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6216 (.I0(x1461), .I1(x1462), .I2(x1463), .I3(n6214), .I4(n6215), .O(n6216));
  LUT3 #(.INIT(8'hE8)) lut_n6217 (.I0(x1470), .I1(x1471), .I2(x1472), .O(n6217));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6218 (.I0(x1461), .I1(x1462), .I2(x1463), .I3(n6214), .I4(n6215), .O(n6218));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6219 (.I0(x1467), .I1(x1468), .I2(x1469), .I3(n6217), .I4(n6218), .O(n6219));
  LUT3 #(.INIT(8'h96)) lut_n6220 (.I0(n6206), .I1(n6209), .I2(n6210), .O(n6220));
  LUT3 #(.INIT(8'hE8)) lut_n6221 (.I0(n6216), .I1(n6219), .I2(n6220), .O(n6221));
  LUT3 #(.INIT(8'hE8)) lut_n6222 (.I0(x1476), .I1(x1477), .I2(x1478), .O(n6222));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6223 (.I0(x1467), .I1(x1468), .I2(x1469), .I3(n6217), .I4(n6218), .O(n6223));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6224 (.I0(x1473), .I1(x1474), .I2(x1475), .I3(n6222), .I4(n6223), .O(n6224));
  LUT3 #(.INIT(8'hE8)) lut_n6225 (.I0(x1482), .I1(x1483), .I2(x1484), .O(n6225));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6226 (.I0(x1473), .I1(x1474), .I2(x1475), .I3(n6222), .I4(n6223), .O(n6226));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6227 (.I0(x1479), .I1(x1480), .I2(x1481), .I3(n6225), .I4(n6226), .O(n6227));
  LUT3 #(.INIT(8'h96)) lut_n6228 (.I0(n6216), .I1(n6219), .I2(n6220), .O(n6228));
  LUT3 #(.INIT(8'hE8)) lut_n6229 (.I0(n6224), .I1(n6227), .I2(n6228), .O(n6229));
  LUT3 #(.INIT(8'h96)) lut_n6230 (.I0(n6203), .I1(n6211), .I2(n6212), .O(n6230));
  LUT3 #(.INIT(8'hE8)) lut_n6231 (.I0(n6221), .I1(n6229), .I2(n6230), .O(n6231));
  LUT3 #(.INIT(8'h96)) lut_n6232 (.I0(n6173), .I1(n6191), .I2(n6192), .O(n6232));
  LUT3 #(.INIT(8'hE8)) lut_n6233 (.I0(n6213), .I1(n6231), .I2(n6232), .O(n6233));
  LUT3 #(.INIT(8'hE8)) lut_n6234 (.I0(x1488), .I1(x1489), .I2(x1490), .O(n6234));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6235 (.I0(x1479), .I1(x1480), .I2(x1481), .I3(n6225), .I4(n6226), .O(n6235));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6236 (.I0(x1485), .I1(x1486), .I2(x1487), .I3(n6234), .I4(n6235), .O(n6236));
  LUT3 #(.INIT(8'hE8)) lut_n6237 (.I0(x1494), .I1(x1495), .I2(x1496), .O(n6237));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6238 (.I0(x1485), .I1(x1486), .I2(x1487), .I3(n6234), .I4(n6235), .O(n6238));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6239 (.I0(x1491), .I1(x1492), .I2(x1493), .I3(n6237), .I4(n6238), .O(n6239));
  LUT3 #(.INIT(8'h96)) lut_n6240 (.I0(n6224), .I1(n6227), .I2(n6228), .O(n6240));
  LUT3 #(.INIT(8'hE8)) lut_n6241 (.I0(n6236), .I1(n6239), .I2(n6240), .O(n6241));
  LUT3 #(.INIT(8'hE8)) lut_n6242 (.I0(x1500), .I1(x1501), .I2(x1502), .O(n6242));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6243 (.I0(x1491), .I1(x1492), .I2(x1493), .I3(n6237), .I4(n6238), .O(n6243));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6244 (.I0(x1497), .I1(x1498), .I2(x1499), .I3(n6242), .I4(n6243), .O(n6244));
  LUT3 #(.INIT(8'hE8)) lut_n6245 (.I0(x1506), .I1(x1507), .I2(x1508), .O(n6245));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6246 (.I0(x1497), .I1(x1498), .I2(x1499), .I3(n6242), .I4(n6243), .O(n6246));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6247 (.I0(x1503), .I1(x1504), .I2(x1505), .I3(n6245), .I4(n6246), .O(n6247));
  LUT3 #(.INIT(8'h96)) lut_n6248 (.I0(n6236), .I1(n6239), .I2(n6240), .O(n6248));
  LUT3 #(.INIT(8'hE8)) lut_n6249 (.I0(n6244), .I1(n6247), .I2(n6248), .O(n6249));
  LUT3 #(.INIT(8'h96)) lut_n6250 (.I0(n6221), .I1(n6229), .I2(n6230), .O(n6250));
  LUT3 #(.INIT(8'hE8)) lut_n6251 (.I0(n6241), .I1(n6249), .I2(n6250), .O(n6251));
  LUT3 #(.INIT(8'hE8)) lut_n6252 (.I0(x1512), .I1(x1513), .I2(x1514), .O(n6252));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6253 (.I0(x1503), .I1(x1504), .I2(x1505), .I3(n6245), .I4(n6246), .O(n6253));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6254 (.I0(x1509), .I1(x1510), .I2(x1511), .I3(n6252), .I4(n6253), .O(n6254));
  LUT3 #(.INIT(8'hE8)) lut_n6255 (.I0(x1518), .I1(x1519), .I2(x1520), .O(n6255));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6256 (.I0(x1509), .I1(x1510), .I2(x1511), .I3(n6252), .I4(n6253), .O(n6256));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6257 (.I0(x1515), .I1(x1516), .I2(x1517), .I3(n6255), .I4(n6256), .O(n6257));
  LUT3 #(.INIT(8'h96)) lut_n6258 (.I0(n6244), .I1(n6247), .I2(n6248), .O(n6258));
  LUT3 #(.INIT(8'hE8)) lut_n6259 (.I0(n6254), .I1(n6257), .I2(n6258), .O(n6259));
  LUT3 #(.INIT(8'hE8)) lut_n6260 (.I0(x1524), .I1(x1525), .I2(x1526), .O(n6260));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6261 (.I0(x1515), .I1(x1516), .I2(x1517), .I3(n6255), .I4(n6256), .O(n6261));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6262 (.I0(x1521), .I1(x1522), .I2(x1523), .I3(n6260), .I4(n6261), .O(n6262));
  LUT3 #(.INIT(8'hE8)) lut_n6263 (.I0(x1530), .I1(x1531), .I2(x1532), .O(n6263));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6264 (.I0(x1521), .I1(x1522), .I2(x1523), .I3(n6260), .I4(n6261), .O(n6264));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6265 (.I0(x1527), .I1(x1528), .I2(x1529), .I3(n6263), .I4(n6264), .O(n6265));
  LUT3 #(.INIT(8'h96)) lut_n6266 (.I0(n6254), .I1(n6257), .I2(n6258), .O(n6266));
  LUT3 #(.INIT(8'hE8)) lut_n6267 (.I0(n6262), .I1(n6265), .I2(n6266), .O(n6267));
  LUT3 #(.INIT(8'h96)) lut_n6268 (.I0(n6241), .I1(n6249), .I2(n6250), .O(n6268));
  LUT3 #(.INIT(8'hE8)) lut_n6269 (.I0(n6259), .I1(n6267), .I2(n6268), .O(n6269));
  LUT3 #(.INIT(8'h96)) lut_n6270 (.I0(n6213), .I1(n6231), .I2(n6232), .O(n6270));
  LUT3 #(.INIT(8'hE8)) lut_n6271 (.I0(n6251), .I1(n6269), .I2(n6270), .O(n6271));
  LUT3 #(.INIT(8'h96)) lut_n6272 (.I0(n6155), .I1(n6193), .I2(n6194), .O(n6272));
  LUT3 #(.INIT(8'hE8)) lut_n6273 (.I0(n6233), .I1(n6271), .I2(n6272), .O(n6273));
  LUT3 #(.INIT(8'h96)) lut_n6274 (.I0(n6037), .I1(n6115), .I2(n6116), .O(n6274));
  LUT3 #(.INIT(8'hE8)) lut_n6275 (.I0(n6195), .I1(n6273), .I2(n6274), .O(n6275));
  LUT3 #(.INIT(8'h96)) lut_n6276 (.I0(n5799), .I1(n5957), .I2(n5958), .O(n6276));
  LUT3 #(.INIT(8'hE8)) lut_n6277 (.I0(n6117), .I1(n6275), .I2(n6276), .O(n6277));
  LUT3 #(.INIT(8'hE8)) lut_n6278 (.I0(n5641), .I1(n5959), .I2(n6277), .O(n6278));
  LUT3 #(.INIT(8'hE8)) lut_n6279 (.I0(x1536), .I1(x1537), .I2(x1538), .O(n6279));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6280 (.I0(x1527), .I1(x1528), .I2(x1529), .I3(n6263), .I4(n6264), .O(n6280));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6281 (.I0(x1533), .I1(x1534), .I2(x1535), .I3(n6279), .I4(n6280), .O(n6281));
  LUT3 #(.INIT(8'hE8)) lut_n6282 (.I0(x1542), .I1(x1543), .I2(x1544), .O(n6282));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6283 (.I0(x1533), .I1(x1534), .I2(x1535), .I3(n6279), .I4(n6280), .O(n6283));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6284 (.I0(x1539), .I1(x1540), .I2(x1541), .I3(n6282), .I4(n6283), .O(n6284));
  LUT3 #(.INIT(8'h96)) lut_n6285 (.I0(n6262), .I1(n6265), .I2(n6266), .O(n6285));
  LUT3 #(.INIT(8'hE8)) lut_n6286 (.I0(n6281), .I1(n6284), .I2(n6285), .O(n6286));
  LUT3 #(.INIT(8'hE8)) lut_n6287 (.I0(x1548), .I1(x1549), .I2(x1550), .O(n6287));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6288 (.I0(x1539), .I1(x1540), .I2(x1541), .I3(n6282), .I4(n6283), .O(n6288));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6289 (.I0(x1545), .I1(x1546), .I2(x1547), .I3(n6287), .I4(n6288), .O(n6289));
  LUT3 #(.INIT(8'hE8)) lut_n6290 (.I0(x1554), .I1(x1555), .I2(x1556), .O(n6290));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6291 (.I0(x1545), .I1(x1546), .I2(x1547), .I3(n6287), .I4(n6288), .O(n6291));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6292 (.I0(x1551), .I1(x1552), .I2(x1553), .I3(n6290), .I4(n6291), .O(n6292));
  LUT3 #(.INIT(8'h96)) lut_n6293 (.I0(n6281), .I1(n6284), .I2(n6285), .O(n6293));
  LUT3 #(.INIT(8'hE8)) lut_n6294 (.I0(n6289), .I1(n6292), .I2(n6293), .O(n6294));
  LUT3 #(.INIT(8'h96)) lut_n6295 (.I0(n6259), .I1(n6267), .I2(n6268), .O(n6295));
  LUT3 #(.INIT(8'hE8)) lut_n6296 (.I0(n6286), .I1(n6294), .I2(n6295), .O(n6296));
  LUT3 #(.INIT(8'hE8)) lut_n6297 (.I0(x1560), .I1(x1561), .I2(x1562), .O(n6297));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6298 (.I0(x1551), .I1(x1552), .I2(x1553), .I3(n6290), .I4(n6291), .O(n6298));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6299 (.I0(x1557), .I1(x1558), .I2(x1559), .I3(n6297), .I4(n6298), .O(n6299));
  LUT3 #(.INIT(8'hE8)) lut_n6300 (.I0(x1566), .I1(x1567), .I2(x1568), .O(n6300));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6301 (.I0(x1557), .I1(x1558), .I2(x1559), .I3(n6297), .I4(n6298), .O(n6301));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6302 (.I0(x1563), .I1(x1564), .I2(x1565), .I3(n6300), .I4(n6301), .O(n6302));
  LUT3 #(.INIT(8'h96)) lut_n6303 (.I0(n6289), .I1(n6292), .I2(n6293), .O(n6303));
  LUT3 #(.INIT(8'hE8)) lut_n6304 (.I0(n6299), .I1(n6302), .I2(n6303), .O(n6304));
  LUT3 #(.INIT(8'hE8)) lut_n6305 (.I0(x1572), .I1(x1573), .I2(x1574), .O(n6305));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6306 (.I0(x1563), .I1(x1564), .I2(x1565), .I3(n6300), .I4(n6301), .O(n6306));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6307 (.I0(x1569), .I1(x1570), .I2(x1571), .I3(n6305), .I4(n6306), .O(n6307));
  LUT3 #(.INIT(8'hE8)) lut_n6308 (.I0(x1578), .I1(x1579), .I2(x1580), .O(n6308));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6309 (.I0(x1569), .I1(x1570), .I2(x1571), .I3(n6305), .I4(n6306), .O(n6309));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6310 (.I0(x1575), .I1(x1576), .I2(x1577), .I3(n6308), .I4(n6309), .O(n6310));
  LUT3 #(.INIT(8'h96)) lut_n6311 (.I0(n6299), .I1(n6302), .I2(n6303), .O(n6311));
  LUT3 #(.INIT(8'hE8)) lut_n6312 (.I0(n6307), .I1(n6310), .I2(n6311), .O(n6312));
  LUT3 #(.INIT(8'h96)) lut_n6313 (.I0(n6286), .I1(n6294), .I2(n6295), .O(n6313));
  LUT3 #(.INIT(8'hE8)) lut_n6314 (.I0(n6304), .I1(n6312), .I2(n6313), .O(n6314));
  LUT3 #(.INIT(8'h96)) lut_n6315 (.I0(n6251), .I1(n6269), .I2(n6270), .O(n6315));
  LUT3 #(.INIT(8'hE8)) lut_n6316 (.I0(n6296), .I1(n6314), .I2(n6315), .O(n6316));
  LUT3 #(.INIT(8'hE8)) lut_n6317 (.I0(x1584), .I1(x1585), .I2(x1586), .O(n6317));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6318 (.I0(x1575), .I1(x1576), .I2(x1577), .I3(n6308), .I4(n6309), .O(n6318));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6319 (.I0(x1581), .I1(x1582), .I2(x1583), .I3(n6317), .I4(n6318), .O(n6319));
  LUT3 #(.INIT(8'hE8)) lut_n6320 (.I0(x1590), .I1(x1591), .I2(x1592), .O(n6320));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6321 (.I0(x1581), .I1(x1582), .I2(x1583), .I3(n6317), .I4(n6318), .O(n6321));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6322 (.I0(x1587), .I1(x1588), .I2(x1589), .I3(n6320), .I4(n6321), .O(n6322));
  LUT3 #(.INIT(8'h96)) lut_n6323 (.I0(n6307), .I1(n6310), .I2(n6311), .O(n6323));
  LUT3 #(.INIT(8'hE8)) lut_n6324 (.I0(n6319), .I1(n6322), .I2(n6323), .O(n6324));
  LUT3 #(.INIT(8'hE8)) lut_n6325 (.I0(x1596), .I1(x1597), .I2(x1598), .O(n6325));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6326 (.I0(x1587), .I1(x1588), .I2(x1589), .I3(n6320), .I4(n6321), .O(n6326));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6327 (.I0(x1593), .I1(x1594), .I2(x1595), .I3(n6325), .I4(n6326), .O(n6327));
  LUT3 #(.INIT(8'hE8)) lut_n6328 (.I0(x1602), .I1(x1603), .I2(x1604), .O(n6328));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6329 (.I0(x1593), .I1(x1594), .I2(x1595), .I3(n6325), .I4(n6326), .O(n6329));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6330 (.I0(x1599), .I1(x1600), .I2(x1601), .I3(n6328), .I4(n6329), .O(n6330));
  LUT3 #(.INIT(8'h96)) lut_n6331 (.I0(n6319), .I1(n6322), .I2(n6323), .O(n6331));
  LUT3 #(.INIT(8'hE8)) lut_n6332 (.I0(n6327), .I1(n6330), .I2(n6331), .O(n6332));
  LUT3 #(.INIT(8'h96)) lut_n6333 (.I0(n6304), .I1(n6312), .I2(n6313), .O(n6333));
  LUT3 #(.INIT(8'hE8)) lut_n6334 (.I0(n6324), .I1(n6332), .I2(n6333), .O(n6334));
  LUT3 #(.INIT(8'hE8)) lut_n6335 (.I0(x1608), .I1(x1609), .I2(x1610), .O(n6335));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6336 (.I0(x1599), .I1(x1600), .I2(x1601), .I3(n6328), .I4(n6329), .O(n6336));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6337 (.I0(x1605), .I1(x1606), .I2(x1607), .I3(n6335), .I4(n6336), .O(n6337));
  LUT3 #(.INIT(8'hE8)) lut_n6338 (.I0(x1614), .I1(x1615), .I2(x1616), .O(n6338));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6339 (.I0(x1605), .I1(x1606), .I2(x1607), .I3(n6335), .I4(n6336), .O(n6339));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6340 (.I0(x1611), .I1(x1612), .I2(x1613), .I3(n6338), .I4(n6339), .O(n6340));
  LUT3 #(.INIT(8'h96)) lut_n6341 (.I0(n6327), .I1(n6330), .I2(n6331), .O(n6341));
  LUT3 #(.INIT(8'hE8)) lut_n6342 (.I0(n6337), .I1(n6340), .I2(n6341), .O(n6342));
  LUT3 #(.INIT(8'hE8)) lut_n6343 (.I0(x1620), .I1(x1621), .I2(x1622), .O(n6343));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6344 (.I0(x1611), .I1(x1612), .I2(x1613), .I3(n6338), .I4(n6339), .O(n6344));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6345 (.I0(x1617), .I1(x1618), .I2(x1619), .I3(n6343), .I4(n6344), .O(n6345));
  LUT3 #(.INIT(8'hE8)) lut_n6346 (.I0(x1626), .I1(x1627), .I2(x1628), .O(n6346));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6347 (.I0(x1617), .I1(x1618), .I2(x1619), .I3(n6343), .I4(n6344), .O(n6347));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6348 (.I0(x1623), .I1(x1624), .I2(x1625), .I3(n6346), .I4(n6347), .O(n6348));
  LUT3 #(.INIT(8'h96)) lut_n6349 (.I0(n6337), .I1(n6340), .I2(n6341), .O(n6349));
  LUT3 #(.INIT(8'hE8)) lut_n6350 (.I0(n6345), .I1(n6348), .I2(n6349), .O(n6350));
  LUT3 #(.INIT(8'h96)) lut_n6351 (.I0(n6324), .I1(n6332), .I2(n6333), .O(n6351));
  LUT3 #(.INIT(8'hE8)) lut_n6352 (.I0(n6342), .I1(n6350), .I2(n6351), .O(n6352));
  LUT3 #(.INIT(8'h96)) lut_n6353 (.I0(n6296), .I1(n6314), .I2(n6315), .O(n6353));
  LUT3 #(.INIT(8'hE8)) lut_n6354 (.I0(n6334), .I1(n6352), .I2(n6353), .O(n6354));
  LUT3 #(.INIT(8'h96)) lut_n6355 (.I0(n6233), .I1(n6271), .I2(n6272), .O(n6355));
  LUT3 #(.INIT(8'hE8)) lut_n6356 (.I0(n6316), .I1(n6354), .I2(n6355), .O(n6356));
  LUT3 #(.INIT(8'hE8)) lut_n6357 (.I0(x1632), .I1(x1633), .I2(x1634), .O(n6357));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6358 (.I0(x1623), .I1(x1624), .I2(x1625), .I3(n6346), .I4(n6347), .O(n6358));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6359 (.I0(x1629), .I1(x1630), .I2(x1631), .I3(n6357), .I4(n6358), .O(n6359));
  LUT3 #(.INIT(8'hE8)) lut_n6360 (.I0(x1638), .I1(x1639), .I2(x1640), .O(n6360));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6361 (.I0(x1629), .I1(x1630), .I2(x1631), .I3(n6357), .I4(n6358), .O(n6361));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6362 (.I0(x1635), .I1(x1636), .I2(x1637), .I3(n6360), .I4(n6361), .O(n6362));
  LUT3 #(.INIT(8'h96)) lut_n6363 (.I0(n6345), .I1(n6348), .I2(n6349), .O(n6363));
  LUT3 #(.INIT(8'hE8)) lut_n6364 (.I0(n6359), .I1(n6362), .I2(n6363), .O(n6364));
  LUT3 #(.INIT(8'hE8)) lut_n6365 (.I0(x1644), .I1(x1645), .I2(x1646), .O(n6365));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6366 (.I0(x1635), .I1(x1636), .I2(x1637), .I3(n6360), .I4(n6361), .O(n6366));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6367 (.I0(x1641), .I1(x1642), .I2(x1643), .I3(n6365), .I4(n6366), .O(n6367));
  LUT3 #(.INIT(8'hE8)) lut_n6368 (.I0(x1650), .I1(x1651), .I2(x1652), .O(n6368));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6369 (.I0(x1641), .I1(x1642), .I2(x1643), .I3(n6365), .I4(n6366), .O(n6369));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6370 (.I0(x1647), .I1(x1648), .I2(x1649), .I3(n6368), .I4(n6369), .O(n6370));
  LUT3 #(.INIT(8'h96)) lut_n6371 (.I0(n6359), .I1(n6362), .I2(n6363), .O(n6371));
  LUT3 #(.INIT(8'hE8)) lut_n6372 (.I0(n6367), .I1(n6370), .I2(n6371), .O(n6372));
  LUT3 #(.INIT(8'h96)) lut_n6373 (.I0(n6342), .I1(n6350), .I2(n6351), .O(n6373));
  LUT3 #(.INIT(8'hE8)) lut_n6374 (.I0(n6364), .I1(n6372), .I2(n6373), .O(n6374));
  LUT3 #(.INIT(8'hE8)) lut_n6375 (.I0(x1656), .I1(x1657), .I2(x1658), .O(n6375));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6376 (.I0(x1647), .I1(x1648), .I2(x1649), .I3(n6368), .I4(n6369), .O(n6376));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6377 (.I0(x1653), .I1(x1654), .I2(x1655), .I3(n6375), .I4(n6376), .O(n6377));
  LUT3 #(.INIT(8'hE8)) lut_n6378 (.I0(x1662), .I1(x1663), .I2(x1664), .O(n6378));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6379 (.I0(x1653), .I1(x1654), .I2(x1655), .I3(n6375), .I4(n6376), .O(n6379));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6380 (.I0(x1659), .I1(x1660), .I2(x1661), .I3(n6378), .I4(n6379), .O(n6380));
  LUT3 #(.INIT(8'h96)) lut_n6381 (.I0(n6367), .I1(n6370), .I2(n6371), .O(n6381));
  LUT3 #(.INIT(8'hE8)) lut_n6382 (.I0(n6377), .I1(n6380), .I2(n6381), .O(n6382));
  LUT3 #(.INIT(8'hE8)) lut_n6383 (.I0(x1668), .I1(x1669), .I2(x1670), .O(n6383));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6384 (.I0(x1659), .I1(x1660), .I2(x1661), .I3(n6378), .I4(n6379), .O(n6384));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6385 (.I0(x1665), .I1(x1666), .I2(x1667), .I3(n6383), .I4(n6384), .O(n6385));
  LUT3 #(.INIT(8'hE8)) lut_n6386 (.I0(x1674), .I1(x1675), .I2(x1676), .O(n6386));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6387 (.I0(x1665), .I1(x1666), .I2(x1667), .I3(n6383), .I4(n6384), .O(n6387));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6388 (.I0(x1671), .I1(x1672), .I2(x1673), .I3(n6386), .I4(n6387), .O(n6388));
  LUT3 #(.INIT(8'h96)) lut_n6389 (.I0(n6377), .I1(n6380), .I2(n6381), .O(n6389));
  LUT3 #(.INIT(8'hE8)) lut_n6390 (.I0(n6385), .I1(n6388), .I2(n6389), .O(n6390));
  LUT3 #(.INIT(8'h96)) lut_n6391 (.I0(n6364), .I1(n6372), .I2(n6373), .O(n6391));
  LUT3 #(.INIT(8'hE8)) lut_n6392 (.I0(n6382), .I1(n6390), .I2(n6391), .O(n6392));
  LUT3 #(.INIT(8'h96)) lut_n6393 (.I0(n6334), .I1(n6352), .I2(n6353), .O(n6393));
  LUT3 #(.INIT(8'hE8)) lut_n6394 (.I0(n6374), .I1(n6392), .I2(n6393), .O(n6394));
  LUT3 #(.INIT(8'hE8)) lut_n6395 (.I0(x1680), .I1(x1681), .I2(x1682), .O(n6395));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6396 (.I0(x1671), .I1(x1672), .I2(x1673), .I3(n6386), .I4(n6387), .O(n6396));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6397 (.I0(x1677), .I1(x1678), .I2(x1679), .I3(n6395), .I4(n6396), .O(n6397));
  LUT3 #(.INIT(8'hE8)) lut_n6398 (.I0(x1686), .I1(x1687), .I2(x1688), .O(n6398));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6399 (.I0(x1677), .I1(x1678), .I2(x1679), .I3(n6395), .I4(n6396), .O(n6399));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6400 (.I0(x1683), .I1(x1684), .I2(x1685), .I3(n6398), .I4(n6399), .O(n6400));
  LUT3 #(.INIT(8'h96)) lut_n6401 (.I0(n6385), .I1(n6388), .I2(n6389), .O(n6401));
  LUT3 #(.INIT(8'hE8)) lut_n6402 (.I0(n6397), .I1(n6400), .I2(n6401), .O(n6402));
  LUT3 #(.INIT(8'hE8)) lut_n6403 (.I0(x1692), .I1(x1693), .I2(x1694), .O(n6403));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6404 (.I0(x1683), .I1(x1684), .I2(x1685), .I3(n6398), .I4(n6399), .O(n6404));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6405 (.I0(x1689), .I1(x1690), .I2(x1691), .I3(n6403), .I4(n6404), .O(n6405));
  LUT3 #(.INIT(8'hE8)) lut_n6406 (.I0(x1698), .I1(x1699), .I2(x1700), .O(n6406));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6407 (.I0(x1689), .I1(x1690), .I2(x1691), .I3(n6403), .I4(n6404), .O(n6407));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6408 (.I0(x1695), .I1(x1696), .I2(x1697), .I3(n6406), .I4(n6407), .O(n6408));
  LUT3 #(.INIT(8'h96)) lut_n6409 (.I0(n6397), .I1(n6400), .I2(n6401), .O(n6409));
  LUT3 #(.INIT(8'hE8)) lut_n6410 (.I0(n6405), .I1(n6408), .I2(n6409), .O(n6410));
  LUT3 #(.INIT(8'h96)) lut_n6411 (.I0(n6382), .I1(n6390), .I2(n6391), .O(n6411));
  LUT3 #(.INIT(8'hE8)) lut_n6412 (.I0(n6402), .I1(n6410), .I2(n6411), .O(n6412));
  LUT3 #(.INIT(8'hE8)) lut_n6413 (.I0(x1704), .I1(x1705), .I2(x1706), .O(n6413));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6414 (.I0(x1695), .I1(x1696), .I2(x1697), .I3(n6406), .I4(n6407), .O(n6414));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6415 (.I0(x1701), .I1(x1702), .I2(x1703), .I3(n6413), .I4(n6414), .O(n6415));
  LUT3 #(.INIT(8'hE8)) lut_n6416 (.I0(x1710), .I1(x1711), .I2(x1712), .O(n6416));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6417 (.I0(x1701), .I1(x1702), .I2(x1703), .I3(n6413), .I4(n6414), .O(n6417));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6418 (.I0(x1707), .I1(x1708), .I2(x1709), .I3(n6416), .I4(n6417), .O(n6418));
  LUT3 #(.INIT(8'h96)) lut_n6419 (.I0(n6405), .I1(n6408), .I2(n6409), .O(n6419));
  LUT3 #(.INIT(8'hE8)) lut_n6420 (.I0(n6415), .I1(n6418), .I2(n6419), .O(n6420));
  LUT3 #(.INIT(8'hE8)) lut_n6421 (.I0(x1716), .I1(x1717), .I2(x1718), .O(n6421));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6422 (.I0(x1707), .I1(x1708), .I2(x1709), .I3(n6416), .I4(n6417), .O(n6422));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6423 (.I0(x1713), .I1(x1714), .I2(x1715), .I3(n6421), .I4(n6422), .O(n6423));
  LUT3 #(.INIT(8'hE8)) lut_n6424 (.I0(x1722), .I1(x1723), .I2(x1724), .O(n6424));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6425 (.I0(x1713), .I1(x1714), .I2(x1715), .I3(n6421), .I4(n6422), .O(n6425));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6426 (.I0(x1719), .I1(x1720), .I2(x1721), .I3(n6424), .I4(n6425), .O(n6426));
  LUT3 #(.INIT(8'h96)) lut_n6427 (.I0(n6415), .I1(n6418), .I2(n6419), .O(n6427));
  LUT3 #(.INIT(8'hE8)) lut_n6428 (.I0(n6423), .I1(n6426), .I2(n6427), .O(n6428));
  LUT3 #(.INIT(8'h96)) lut_n6429 (.I0(n6402), .I1(n6410), .I2(n6411), .O(n6429));
  LUT3 #(.INIT(8'hE8)) lut_n6430 (.I0(n6420), .I1(n6428), .I2(n6429), .O(n6430));
  LUT3 #(.INIT(8'h96)) lut_n6431 (.I0(n6374), .I1(n6392), .I2(n6393), .O(n6431));
  LUT3 #(.INIT(8'hE8)) lut_n6432 (.I0(n6412), .I1(n6430), .I2(n6431), .O(n6432));
  LUT3 #(.INIT(8'h96)) lut_n6433 (.I0(n6316), .I1(n6354), .I2(n6355), .O(n6433));
  LUT3 #(.INIT(8'hE8)) lut_n6434 (.I0(n6394), .I1(n6432), .I2(n6433), .O(n6434));
  LUT3 #(.INIT(8'h96)) lut_n6435 (.I0(n6195), .I1(n6273), .I2(n6274), .O(n6435));
  LUT3 #(.INIT(8'hE8)) lut_n6436 (.I0(n6356), .I1(n6434), .I2(n6435), .O(n6436));
  LUT3 #(.INIT(8'hE8)) lut_n6437 (.I0(x1728), .I1(x1729), .I2(x1730), .O(n6437));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6438 (.I0(x1719), .I1(x1720), .I2(x1721), .I3(n6424), .I4(n6425), .O(n6438));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6439 (.I0(x1725), .I1(x1726), .I2(x1727), .I3(n6437), .I4(n6438), .O(n6439));
  LUT3 #(.INIT(8'hE8)) lut_n6440 (.I0(x1734), .I1(x1735), .I2(x1736), .O(n6440));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6441 (.I0(x1725), .I1(x1726), .I2(x1727), .I3(n6437), .I4(n6438), .O(n6441));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6442 (.I0(x1731), .I1(x1732), .I2(x1733), .I3(n6440), .I4(n6441), .O(n6442));
  LUT3 #(.INIT(8'h96)) lut_n6443 (.I0(n6423), .I1(n6426), .I2(n6427), .O(n6443));
  LUT3 #(.INIT(8'hE8)) lut_n6444 (.I0(n6439), .I1(n6442), .I2(n6443), .O(n6444));
  LUT3 #(.INIT(8'hE8)) lut_n6445 (.I0(x1740), .I1(x1741), .I2(x1742), .O(n6445));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6446 (.I0(x1731), .I1(x1732), .I2(x1733), .I3(n6440), .I4(n6441), .O(n6446));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6447 (.I0(x1737), .I1(x1738), .I2(x1739), .I3(n6445), .I4(n6446), .O(n6447));
  LUT3 #(.INIT(8'hE8)) lut_n6448 (.I0(x1746), .I1(x1747), .I2(x1748), .O(n6448));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6449 (.I0(x1737), .I1(x1738), .I2(x1739), .I3(n6445), .I4(n6446), .O(n6449));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6450 (.I0(x1743), .I1(x1744), .I2(x1745), .I3(n6448), .I4(n6449), .O(n6450));
  LUT3 #(.INIT(8'h96)) lut_n6451 (.I0(n6439), .I1(n6442), .I2(n6443), .O(n6451));
  LUT3 #(.INIT(8'hE8)) lut_n6452 (.I0(n6447), .I1(n6450), .I2(n6451), .O(n6452));
  LUT3 #(.INIT(8'h96)) lut_n6453 (.I0(n6420), .I1(n6428), .I2(n6429), .O(n6453));
  LUT3 #(.INIT(8'hE8)) lut_n6454 (.I0(n6444), .I1(n6452), .I2(n6453), .O(n6454));
  LUT3 #(.INIT(8'hE8)) lut_n6455 (.I0(x1752), .I1(x1753), .I2(x1754), .O(n6455));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6456 (.I0(x1743), .I1(x1744), .I2(x1745), .I3(n6448), .I4(n6449), .O(n6456));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6457 (.I0(x1749), .I1(x1750), .I2(x1751), .I3(n6455), .I4(n6456), .O(n6457));
  LUT3 #(.INIT(8'hE8)) lut_n6458 (.I0(x1758), .I1(x1759), .I2(x1760), .O(n6458));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6459 (.I0(x1749), .I1(x1750), .I2(x1751), .I3(n6455), .I4(n6456), .O(n6459));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6460 (.I0(x1755), .I1(x1756), .I2(x1757), .I3(n6458), .I4(n6459), .O(n6460));
  LUT3 #(.INIT(8'h96)) lut_n6461 (.I0(n6447), .I1(n6450), .I2(n6451), .O(n6461));
  LUT3 #(.INIT(8'hE8)) lut_n6462 (.I0(n6457), .I1(n6460), .I2(n6461), .O(n6462));
  LUT3 #(.INIT(8'hE8)) lut_n6463 (.I0(x1764), .I1(x1765), .I2(x1766), .O(n6463));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6464 (.I0(x1755), .I1(x1756), .I2(x1757), .I3(n6458), .I4(n6459), .O(n6464));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6465 (.I0(x1761), .I1(x1762), .I2(x1763), .I3(n6463), .I4(n6464), .O(n6465));
  LUT3 #(.INIT(8'hE8)) lut_n6466 (.I0(x1770), .I1(x1771), .I2(x1772), .O(n6466));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6467 (.I0(x1761), .I1(x1762), .I2(x1763), .I3(n6463), .I4(n6464), .O(n6467));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6468 (.I0(x1767), .I1(x1768), .I2(x1769), .I3(n6466), .I4(n6467), .O(n6468));
  LUT3 #(.INIT(8'h96)) lut_n6469 (.I0(n6457), .I1(n6460), .I2(n6461), .O(n6469));
  LUT3 #(.INIT(8'hE8)) lut_n6470 (.I0(n6465), .I1(n6468), .I2(n6469), .O(n6470));
  LUT3 #(.INIT(8'h96)) lut_n6471 (.I0(n6444), .I1(n6452), .I2(n6453), .O(n6471));
  LUT3 #(.INIT(8'hE8)) lut_n6472 (.I0(n6462), .I1(n6470), .I2(n6471), .O(n6472));
  LUT3 #(.INIT(8'h96)) lut_n6473 (.I0(n6412), .I1(n6430), .I2(n6431), .O(n6473));
  LUT3 #(.INIT(8'hE8)) lut_n6474 (.I0(n6454), .I1(n6472), .I2(n6473), .O(n6474));
  LUT3 #(.INIT(8'hE8)) lut_n6475 (.I0(x1776), .I1(x1777), .I2(x1778), .O(n6475));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6476 (.I0(x1767), .I1(x1768), .I2(x1769), .I3(n6466), .I4(n6467), .O(n6476));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6477 (.I0(x1773), .I1(x1774), .I2(x1775), .I3(n6475), .I4(n6476), .O(n6477));
  LUT3 #(.INIT(8'hE8)) lut_n6478 (.I0(x1782), .I1(x1783), .I2(x1784), .O(n6478));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6479 (.I0(x1773), .I1(x1774), .I2(x1775), .I3(n6475), .I4(n6476), .O(n6479));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6480 (.I0(x1779), .I1(x1780), .I2(x1781), .I3(n6478), .I4(n6479), .O(n6480));
  LUT3 #(.INIT(8'h96)) lut_n6481 (.I0(n6465), .I1(n6468), .I2(n6469), .O(n6481));
  LUT3 #(.INIT(8'hE8)) lut_n6482 (.I0(n6477), .I1(n6480), .I2(n6481), .O(n6482));
  LUT3 #(.INIT(8'hE8)) lut_n6483 (.I0(x1788), .I1(x1789), .I2(x1790), .O(n6483));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6484 (.I0(x1779), .I1(x1780), .I2(x1781), .I3(n6478), .I4(n6479), .O(n6484));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6485 (.I0(x1785), .I1(x1786), .I2(x1787), .I3(n6483), .I4(n6484), .O(n6485));
  LUT3 #(.INIT(8'hE8)) lut_n6486 (.I0(x1794), .I1(x1795), .I2(x1796), .O(n6486));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6487 (.I0(x1785), .I1(x1786), .I2(x1787), .I3(n6483), .I4(n6484), .O(n6487));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6488 (.I0(x1791), .I1(x1792), .I2(x1793), .I3(n6486), .I4(n6487), .O(n6488));
  LUT3 #(.INIT(8'h96)) lut_n6489 (.I0(n6477), .I1(n6480), .I2(n6481), .O(n6489));
  LUT3 #(.INIT(8'hE8)) lut_n6490 (.I0(n6485), .I1(n6488), .I2(n6489), .O(n6490));
  LUT3 #(.INIT(8'h96)) lut_n6491 (.I0(n6462), .I1(n6470), .I2(n6471), .O(n6491));
  LUT3 #(.INIT(8'hE8)) lut_n6492 (.I0(n6482), .I1(n6490), .I2(n6491), .O(n6492));
  LUT3 #(.INIT(8'hE8)) lut_n6493 (.I0(x1800), .I1(x1801), .I2(x1802), .O(n6493));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6494 (.I0(x1791), .I1(x1792), .I2(x1793), .I3(n6486), .I4(n6487), .O(n6494));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6495 (.I0(x1797), .I1(x1798), .I2(x1799), .I3(n6493), .I4(n6494), .O(n6495));
  LUT3 #(.INIT(8'hE8)) lut_n6496 (.I0(x1806), .I1(x1807), .I2(x1808), .O(n6496));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6497 (.I0(x1797), .I1(x1798), .I2(x1799), .I3(n6493), .I4(n6494), .O(n6497));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6498 (.I0(x1803), .I1(x1804), .I2(x1805), .I3(n6496), .I4(n6497), .O(n6498));
  LUT3 #(.INIT(8'h96)) lut_n6499 (.I0(n6485), .I1(n6488), .I2(n6489), .O(n6499));
  LUT3 #(.INIT(8'hE8)) lut_n6500 (.I0(n6495), .I1(n6498), .I2(n6499), .O(n6500));
  LUT3 #(.INIT(8'hE8)) lut_n6501 (.I0(x1812), .I1(x1813), .I2(x1814), .O(n6501));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6502 (.I0(x1803), .I1(x1804), .I2(x1805), .I3(n6496), .I4(n6497), .O(n6502));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6503 (.I0(x1809), .I1(x1810), .I2(x1811), .I3(n6501), .I4(n6502), .O(n6503));
  LUT3 #(.INIT(8'hE8)) lut_n6504 (.I0(x1818), .I1(x1819), .I2(x1820), .O(n6504));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6505 (.I0(x1809), .I1(x1810), .I2(x1811), .I3(n6501), .I4(n6502), .O(n6505));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6506 (.I0(x1815), .I1(x1816), .I2(x1817), .I3(n6504), .I4(n6505), .O(n6506));
  LUT3 #(.INIT(8'h96)) lut_n6507 (.I0(n6495), .I1(n6498), .I2(n6499), .O(n6507));
  LUT3 #(.INIT(8'hE8)) lut_n6508 (.I0(n6503), .I1(n6506), .I2(n6507), .O(n6508));
  LUT3 #(.INIT(8'h96)) lut_n6509 (.I0(n6482), .I1(n6490), .I2(n6491), .O(n6509));
  LUT3 #(.INIT(8'hE8)) lut_n6510 (.I0(n6500), .I1(n6508), .I2(n6509), .O(n6510));
  LUT3 #(.INIT(8'h96)) lut_n6511 (.I0(n6454), .I1(n6472), .I2(n6473), .O(n6511));
  LUT3 #(.INIT(8'hE8)) lut_n6512 (.I0(n6492), .I1(n6510), .I2(n6511), .O(n6512));
  LUT3 #(.INIT(8'h96)) lut_n6513 (.I0(n6394), .I1(n6432), .I2(n6433), .O(n6513));
  LUT3 #(.INIT(8'hE8)) lut_n6514 (.I0(n6474), .I1(n6512), .I2(n6513), .O(n6514));
  LUT3 #(.INIT(8'hE8)) lut_n6515 (.I0(x1824), .I1(x1825), .I2(x1826), .O(n6515));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6516 (.I0(x1815), .I1(x1816), .I2(x1817), .I3(n6504), .I4(n6505), .O(n6516));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6517 (.I0(x1821), .I1(x1822), .I2(x1823), .I3(n6515), .I4(n6516), .O(n6517));
  LUT3 #(.INIT(8'hE8)) lut_n6518 (.I0(x1830), .I1(x1831), .I2(x1832), .O(n6518));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6519 (.I0(x1821), .I1(x1822), .I2(x1823), .I3(n6515), .I4(n6516), .O(n6519));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6520 (.I0(x1827), .I1(x1828), .I2(x1829), .I3(n6518), .I4(n6519), .O(n6520));
  LUT3 #(.INIT(8'h96)) lut_n6521 (.I0(n6503), .I1(n6506), .I2(n6507), .O(n6521));
  LUT3 #(.INIT(8'hE8)) lut_n6522 (.I0(n6517), .I1(n6520), .I2(n6521), .O(n6522));
  LUT3 #(.INIT(8'hE8)) lut_n6523 (.I0(x1836), .I1(x1837), .I2(x1838), .O(n6523));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6524 (.I0(x1827), .I1(x1828), .I2(x1829), .I3(n6518), .I4(n6519), .O(n6524));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6525 (.I0(x1833), .I1(x1834), .I2(x1835), .I3(n6523), .I4(n6524), .O(n6525));
  LUT3 #(.INIT(8'hE8)) lut_n6526 (.I0(x1842), .I1(x1843), .I2(x1844), .O(n6526));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6527 (.I0(x1833), .I1(x1834), .I2(x1835), .I3(n6523), .I4(n6524), .O(n6527));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6528 (.I0(x1839), .I1(x1840), .I2(x1841), .I3(n6526), .I4(n6527), .O(n6528));
  LUT3 #(.INIT(8'h96)) lut_n6529 (.I0(n6517), .I1(n6520), .I2(n6521), .O(n6529));
  LUT3 #(.INIT(8'hE8)) lut_n6530 (.I0(n6525), .I1(n6528), .I2(n6529), .O(n6530));
  LUT3 #(.INIT(8'h96)) lut_n6531 (.I0(n6500), .I1(n6508), .I2(n6509), .O(n6531));
  LUT3 #(.INIT(8'hE8)) lut_n6532 (.I0(n6522), .I1(n6530), .I2(n6531), .O(n6532));
  LUT3 #(.INIT(8'hE8)) lut_n6533 (.I0(x1848), .I1(x1849), .I2(x1850), .O(n6533));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6534 (.I0(x1839), .I1(x1840), .I2(x1841), .I3(n6526), .I4(n6527), .O(n6534));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6535 (.I0(x1845), .I1(x1846), .I2(x1847), .I3(n6533), .I4(n6534), .O(n6535));
  LUT3 #(.INIT(8'hE8)) lut_n6536 (.I0(x1854), .I1(x1855), .I2(x1856), .O(n6536));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6537 (.I0(x1845), .I1(x1846), .I2(x1847), .I3(n6533), .I4(n6534), .O(n6537));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6538 (.I0(x1851), .I1(x1852), .I2(x1853), .I3(n6536), .I4(n6537), .O(n6538));
  LUT3 #(.INIT(8'h96)) lut_n6539 (.I0(n6525), .I1(n6528), .I2(n6529), .O(n6539));
  LUT3 #(.INIT(8'hE8)) lut_n6540 (.I0(n6535), .I1(n6538), .I2(n6539), .O(n6540));
  LUT3 #(.INIT(8'hE8)) lut_n6541 (.I0(x1860), .I1(x1861), .I2(x1862), .O(n6541));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6542 (.I0(x1851), .I1(x1852), .I2(x1853), .I3(n6536), .I4(n6537), .O(n6542));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6543 (.I0(x1857), .I1(x1858), .I2(x1859), .I3(n6541), .I4(n6542), .O(n6543));
  LUT3 #(.INIT(8'hE8)) lut_n6544 (.I0(x1866), .I1(x1867), .I2(x1868), .O(n6544));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6545 (.I0(x1857), .I1(x1858), .I2(x1859), .I3(n6541), .I4(n6542), .O(n6545));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6546 (.I0(x1863), .I1(x1864), .I2(x1865), .I3(n6544), .I4(n6545), .O(n6546));
  LUT3 #(.INIT(8'h96)) lut_n6547 (.I0(n6535), .I1(n6538), .I2(n6539), .O(n6547));
  LUT3 #(.INIT(8'hE8)) lut_n6548 (.I0(n6543), .I1(n6546), .I2(n6547), .O(n6548));
  LUT3 #(.INIT(8'h96)) lut_n6549 (.I0(n6522), .I1(n6530), .I2(n6531), .O(n6549));
  LUT3 #(.INIT(8'hE8)) lut_n6550 (.I0(n6540), .I1(n6548), .I2(n6549), .O(n6550));
  LUT3 #(.INIT(8'h96)) lut_n6551 (.I0(n6492), .I1(n6510), .I2(n6511), .O(n6551));
  LUT3 #(.INIT(8'hE8)) lut_n6552 (.I0(n6532), .I1(n6550), .I2(n6551), .O(n6552));
  LUT3 #(.INIT(8'hE8)) lut_n6553 (.I0(x1872), .I1(x1873), .I2(x1874), .O(n6553));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6554 (.I0(x1863), .I1(x1864), .I2(x1865), .I3(n6544), .I4(n6545), .O(n6554));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6555 (.I0(x1869), .I1(x1870), .I2(x1871), .I3(n6553), .I4(n6554), .O(n6555));
  LUT3 #(.INIT(8'hE8)) lut_n6556 (.I0(x1878), .I1(x1879), .I2(x1880), .O(n6556));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6557 (.I0(x1869), .I1(x1870), .I2(x1871), .I3(n6553), .I4(n6554), .O(n6557));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6558 (.I0(x1875), .I1(x1876), .I2(x1877), .I3(n6556), .I4(n6557), .O(n6558));
  LUT3 #(.INIT(8'h96)) lut_n6559 (.I0(n6543), .I1(n6546), .I2(n6547), .O(n6559));
  LUT3 #(.INIT(8'hE8)) lut_n6560 (.I0(n6555), .I1(n6558), .I2(n6559), .O(n6560));
  LUT3 #(.INIT(8'hE8)) lut_n6561 (.I0(x1884), .I1(x1885), .I2(x1886), .O(n6561));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6562 (.I0(x1875), .I1(x1876), .I2(x1877), .I3(n6556), .I4(n6557), .O(n6562));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6563 (.I0(x1881), .I1(x1882), .I2(x1883), .I3(n6561), .I4(n6562), .O(n6563));
  LUT3 #(.INIT(8'hE8)) lut_n6564 (.I0(x1890), .I1(x1891), .I2(x1892), .O(n6564));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6565 (.I0(x1881), .I1(x1882), .I2(x1883), .I3(n6561), .I4(n6562), .O(n6565));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6566 (.I0(x1887), .I1(x1888), .I2(x1889), .I3(n6564), .I4(n6565), .O(n6566));
  LUT3 #(.INIT(8'h96)) lut_n6567 (.I0(n6555), .I1(n6558), .I2(n6559), .O(n6567));
  LUT3 #(.INIT(8'hE8)) lut_n6568 (.I0(n6563), .I1(n6566), .I2(n6567), .O(n6568));
  LUT3 #(.INIT(8'h96)) lut_n6569 (.I0(n6540), .I1(n6548), .I2(n6549), .O(n6569));
  LUT3 #(.INIT(8'hE8)) lut_n6570 (.I0(n6560), .I1(n6568), .I2(n6569), .O(n6570));
  LUT3 #(.INIT(8'hE8)) lut_n6571 (.I0(x1896), .I1(x1897), .I2(x1898), .O(n6571));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6572 (.I0(x1887), .I1(x1888), .I2(x1889), .I3(n6564), .I4(n6565), .O(n6572));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6573 (.I0(x1893), .I1(x1894), .I2(x1895), .I3(n6571), .I4(n6572), .O(n6573));
  LUT3 #(.INIT(8'hE8)) lut_n6574 (.I0(x1902), .I1(x1903), .I2(x1904), .O(n6574));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6575 (.I0(x1893), .I1(x1894), .I2(x1895), .I3(n6571), .I4(n6572), .O(n6575));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6576 (.I0(x1899), .I1(x1900), .I2(x1901), .I3(n6574), .I4(n6575), .O(n6576));
  LUT3 #(.INIT(8'h96)) lut_n6577 (.I0(n6563), .I1(n6566), .I2(n6567), .O(n6577));
  LUT3 #(.INIT(8'hE8)) lut_n6578 (.I0(n6573), .I1(n6576), .I2(n6577), .O(n6578));
  LUT3 #(.INIT(8'hE8)) lut_n6579 (.I0(x1908), .I1(x1909), .I2(x1910), .O(n6579));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6580 (.I0(x1899), .I1(x1900), .I2(x1901), .I3(n6574), .I4(n6575), .O(n6580));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6581 (.I0(x1905), .I1(x1906), .I2(x1907), .I3(n6579), .I4(n6580), .O(n6581));
  LUT3 #(.INIT(8'hE8)) lut_n6582 (.I0(x1914), .I1(x1915), .I2(x1916), .O(n6582));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6583 (.I0(x1905), .I1(x1906), .I2(x1907), .I3(n6579), .I4(n6580), .O(n6583));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6584 (.I0(x1911), .I1(x1912), .I2(x1913), .I3(n6582), .I4(n6583), .O(n6584));
  LUT3 #(.INIT(8'h96)) lut_n6585 (.I0(n6573), .I1(n6576), .I2(n6577), .O(n6585));
  LUT3 #(.INIT(8'hE8)) lut_n6586 (.I0(n6581), .I1(n6584), .I2(n6585), .O(n6586));
  LUT3 #(.INIT(8'h96)) lut_n6587 (.I0(n6560), .I1(n6568), .I2(n6569), .O(n6587));
  LUT3 #(.INIT(8'hE8)) lut_n6588 (.I0(n6578), .I1(n6586), .I2(n6587), .O(n6588));
  LUT3 #(.INIT(8'h96)) lut_n6589 (.I0(n6532), .I1(n6550), .I2(n6551), .O(n6589));
  LUT3 #(.INIT(8'hE8)) lut_n6590 (.I0(n6570), .I1(n6588), .I2(n6589), .O(n6590));
  LUT3 #(.INIT(8'h96)) lut_n6591 (.I0(n6474), .I1(n6512), .I2(n6513), .O(n6591));
  LUT3 #(.INIT(8'hE8)) lut_n6592 (.I0(n6552), .I1(n6590), .I2(n6591), .O(n6592));
  LUT3 #(.INIT(8'h96)) lut_n6593 (.I0(n6356), .I1(n6434), .I2(n6435), .O(n6593));
  LUT3 #(.INIT(8'hE8)) lut_n6594 (.I0(n6514), .I1(n6592), .I2(n6593), .O(n6594));
  LUT3 #(.INIT(8'h96)) lut_n6595 (.I0(n6117), .I1(n6275), .I2(n6276), .O(n6595));
  LUT3 #(.INIT(8'hE8)) lut_n6596 (.I0(n6436), .I1(n6594), .I2(n6595), .O(n6596));
  LUT3 #(.INIT(8'hE8)) lut_n6597 (.I0(x1920), .I1(x1921), .I2(x1922), .O(n6597));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6598 (.I0(x1911), .I1(x1912), .I2(x1913), .I3(n6582), .I4(n6583), .O(n6598));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6599 (.I0(x1917), .I1(x1918), .I2(x1919), .I3(n6597), .I4(n6598), .O(n6599));
  LUT3 #(.INIT(8'hE8)) lut_n6600 (.I0(x1926), .I1(x1927), .I2(x1928), .O(n6600));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6601 (.I0(x1917), .I1(x1918), .I2(x1919), .I3(n6597), .I4(n6598), .O(n6601));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6602 (.I0(x1923), .I1(x1924), .I2(x1925), .I3(n6600), .I4(n6601), .O(n6602));
  LUT3 #(.INIT(8'h96)) lut_n6603 (.I0(n6581), .I1(n6584), .I2(n6585), .O(n6603));
  LUT3 #(.INIT(8'hE8)) lut_n6604 (.I0(n6599), .I1(n6602), .I2(n6603), .O(n6604));
  LUT3 #(.INIT(8'hE8)) lut_n6605 (.I0(x1932), .I1(x1933), .I2(x1934), .O(n6605));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6606 (.I0(x1923), .I1(x1924), .I2(x1925), .I3(n6600), .I4(n6601), .O(n6606));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6607 (.I0(x1929), .I1(x1930), .I2(x1931), .I3(n6605), .I4(n6606), .O(n6607));
  LUT3 #(.INIT(8'hE8)) lut_n6608 (.I0(x1938), .I1(x1939), .I2(x1940), .O(n6608));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6609 (.I0(x1929), .I1(x1930), .I2(x1931), .I3(n6605), .I4(n6606), .O(n6609));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6610 (.I0(x1935), .I1(x1936), .I2(x1937), .I3(n6608), .I4(n6609), .O(n6610));
  LUT3 #(.INIT(8'h96)) lut_n6611 (.I0(n6599), .I1(n6602), .I2(n6603), .O(n6611));
  LUT3 #(.INIT(8'hE8)) lut_n6612 (.I0(n6607), .I1(n6610), .I2(n6611), .O(n6612));
  LUT3 #(.INIT(8'h96)) lut_n6613 (.I0(n6578), .I1(n6586), .I2(n6587), .O(n6613));
  LUT3 #(.INIT(8'hE8)) lut_n6614 (.I0(n6604), .I1(n6612), .I2(n6613), .O(n6614));
  LUT3 #(.INIT(8'hE8)) lut_n6615 (.I0(x1944), .I1(x1945), .I2(x1946), .O(n6615));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6616 (.I0(x1935), .I1(x1936), .I2(x1937), .I3(n6608), .I4(n6609), .O(n6616));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6617 (.I0(x1941), .I1(x1942), .I2(x1943), .I3(n6615), .I4(n6616), .O(n6617));
  LUT3 #(.INIT(8'hE8)) lut_n6618 (.I0(x1950), .I1(x1951), .I2(x1952), .O(n6618));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6619 (.I0(x1941), .I1(x1942), .I2(x1943), .I3(n6615), .I4(n6616), .O(n6619));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6620 (.I0(x1947), .I1(x1948), .I2(x1949), .I3(n6618), .I4(n6619), .O(n6620));
  LUT3 #(.INIT(8'h96)) lut_n6621 (.I0(n6607), .I1(n6610), .I2(n6611), .O(n6621));
  LUT3 #(.INIT(8'hE8)) lut_n6622 (.I0(n6617), .I1(n6620), .I2(n6621), .O(n6622));
  LUT3 #(.INIT(8'hE8)) lut_n6623 (.I0(x1956), .I1(x1957), .I2(x1958), .O(n6623));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6624 (.I0(x1947), .I1(x1948), .I2(x1949), .I3(n6618), .I4(n6619), .O(n6624));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6625 (.I0(x1953), .I1(x1954), .I2(x1955), .I3(n6623), .I4(n6624), .O(n6625));
  LUT3 #(.INIT(8'hE8)) lut_n6626 (.I0(x1962), .I1(x1963), .I2(x1964), .O(n6626));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6627 (.I0(x1953), .I1(x1954), .I2(x1955), .I3(n6623), .I4(n6624), .O(n6627));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6628 (.I0(x1959), .I1(x1960), .I2(x1961), .I3(n6626), .I4(n6627), .O(n6628));
  LUT3 #(.INIT(8'h96)) lut_n6629 (.I0(n6617), .I1(n6620), .I2(n6621), .O(n6629));
  LUT3 #(.INIT(8'hE8)) lut_n6630 (.I0(n6625), .I1(n6628), .I2(n6629), .O(n6630));
  LUT3 #(.INIT(8'h96)) lut_n6631 (.I0(n6604), .I1(n6612), .I2(n6613), .O(n6631));
  LUT3 #(.INIT(8'hE8)) lut_n6632 (.I0(n6622), .I1(n6630), .I2(n6631), .O(n6632));
  LUT3 #(.INIT(8'h96)) lut_n6633 (.I0(n6570), .I1(n6588), .I2(n6589), .O(n6633));
  LUT3 #(.INIT(8'hE8)) lut_n6634 (.I0(n6614), .I1(n6632), .I2(n6633), .O(n6634));
  LUT3 #(.INIT(8'hE8)) lut_n6635 (.I0(x1968), .I1(x1969), .I2(x1970), .O(n6635));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6636 (.I0(x1959), .I1(x1960), .I2(x1961), .I3(n6626), .I4(n6627), .O(n6636));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6637 (.I0(x1965), .I1(x1966), .I2(x1967), .I3(n6635), .I4(n6636), .O(n6637));
  LUT3 #(.INIT(8'hE8)) lut_n6638 (.I0(x1974), .I1(x1975), .I2(x1976), .O(n6638));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6639 (.I0(x1965), .I1(x1966), .I2(x1967), .I3(n6635), .I4(n6636), .O(n6639));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6640 (.I0(x1971), .I1(x1972), .I2(x1973), .I3(n6638), .I4(n6639), .O(n6640));
  LUT3 #(.INIT(8'h96)) lut_n6641 (.I0(n6625), .I1(n6628), .I2(n6629), .O(n6641));
  LUT3 #(.INIT(8'hE8)) lut_n6642 (.I0(n6637), .I1(n6640), .I2(n6641), .O(n6642));
  LUT3 #(.INIT(8'hE8)) lut_n6643 (.I0(x1980), .I1(x1981), .I2(x1982), .O(n6643));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6644 (.I0(x1971), .I1(x1972), .I2(x1973), .I3(n6638), .I4(n6639), .O(n6644));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6645 (.I0(x1977), .I1(x1978), .I2(x1979), .I3(n6643), .I4(n6644), .O(n6645));
  LUT3 #(.INIT(8'hE8)) lut_n6646 (.I0(x1986), .I1(x1987), .I2(x1988), .O(n6646));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6647 (.I0(x1977), .I1(x1978), .I2(x1979), .I3(n6643), .I4(n6644), .O(n6647));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6648 (.I0(x1983), .I1(x1984), .I2(x1985), .I3(n6646), .I4(n6647), .O(n6648));
  LUT3 #(.INIT(8'h96)) lut_n6649 (.I0(n6637), .I1(n6640), .I2(n6641), .O(n6649));
  LUT3 #(.INIT(8'hE8)) lut_n6650 (.I0(n6645), .I1(n6648), .I2(n6649), .O(n6650));
  LUT3 #(.INIT(8'h96)) lut_n6651 (.I0(n6622), .I1(n6630), .I2(n6631), .O(n6651));
  LUT3 #(.INIT(8'hE8)) lut_n6652 (.I0(n6642), .I1(n6650), .I2(n6651), .O(n6652));
  LUT3 #(.INIT(8'hE8)) lut_n6653 (.I0(x1992), .I1(x1993), .I2(x1994), .O(n6653));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6654 (.I0(x1983), .I1(x1984), .I2(x1985), .I3(n6646), .I4(n6647), .O(n6654));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6655 (.I0(x1989), .I1(x1990), .I2(x1991), .I3(n6653), .I4(n6654), .O(n6655));
  LUT3 #(.INIT(8'hE8)) lut_n6656 (.I0(x1998), .I1(x1999), .I2(x2000), .O(n6656));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6657 (.I0(x1989), .I1(x1990), .I2(x1991), .I3(n6653), .I4(n6654), .O(n6657));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6658 (.I0(x1995), .I1(x1996), .I2(x1997), .I3(n6656), .I4(n6657), .O(n6658));
  LUT3 #(.INIT(8'h96)) lut_n6659 (.I0(n6645), .I1(n6648), .I2(n6649), .O(n6659));
  LUT3 #(.INIT(8'hE8)) lut_n6660 (.I0(n6655), .I1(n6658), .I2(n6659), .O(n6660));
  LUT3 #(.INIT(8'hE8)) lut_n6661 (.I0(x2004), .I1(x2005), .I2(x2006), .O(n6661));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6662 (.I0(x1995), .I1(x1996), .I2(x1997), .I3(n6656), .I4(n6657), .O(n6662));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6663 (.I0(x2001), .I1(x2002), .I2(x2003), .I3(n6661), .I4(n6662), .O(n6663));
  LUT3 #(.INIT(8'hE8)) lut_n6664 (.I0(x2010), .I1(x2011), .I2(x2012), .O(n6664));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6665 (.I0(x2001), .I1(x2002), .I2(x2003), .I3(n6661), .I4(n6662), .O(n6665));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6666 (.I0(x2007), .I1(x2008), .I2(x2009), .I3(n6664), .I4(n6665), .O(n6666));
  LUT3 #(.INIT(8'h96)) lut_n6667 (.I0(n6655), .I1(n6658), .I2(n6659), .O(n6667));
  LUT3 #(.INIT(8'hE8)) lut_n6668 (.I0(n6663), .I1(n6666), .I2(n6667), .O(n6668));
  LUT3 #(.INIT(8'h96)) lut_n6669 (.I0(n6642), .I1(n6650), .I2(n6651), .O(n6669));
  LUT3 #(.INIT(8'hE8)) lut_n6670 (.I0(n6660), .I1(n6668), .I2(n6669), .O(n6670));
  LUT3 #(.INIT(8'h96)) lut_n6671 (.I0(n6614), .I1(n6632), .I2(n6633), .O(n6671));
  LUT3 #(.INIT(8'hE8)) lut_n6672 (.I0(n6652), .I1(n6670), .I2(n6671), .O(n6672));
  LUT3 #(.INIT(8'h96)) lut_n6673 (.I0(n6552), .I1(n6590), .I2(n6591), .O(n6673));
  LUT3 #(.INIT(8'hE8)) lut_n6674 (.I0(n6634), .I1(n6672), .I2(n6673), .O(n6674));
  LUT3 #(.INIT(8'hE8)) lut_n6675 (.I0(x2016), .I1(x2017), .I2(x2018), .O(n6675));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6676 (.I0(x2007), .I1(x2008), .I2(x2009), .I3(n6664), .I4(n6665), .O(n6676));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6677 (.I0(x2013), .I1(x2014), .I2(x2015), .I3(n6675), .I4(n6676), .O(n6677));
  LUT3 #(.INIT(8'hE8)) lut_n6678 (.I0(x2022), .I1(x2023), .I2(x2024), .O(n6678));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6679 (.I0(x2013), .I1(x2014), .I2(x2015), .I3(n6675), .I4(n6676), .O(n6679));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6680 (.I0(x2019), .I1(x2020), .I2(x2021), .I3(n6678), .I4(n6679), .O(n6680));
  LUT3 #(.INIT(8'h96)) lut_n6681 (.I0(n6663), .I1(n6666), .I2(n6667), .O(n6681));
  LUT3 #(.INIT(8'hE8)) lut_n6682 (.I0(n6677), .I1(n6680), .I2(n6681), .O(n6682));
  LUT3 #(.INIT(8'hE8)) lut_n6683 (.I0(x2028), .I1(x2029), .I2(x2030), .O(n6683));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6684 (.I0(x2019), .I1(x2020), .I2(x2021), .I3(n6678), .I4(n6679), .O(n6684));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6685 (.I0(x2025), .I1(x2026), .I2(x2027), .I3(n6683), .I4(n6684), .O(n6685));
  LUT3 #(.INIT(8'hE8)) lut_n6686 (.I0(x2034), .I1(x2035), .I2(x2036), .O(n6686));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6687 (.I0(x2025), .I1(x2026), .I2(x2027), .I3(n6683), .I4(n6684), .O(n6687));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6688 (.I0(x2031), .I1(x2032), .I2(x2033), .I3(n6686), .I4(n6687), .O(n6688));
  LUT3 #(.INIT(8'h96)) lut_n6689 (.I0(n6677), .I1(n6680), .I2(n6681), .O(n6689));
  LUT3 #(.INIT(8'hE8)) lut_n6690 (.I0(n6685), .I1(n6688), .I2(n6689), .O(n6690));
  LUT3 #(.INIT(8'h96)) lut_n6691 (.I0(n6660), .I1(n6668), .I2(n6669), .O(n6691));
  LUT3 #(.INIT(8'hE8)) lut_n6692 (.I0(n6682), .I1(n6690), .I2(n6691), .O(n6692));
  LUT3 #(.INIT(8'hE8)) lut_n6693 (.I0(x2040), .I1(x2041), .I2(x2042), .O(n6693));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6694 (.I0(x2031), .I1(x2032), .I2(x2033), .I3(n6686), .I4(n6687), .O(n6694));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6695 (.I0(x2037), .I1(x2038), .I2(x2039), .I3(n6693), .I4(n6694), .O(n6695));
  LUT3 #(.INIT(8'hE8)) lut_n6696 (.I0(x2046), .I1(x2047), .I2(x2048), .O(n6696));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6697 (.I0(x2037), .I1(x2038), .I2(x2039), .I3(n6693), .I4(n6694), .O(n6697));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6698 (.I0(x2043), .I1(x2044), .I2(x2045), .I3(n6696), .I4(n6697), .O(n6698));
  LUT3 #(.INIT(8'h96)) lut_n6699 (.I0(n6685), .I1(n6688), .I2(n6689), .O(n6699));
  LUT3 #(.INIT(8'hE8)) lut_n6700 (.I0(n6695), .I1(n6698), .I2(n6699), .O(n6700));
  LUT3 #(.INIT(8'hE8)) lut_n6701 (.I0(x2052), .I1(x2053), .I2(x2054), .O(n6701));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6702 (.I0(x2043), .I1(x2044), .I2(x2045), .I3(n6696), .I4(n6697), .O(n6702));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6703 (.I0(x2049), .I1(x2050), .I2(x2051), .I3(n6701), .I4(n6702), .O(n6703));
  LUT3 #(.INIT(8'hE8)) lut_n6704 (.I0(x2058), .I1(x2059), .I2(x2060), .O(n6704));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6705 (.I0(x2049), .I1(x2050), .I2(x2051), .I3(n6701), .I4(n6702), .O(n6705));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6706 (.I0(x2055), .I1(x2056), .I2(x2057), .I3(n6704), .I4(n6705), .O(n6706));
  LUT3 #(.INIT(8'h96)) lut_n6707 (.I0(n6695), .I1(n6698), .I2(n6699), .O(n6707));
  LUT3 #(.INIT(8'hE8)) lut_n6708 (.I0(n6703), .I1(n6706), .I2(n6707), .O(n6708));
  LUT3 #(.INIT(8'h96)) lut_n6709 (.I0(n6682), .I1(n6690), .I2(n6691), .O(n6709));
  LUT3 #(.INIT(8'hE8)) lut_n6710 (.I0(n6700), .I1(n6708), .I2(n6709), .O(n6710));
  LUT3 #(.INIT(8'h96)) lut_n6711 (.I0(n6652), .I1(n6670), .I2(n6671), .O(n6711));
  LUT3 #(.INIT(8'hE8)) lut_n6712 (.I0(n6692), .I1(n6710), .I2(n6711), .O(n6712));
  LUT3 #(.INIT(8'hE8)) lut_n6713 (.I0(x2064), .I1(x2065), .I2(x2066), .O(n6713));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6714 (.I0(x2055), .I1(x2056), .I2(x2057), .I3(n6704), .I4(n6705), .O(n6714));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6715 (.I0(x2061), .I1(x2062), .I2(x2063), .I3(n6713), .I4(n6714), .O(n6715));
  LUT3 #(.INIT(8'hE8)) lut_n6716 (.I0(x2070), .I1(x2071), .I2(x2072), .O(n6716));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6717 (.I0(x2061), .I1(x2062), .I2(x2063), .I3(n6713), .I4(n6714), .O(n6717));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6718 (.I0(x2067), .I1(x2068), .I2(x2069), .I3(n6716), .I4(n6717), .O(n6718));
  LUT3 #(.INIT(8'h96)) lut_n6719 (.I0(n6703), .I1(n6706), .I2(n6707), .O(n6719));
  LUT3 #(.INIT(8'hE8)) lut_n6720 (.I0(n6715), .I1(n6718), .I2(n6719), .O(n6720));
  LUT3 #(.INIT(8'hE8)) lut_n6721 (.I0(x2076), .I1(x2077), .I2(x2078), .O(n6721));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6722 (.I0(x2067), .I1(x2068), .I2(x2069), .I3(n6716), .I4(n6717), .O(n6722));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6723 (.I0(x2073), .I1(x2074), .I2(x2075), .I3(n6721), .I4(n6722), .O(n6723));
  LUT3 #(.INIT(8'hE8)) lut_n6724 (.I0(x2082), .I1(x2083), .I2(x2084), .O(n6724));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6725 (.I0(x2073), .I1(x2074), .I2(x2075), .I3(n6721), .I4(n6722), .O(n6725));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6726 (.I0(x2079), .I1(x2080), .I2(x2081), .I3(n6724), .I4(n6725), .O(n6726));
  LUT3 #(.INIT(8'h96)) lut_n6727 (.I0(n6715), .I1(n6718), .I2(n6719), .O(n6727));
  LUT3 #(.INIT(8'hE8)) lut_n6728 (.I0(n6723), .I1(n6726), .I2(n6727), .O(n6728));
  LUT3 #(.INIT(8'h96)) lut_n6729 (.I0(n6700), .I1(n6708), .I2(n6709), .O(n6729));
  LUT3 #(.INIT(8'hE8)) lut_n6730 (.I0(n6720), .I1(n6728), .I2(n6729), .O(n6730));
  LUT3 #(.INIT(8'hE8)) lut_n6731 (.I0(x2088), .I1(x2089), .I2(x2090), .O(n6731));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6732 (.I0(x2079), .I1(x2080), .I2(x2081), .I3(n6724), .I4(n6725), .O(n6732));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6733 (.I0(x2085), .I1(x2086), .I2(x2087), .I3(n6731), .I4(n6732), .O(n6733));
  LUT3 #(.INIT(8'hE8)) lut_n6734 (.I0(x2094), .I1(x2095), .I2(x2096), .O(n6734));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6735 (.I0(x2085), .I1(x2086), .I2(x2087), .I3(n6731), .I4(n6732), .O(n6735));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6736 (.I0(x2091), .I1(x2092), .I2(x2093), .I3(n6734), .I4(n6735), .O(n6736));
  LUT3 #(.INIT(8'h96)) lut_n6737 (.I0(n6723), .I1(n6726), .I2(n6727), .O(n6737));
  LUT3 #(.INIT(8'hE8)) lut_n6738 (.I0(n6733), .I1(n6736), .I2(n6737), .O(n6738));
  LUT3 #(.INIT(8'hE8)) lut_n6739 (.I0(x2100), .I1(x2101), .I2(x2102), .O(n6739));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6740 (.I0(x2091), .I1(x2092), .I2(x2093), .I3(n6734), .I4(n6735), .O(n6740));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6741 (.I0(x2097), .I1(x2098), .I2(x2099), .I3(n6739), .I4(n6740), .O(n6741));
  LUT3 #(.INIT(8'hE8)) lut_n6742 (.I0(x2106), .I1(x2107), .I2(x2108), .O(n6742));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6743 (.I0(x2097), .I1(x2098), .I2(x2099), .I3(n6739), .I4(n6740), .O(n6743));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6744 (.I0(x2103), .I1(x2104), .I2(x2105), .I3(n6742), .I4(n6743), .O(n6744));
  LUT3 #(.INIT(8'h96)) lut_n6745 (.I0(n6733), .I1(n6736), .I2(n6737), .O(n6745));
  LUT3 #(.INIT(8'hE8)) lut_n6746 (.I0(n6741), .I1(n6744), .I2(n6745), .O(n6746));
  LUT3 #(.INIT(8'h96)) lut_n6747 (.I0(n6720), .I1(n6728), .I2(n6729), .O(n6747));
  LUT3 #(.INIT(8'hE8)) lut_n6748 (.I0(n6738), .I1(n6746), .I2(n6747), .O(n6748));
  LUT3 #(.INIT(8'h96)) lut_n6749 (.I0(n6692), .I1(n6710), .I2(n6711), .O(n6749));
  LUT3 #(.INIT(8'hE8)) lut_n6750 (.I0(n6730), .I1(n6748), .I2(n6749), .O(n6750));
  LUT3 #(.INIT(8'h96)) lut_n6751 (.I0(n6634), .I1(n6672), .I2(n6673), .O(n6751));
  LUT3 #(.INIT(8'hE8)) lut_n6752 (.I0(n6712), .I1(n6750), .I2(n6751), .O(n6752));
  LUT3 #(.INIT(8'h96)) lut_n6753 (.I0(n6514), .I1(n6592), .I2(n6593), .O(n6753));
  LUT3 #(.INIT(8'hE8)) lut_n6754 (.I0(n6674), .I1(n6752), .I2(n6753), .O(n6754));
  LUT3 #(.INIT(8'hE8)) lut_n6755 (.I0(x2112), .I1(x2113), .I2(x2114), .O(n6755));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6756 (.I0(x2103), .I1(x2104), .I2(x2105), .I3(n6742), .I4(n6743), .O(n6756));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6757 (.I0(x2109), .I1(x2110), .I2(x2111), .I3(n6755), .I4(n6756), .O(n6757));
  LUT3 #(.INIT(8'hE8)) lut_n6758 (.I0(x2118), .I1(x2119), .I2(x2120), .O(n6758));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6759 (.I0(x2109), .I1(x2110), .I2(x2111), .I3(n6755), .I4(n6756), .O(n6759));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6760 (.I0(x2115), .I1(x2116), .I2(x2117), .I3(n6758), .I4(n6759), .O(n6760));
  LUT3 #(.INIT(8'h96)) lut_n6761 (.I0(n6741), .I1(n6744), .I2(n6745), .O(n6761));
  LUT3 #(.INIT(8'hE8)) lut_n6762 (.I0(n6757), .I1(n6760), .I2(n6761), .O(n6762));
  LUT3 #(.INIT(8'hE8)) lut_n6763 (.I0(x2124), .I1(x2125), .I2(x2126), .O(n6763));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6764 (.I0(x2115), .I1(x2116), .I2(x2117), .I3(n6758), .I4(n6759), .O(n6764));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6765 (.I0(x2121), .I1(x2122), .I2(x2123), .I3(n6763), .I4(n6764), .O(n6765));
  LUT3 #(.INIT(8'hE8)) lut_n6766 (.I0(x2130), .I1(x2131), .I2(x2132), .O(n6766));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6767 (.I0(x2121), .I1(x2122), .I2(x2123), .I3(n6763), .I4(n6764), .O(n6767));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6768 (.I0(x2127), .I1(x2128), .I2(x2129), .I3(n6766), .I4(n6767), .O(n6768));
  LUT3 #(.INIT(8'h96)) lut_n6769 (.I0(n6757), .I1(n6760), .I2(n6761), .O(n6769));
  LUT3 #(.INIT(8'hE8)) lut_n6770 (.I0(n6765), .I1(n6768), .I2(n6769), .O(n6770));
  LUT3 #(.INIT(8'h96)) lut_n6771 (.I0(n6738), .I1(n6746), .I2(n6747), .O(n6771));
  LUT3 #(.INIT(8'hE8)) lut_n6772 (.I0(n6762), .I1(n6770), .I2(n6771), .O(n6772));
  LUT3 #(.INIT(8'hE8)) lut_n6773 (.I0(x2136), .I1(x2137), .I2(x2138), .O(n6773));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6774 (.I0(x2127), .I1(x2128), .I2(x2129), .I3(n6766), .I4(n6767), .O(n6774));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6775 (.I0(x2133), .I1(x2134), .I2(x2135), .I3(n6773), .I4(n6774), .O(n6775));
  LUT3 #(.INIT(8'hE8)) lut_n6776 (.I0(x2142), .I1(x2143), .I2(x2144), .O(n6776));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6777 (.I0(x2133), .I1(x2134), .I2(x2135), .I3(n6773), .I4(n6774), .O(n6777));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6778 (.I0(x2139), .I1(x2140), .I2(x2141), .I3(n6776), .I4(n6777), .O(n6778));
  LUT3 #(.INIT(8'h96)) lut_n6779 (.I0(n6765), .I1(n6768), .I2(n6769), .O(n6779));
  LUT3 #(.INIT(8'hE8)) lut_n6780 (.I0(n6775), .I1(n6778), .I2(n6779), .O(n6780));
  LUT3 #(.INIT(8'hE8)) lut_n6781 (.I0(x2148), .I1(x2149), .I2(x2150), .O(n6781));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6782 (.I0(x2139), .I1(x2140), .I2(x2141), .I3(n6776), .I4(n6777), .O(n6782));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6783 (.I0(x2145), .I1(x2146), .I2(x2147), .I3(n6781), .I4(n6782), .O(n6783));
  LUT3 #(.INIT(8'hE8)) lut_n6784 (.I0(x2154), .I1(x2155), .I2(x2156), .O(n6784));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6785 (.I0(x2145), .I1(x2146), .I2(x2147), .I3(n6781), .I4(n6782), .O(n6785));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6786 (.I0(x2151), .I1(x2152), .I2(x2153), .I3(n6784), .I4(n6785), .O(n6786));
  LUT3 #(.INIT(8'h96)) lut_n6787 (.I0(n6775), .I1(n6778), .I2(n6779), .O(n6787));
  LUT3 #(.INIT(8'hE8)) lut_n6788 (.I0(n6783), .I1(n6786), .I2(n6787), .O(n6788));
  LUT3 #(.INIT(8'h96)) lut_n6789 (.I0(n6762), .I1(n6770), .I2(n6771), .O(n6789));
  LUT3 #(.INIT(8'hE8)) lut_n6790 (.I0(n6780), .I1(n6788), .I2(n6789), .O(n6790));
  LUT3 #(.INIT(8'h96)) lut_n6791 (.I0(n6730), .I1(n6748), .I2(n6749), .O(n6791));
  LUT3 #(.INIT(8'hE8)) lut_n6792 (.I0(n6772), .I1(n6790), .I2(n6791), .O(n6792));
  LUT3 #(.INIT(8'hE8)) lut_n6793 (.I0(x2160), .I1(x2161), .I2(x2162), .O(n6793));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6794 (.I0(x2151), .I1(x2152), .I2(x2153), .I3(n6784), .I4(n6785), .O(n6794));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6795 (.I0(x2157), .I1(x2158), .I2(x2159), .I3(n6793), .I4(n6794), .O(n6795));
  LUT3 #(.INIT(8'hE8)) lut_n6796 (.I0(x2166), .I1(x2167), .I2(x2168), .O(n6796));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6797 (.I0(x2157), .I1(x2158), .I2(x2159), .I3(n6793), .I4(n6794), .O(n6797));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6798 (.I0(x2163), .I1(x2164), .I2(x2165), .I3(n6796), .I4(n6797), .O(n6798));
  LUT3 #(.INIT(8'h96)) lut_n6799 (.I0(n6783), .I1(n6786), .I2(n6787), .O(n6799));
  LUT3 #(.INIT(8'hE8)) lut_n6800 (.I0(n6795), .I1(n6798), .I2(n6799), .O(n6800));
  LUT3 #(.INIT(8'hE8)) lut_n6801 (.I0(x2172), .I1(x2173), .I2(x2174), .O(n6801));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6802 (.I0(x2163), .I1(x2164), .I2(x2165), .I3(n6796), .I4(n6797), .O(n6802));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6803 (.I0(x2169), .I1(x2170), .I2(x2171), .I3(n6801), .I4(n6802), .O(n6803));
  LUT3 #(.INIT(8'hE8)) lut_n6804 (.I0(x2178), .I1(x2179), .I2(x2180), .O(n6804));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6805 (.I0(x2169), .I1(x2170), .I2(x2171), .I3(n6801), .I4(n6802), .O(n6805));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6806 (.I0(x2175), .I1(x2176), .I2(x2177), .I3(n6804), .I4(n6805), .O(n6806));
  LUT3 #(.INIT(8'h96)) lut_n6807 (.I0(n6795), .I1(n6798), .I2(n6799), .O(n6807));
  LUT3 #(.INIT(8'hE8)) lut_n6808 (.I0(n6803), .I1(n6806), .I2(n6807), .O(n6808));
  LUT3 #(.INIT(8'h96)) lut_n6809 (.I0(n6780), .I1(n6788), .I2(n6789), .O(n6809));
  LUT3 #(.INIT(8'hE8)) lut_n6810 (.I0(n6800), .I1(n6808), .I2(n6809), .O(n6810));
  LUT3 #(.INIT(8'hE8)) lut_n6811 (.I0(x2184), .I1(x2185), .I2(x2186), .O(n6811));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6812 (.I0(x2175), .I1(x2176), .I2(x2177), .I3(n6804), .I4(n6805), .O(n6812));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6813 (.I0(x2181), .I1(x2182), .I2(x2183), .I3(n6811), .I4(n6812), .O(n6813));
  LUT3 #(.INIT(8'hE8)) lut_n6814 (.I0(x2190), .I1(x2191), .I2(x2192), .O(n6814));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6815 (.I0(x2181), .I1(x2182), .I2(x2183), .I3(n6811), .I4(n6812), .O(n6815));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6816 (.I0(x2187), .I1(x2188), .I2(x2189), .I3(n6814), .I4(n6815), .O(n6816));
  LUT3 #(.INIT(8'h96)) lut_n6817 (.I0(n6803), .I1(n6806), .I2(n6807), .O(n6817));
  LUT3 #(.INIT(8'hE8)) lut_n6818 (.I0(n6813), .I1(n6816), .I2(n6817), .O(n6818));
  LUT3 #(.INIT(8'hE8)) lut_n6819 (.I0(x2196), .I1(x2197), .I2(x2198), .O(n6819));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6820 (.I0(x2187), .I1(x2188), .I2(x2189), .I3(n6814), .I4(n6815), .O(n6820));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6821 (.I0(x2193), .I1(x2194), .I2(x2195), .I3(n6819), .I4(n6820), .O(n6821));
  LUT3 #(.INIT(8'hE8)) lut_n6822 (.I0(x2202), .I1(x2203), .I2(x2204), .O(n6822));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6823 (.I0(x2193), .I1(x2194), .I2(x2195), .I3(n6819), .I4(n6820), .O(n6823));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6824 (.I0(x2199), .I1(x2200), .I2(x2201), .I3(n6822), .I4(n6823), .O(n6824));
  LUT3 #(.INIT(8'h96)) lut_n6825 (.I0(n6813), .I1(n6816), .I2(n6817), .O(n6825));
  LUT3 #(.INIT(8'hE8)) lut_n6826 (.I0(n6821), .I1(n6824), .I2(n6825), .O(n6826));
  LUT3 #(.INIT(8'h96)) lut_n6827 (.I0(n6800), .I1(n6808), .I2(n6809), .O(n6827));
  LUT3 #(.INIT(8'hE8)) lut_n6828 (.I0(n6818), .I1(n6826), .I2(n6827), .O(n6828));
  LUT3 #(.INIT(8'h96)) lut_n6829 (.I0(n6772), .I1(n6790), .I2(n6791), .O(n6829));
  LUT3 #(.INIT(8'hE8)) lut_n6830 (.I0(n6810), .I1(n6828), .I2(n6829), .O(n6830));
  LUT3 #(.INIT(8'h96)) lut_n6831 (.I0(n6712), .I1(n6750), .I2(n6751), .O(n6831));
  LUT3 #(.INIT(8'hE8)) lut_n6832 (.I0(n6792), .I1(n6830), .I2(n6831), .O(n6832));
  LUT3 #(.INIT(8'hE8)) lut_n6833 (.I0(x2208), .I1(x2209), .I2(x2210), .O(n6833));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6834 (.I0(x2199), .I1(x2200), .I2(x2201), .I3(n6822), .I4(n6823), .O(n6834));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6835 (.I0(x2205), .I1(x2206), .I2(x2207), .I3(n6833), .I4(n6834), .O(n6835));
  LUT3 #(.INIT(8'hE8)) lut_n6836 (.I0(x2214), .I1(x2215), .I2(x2216), .O(n6836));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6837 (.I0(x2205), .I1(x2206), .I2(x2207), .I3(n6833), .I4(n6834), .O(n6837));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6838 (.I0(x2211), .I1(x2212), .I2(x2213), .I3(n6836), .I4(n6837), .O(n6838));
  LUT3 #(.INIT(8'h96)) lut_n6839 (.I0(n6821), .I1(n6824), .I2(n6825), .O(n6839));
  LUT3 #(.INIT(8'hE8)) lut_n6840 (.I0(n6835), .I1(n6838), .I2(n6839), .O(n6840));
  LUT3 #(.INIT(8'hE8)) lut_n6841 (.I0(x2220), .I1(x2221), .I2(x2222), .O(n6841));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6842 (.I0(x2211), .I1(x2212), .I2(x2213), .I3(n6836), .I4(n6837), .O(n6842));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6843 (.I0(x2217), .I1(x2218), .I2(x2219), .I3(n6841), .I4(n6842), .O(n6843));
  LUT3 #(.INIT(8'hE8)) lut_n6844 (.I0(x2226), .I1(x2227), .I2(x2228), .O(n6844));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6845 (.I0(x2217), .I1(x2218), .I2(x2219), .I3(n6841), .I4(n6842), .O(n6845));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6846 (.I0(x2223), .I1(x2224), .I2(x2225), .I3(n6844), .I4(n6845), .O(n6846));
  LUT3 #(.INIT(8'h96)) lut_n6847 (.I0(n6835), .I1(n6838), .I2(n6839), .O(n6847));
  LUT3 #(.INIT(8'hE8)) lut_n6848 (.I0(n6843), .I1(n6846), .I2(n6847), .O(n6848));
  LUT3 #(.INIT(8'h96)) lut_n6849 (.I0(n6818), .I1(n6826), .I2(n6827), .O(n6849));
  LUT3 #(.INIT(8'hE8)) lut_n6850 (.I0(n6840), .I1(n6848), .I2(n6849), .O(n6850));
  LUT3 #(.INIT(8'hE8)) lut_n6851 (.I0(x2232), .I1(x2233), .I2(x2234), .O(n6851));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6852 (.I0(x2223), .I1(x2224), .I2(x2225), .I3(n6844), .I4(n6845), .O(n6852));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6853 (.I0(x2229), .I1(x2230), .I2(x2231), .I3(n6851), .I4(n6852), .O(n6853));
  LUT3 #(.INIT(8'hE8)) lut_n6854 (.I0(x2238), .I1(x2239), .I2(x2240), .O(n6854));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6855 (.I0(x2229), .I1(x2230), .I2(x2231), .I3(n6851), .I4(n6852), .O(n6855));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6856 (.I0(x2235), .I1(x2236), .I2(x2237), .I3(n6854), .I4(n6855), .O(n6856));
  LUT3 #(.INIT(8'h96)) lut_n6857 (.I0(n6843), .I1(n6846), .I2(n6847), .O(n6857));
  LUT3 #(.INIT(8'hE8)) lut_n6858 (.I0(n6853), .I1(n6856), .I2(n6857), .O(n6858));
  LUT3 #(.INIT(8'hE8)) lut_n6859 (.I0(x2244), .I1(x2245), .I2(x2246), .O(n6859));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6860 (.I0(x2235), .I1(x2236), .I2(x2237), .I3(n6854), .I4(n6855), .O(n6860));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6861 (.I0(x2241), .I1(x2242), .I2(x2243), .I3(n6859), .I4(n6860), .O(n6861));
  LUT3 #(.INIT(8'hE8)) lut_n6862 (.I0(x2250), .I1(x2251), .I2(x2252), .O(n6862));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6863 (.I0(x2241), .I1(x2242), .I2(x2243), .I3(n6859), .I4(n6860), .O(n6863));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6864 (.I0(x2247), .I1(x2248), .I2(x2249), .I3(n6862), .I4(n6863), .O(n6864));
  LUT3 #(.INIT(8'h96)) lut_n6865 (.I0(n6853), .I1(n6856), .I2(n6857), .O(n6865));
  LUT3 #(.INIT(8'hE8)) lut_n6866 (.I0(n6861), .I1(n6864), .I2(n6865), .O(n6866));
  LUT3 #(.INIT(8'h96)) lut_n6867 (.I0(n6840), .I1(n6848), .I2(n6849), .O(n6867));
  LUT3 #(.INIT(8'hE8)) lut_n6868 (.I0(n6858), .I1(n6866), .I2(n6867), .O(n6868));
  LUT3 #(.INIT(8'h96)) lut_n6869 (.I0(n6810), .I1(n6828), .I2(n6829), .O(n6869));
  LUT3 #(.INIT(8'hE8)) lut_n6870 (.I0(n6850), .I1(n6868), .I2(n6869), .O(n6870));
  LUT3 #(.INIT(8'hE8)) lut_n6871 (.I0(x2256), .I1(x2257), .I2(x2258), .O(n6871));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6872 (.I0(x2247), .I1(x2248), .I2(x2249), .I3(n6862), .I4(n6863), .O(n6872));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6873 (.I0(x2253), .I1(x2254), .I2(x2255), .I3(n6871), .I4(n6872), .O(n6873));
  LUT3 #(.INIT(8'hE8)) lut_n6874 (.I0(x2262), .I1(x2263), .I2(x2264), .O(n6874));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6875 (.I0(x2253), .I1(x2254), .I2(x2255), .I3(n6871), .I4(n6872), .O(n6875));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6876 (.I0(x2259), .I1(x2260), .I2(x2261), .I3(n6874), .I4(n6875), .O(n6876));
  LUT3 #(.INIT(8'h96)) lut_n6877 (.I0(n6861), .I1(n6864), .I2(n6865), .O(n6877));
  LUT3 #(.INIT(8'hE8)) lut_n6878 (.I0(n6873), .I1(n6876), .I2(n6877), .O(n6878));
  LUT3 #(.INIT(8'hE8)) lut_n6879 (.I0(x2268), .I1(x2269), .I2(x2270), .O(n6879));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6880 (.I0(x2259), .I1(x2260), .I2(x2261), .I3(n6874), .I4(n6875), .O(n6880));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6881 (.I0(x2265), .I1(x2266), .I2(x2267), .I3(n6879), .I4(n6880), .O(n6881));
  LUT3 #(.INIT(8'hE8)) lut_n6882 (.I0(x2274), .I1(x2275), .I2(x2276), .O(n6882));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6883 (.I0(x2265), .I1(x2266), .I2(x2267), .I3(n6879), .I4(n6880), .O(n6883));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6884 (.I0(x2271), .I1(x2272), .I2(x2273), .I3(n6882), .I4(n6883), .O(n6884));
  LUT3 #(.INIT(8'h96)) lut_n6885 (.I0(n6873), .I1(n6876), .I2(n6877), .O(n6885));
  LUT3 #(.INIT(8'hE8)) lut_n6886 (.I0(n6881), .I1(n6884), .I2(n6885), .O(n6886));
  LUT3 #(.INIT(8'h96)) lut_n6887 (.I0(n6858), .I1(n6866), .I2(n6867), .O(n6887));
  LUT3 #(.INIT(8'hE8)) lut_n6888 (.I0(n6878), .I1(n6886), .I2(n6887), .O(n6888));
  LUT3 #(.INIT(8'hE8)) lut_n6889 (.I0(x2280), .I1(x2281), .I2(x2282), .O(n6889));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6890 (.I0(x2271), .I1(x2272), .I2(x2273), .I3(n6882), .I4(n6883), .O(n6890));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6891 (.I0(x2277), .I1(x2278), .I2(x2279), .I3(n6889), .I4(n6890), .O(n6891));
  LUT3 #(.INIT(8'hE8)) lut_n6892 (.I0(x2286), .I1(x2287), .I2(x2288), .O(n6892));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6893 (.I0(x2277), .I1(x2278), .I2(x2279), .I3(n6889), .I4(n6890), .O(n6893));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6894 (.I0(x2283), .I1(x2284), .I2(x2285), .I3(n6892), .I4(n6893), .O(n6894));
  LUT3 #(.INIT(8'h96)) lut_n6895 (.I0(n6881), .I1(n6884), .I2(n6885), .O(n6895));
  LUT3 #(.INIT(8'hE8)) lut_n6896 (.I0(n6891), .I1(n6894), .I2(n6895), .O(n6896));
  LUT3 #(.INIT(8'hE8)) lut_n6897 (.I0(x2292), .I1(x2293), .I2(x2294), .O(n6897));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6898 (.I0(x2283), .I1(x2284), .I2(x2285), .I3(n6892), .I4(n6893), .O(n6898));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6899 (.I0(x2289), .I1(x2290), .I2(x2291), .I3(n6897), .I4(n6898), .O(n6899));
  LUT3 #(.INIT(8'hE8)) lut_n6900 (.I0(x2298), .I1(x2299), .I2(x2300), .O(n6900));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6901 (.I0(x2289), .I1(x2290), .I2(x2291), .I3(n6897), .I4(n6898), .O(n6901));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6902 (.I0(x2295), .I1(x2296), .I2(x2297), .I3(n6900), .I4(n6901), .O(n6902));
  LUT3 #(.INIT(8'h96)) lut_n6903 (.I0(n6891), .I1(n6894), .I2(n6895), .O(n6903));
  LUT3 #(.INIT(8'hE8)) lut_n6904 (.I0(n6899), .I1(n6902), .I2(n6903), .O(n6904));
  LUT3 #(.INIT(8'h96)) lut_n6905 (.I0(n6878), .I1(n6886), .I2(n6887), .O(n6905));
  LUT3 #(.INIT(8'hE8)) lut_n6906 (.I0(n6896), .I1(n6904), .I2(n6905), .O(n6906));
  LUT3 #(.INIT(8'h96)) lut_n6907 (.I0(n6850), .I1(n6868), .I2(n6869), .O(n6907));
  LUT3 #(.INIT(8'hE8)) lut_n6908 (.I0(n6888), .I1(n6906), .I2(n6907), .O(n6908));
  LUT3 #(.INIT(8'h96)) lut_n6909 (.I0(n6792), .I1(n6830), .I2(n6831), .O(n6909));
  LUT3 #(.INIT(8'hE8)) lut_n6910 (.I0(n6870), .I1(n6908), .I2(n6909), .O(n6910));
  LUT3 #(.INIT(8'h96)) lut_n6911 (.I0(n6674), .I1(n6752), .I2(n6753), .O(n6911));
  LUT3 #(.INIT(8'hE8)) lut_n6912 (.I0(n6832), .I1(n6910), .I2(n6911), .O(n6912));
  LUT3 #(.INIT(8'h96)) lut_n6913 (.I0(n6436), .I1(n6594), .I2(n6595), .O(n6913));
  LUT3 #(.INIT(8'hE8)) lut_n6914 (.I0(n6754), .I1(n6912), .I2(n6913), .O(n6914));
  LUT3 #(.INIT(8'h96)) lut_n6915 (.I0(n5641), .I1(n5959), .I2(n6277), .O(n6915));
  LUT3 #(.INIT(8'hE8)) lut_n6916 (.I0(n6596), .I1(n6914), .I2(n6915), .O(n6916));
  LUT3 #(.INIT(8'hE8)) lut_n6917 (.I0(x2304), .I1(x2305), .I2(x2306), .O(n6917));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6918 (.I0(x2295), .I1(x2296), .I2(x2297), .I3(n6900), .I4(n6901), .O(n6918));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6919 (.I0(x2301), .I1(x2302), .I2(x2303), .I3(n6917), .I4(n6918), .O(n6919));
  LUT3 #(.INIT(8'hE8)) lut_n6920 (.I0(x2310), .I1(x2311), .I2(x2312), .O(n6920));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6921 (.I0(x2301), .I1(x2302), .I2(x2303), .I3(n6917), .I4(n6918), .O(n6921));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6922 (.I0(x2307), .I1(x2308), .I2(x2309), .I3(n6920), .I4(n6921), .O(n6922));
  LUT3 #(.INIT(8'h96)) lut_n6923 (.I0(n6899), .I1(n6902), .I2(n6903), .O(n6923));
  LUT3 #(.INIT(8'hE8)) lut_n6924 (.I0(n6919), .I1(n6922), .I2(n6923), .O(n6924));
  LUT3 #(.INIT(8'hE8)) lut_n6925 (.I0(x2316), .I1(x2317), .I2(x2318), .O(n6925));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6926 (.I0(x2307), .I1(x2308), .I2(x2309), .I3(n6920), .I4(n6921), .O(n6926));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6927 (.I0(x2313), .I1(x2314), .I2(x2315), .I3(n6925), .I4(n6926), .O(n6927));
  LUT3 #(.INIT(8'hE8)) lut_n6928 (.I0(x2322), .I1(x2323), .I2(x2324), .O(n6928));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6929 (.I0(x2313), .I1(x2314), .I2(x2315), .I3(n6925), .I4(n6926), .O(n6929));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6930 (.I0(x2319), .I1(x2320), .I2(x2321), .I3(n6928), .I4(n6929), .O(n6930));
  LUT3 #(.INIT(8'h96)) lut_n6931 (.I0(n6919), .I1(n6922), .I2(n6923), .O(n6931));
  LUT3 #(.INIT(8'hE8)) lut_n6932 (.I0(n6927), .I1(n6930), .I2(n6931), .O(n6932));
  LUT3 #(.INIT(8'h96)) lut_n6933 (.I0(n6896), .I1(n6904), .I2(n6905), .O(n6933));
  LUT3 #(.INIT(8'hE8)) lut_n6934 (.I0(n6924), .I1(n6932), .I2(n6933), .O(n6934));
  LUT3 #(.INIT(8'hE8)) lut_n6935 (.I0(x2328), .I1(x2329), .I2(x2330), .O(n6935));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6936 (.I0(x2319), .I1(x2320), .I2(x2321), .I3(n6928), .I4(n6929), .O(n6936));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6937 (.I0(x2325), .I1(x2326), .I2(x2327), .I3(n6935), .I4(n6936), .O(n6937));
  LUT3 #(.INIT(8'hE8)) lut_n6938 (.I0(x2334), .I1(x2335), .I2(x2336), .O(n6938));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6939 (.I0(x2325), .I1(x2326), .I2(x2327), .I3(n6935), .I4(n6936), .O(n6939));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6940 (.I0(x2331), .I1(x2332), .I2(x2333), .I3(n6938), .I4(n6939), .O(n6940));
  LUT3 #(.INIT(8'h96)) lut_n6941 (.I0(n6927), .I1(n6930), .I2(n6931), .O(n6941));
  LUT3 #(.INIT(8'hE8)) lut_n6942 (.I0(n6937), .I1(n6940), .I2(n6941), .O(n6942));
  LUT3 #(.INIT(8'hE8)) lut_n6943 (.I0(x2340), .I1(x2341), .I2(x2342), .O(n6943));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6944 (.I0(x2331), .I1(x2332), .I2(x2333), .I3(n6938), .I4(n6939), .O(n6944));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6945 (.I0(x2337), .I1(x2338), .I2(x2339), .I3(n6943), .I4(n6944), .O(n6945));
  LUT3 #(.INIT(8'hE8)) lut_n6946 (.I0(x2346), .I1(x2347), .I2(x2348), .O(n6946));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6947 (.I0(x2337), .I1(x2338), .I2(x2339), .I3(n6943), .I4(n6944), .O(n6947));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6948 (.I0(x2343), .I1(x2344), .I2(x2345), .I3(n6946), .I4(n6947), .O(n6948));
  LUT3 #(.INIT(8'h96)) lut_n6949 (.I0(n6937), .I1(n6940), .I2(n6941), .O(n6949));
  LUT3 #(.INIT(8'hE8)) lut_n6950 (.I0(n6945), .I1(n6948), .I2(n6949), .O(n6950));
  LUT3 #(.INIT(8'h96)) lut_n6951 (.I0(n6924), .I1(n6932), .I2(n6933), .O(n6951));
  LUT3 #(.INIT(8'hE8)) lut_n6952 (.I0(n6942), .I1(n6950), .I2(n6951), .O(n6952));
  LUT3 #(.INIT(8'h96)) lut_n6953 (.I0(n6888), .I1(n6906), .I2(n6907), .O(n6953));
  LUT3 #(.INIT(8'hE8)) lut_n6954 (.I0(n6934), .I1(n6952), .I2(n6953), .O(n6954));
  LUT3 #(.INIT(8'hE8)) lut_n6955 (.I0(x2352), .I1(x2353), .I2(x2354), .O(n6955));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6956 (.I0(x2343), .I1(x2344), .I2(x2345), .I3(n6946), .I4(n6947), .O(n6956));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6957 (.I0(x2349), .I1(x2350), .I2(x2351), .I3(n6955), .I4(n6956), .O(n6957));
  LUT3 #(.INIT(8'hE8)) lut_n6958 (.I0(x2358), .I1(x2359), .I2(x2360), .O(n6958));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6959 (.I0(x2349), .I1(x2350), .I2(x2351), .I3(n6955), .I4(n6956), .O(n6959));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6960 (.I0(x2355), .I1(x2356), .I2(x2357), .I3(n6958), .I4(n6959), .O(n6960));
  LUT3 #(.INIT(8'h96)) lut_n6961 (.I0(n6945), .I1(n6948), .I2(n6949), .O(n6961));
  LUT3 #(.INIT(8'hE8)) lut_n6962 (.I0(n6957), .I1(n6960), .I2(n6961), .O(n6962));
  LUT3 #(.INIT(8'hE8)) lut_n6963 (.I0(x2364), .I1(x2365), .I2(x2366), .O(n6963));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6964 (.I0(x2355), .I1(x2356), .I2(x2357), .I3(n6958), .I4(n6959), .O(n6964));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6965 (.I0(x2361), .I1(x2362), .I2(x2363), .I3(n6963), .I4(n6964), .O(n6965));
  LUT3 #(.INIT(8'hE8)) lut_n6966 (.I0(x2370), .I1(x2371), .I2(x2372), .O(n6966));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6967 (.I0(x2361), .I1(x2362), .I2(x2363), .I3(n6963), .I4(n6964), .O(n6967));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6968 (.I0(x2367), .I1(x2368), .I2(x2369), .I3(n6966), .I4(n6967), .O(n6968));
  LUT3 #(.INIT(8'h96)) lut_n6969 (.I0(n6957), .I1(n6960), .I2(n6961), .O(n6969));
  LUT3 #(.INIT(8'hE8)) lut_n6970 (.I0(n6965), .I1(n6968), .I2(n6969), .O(n6970));
  LUT3 #(.INIT(8'h96)) lut_n6971 (.I0(n6942), .I1(n6950), .I2(n6951), .O(n6971));
  LUT3 #(.INIT(8'hE8)) lut_n6972 (.I0(n6962), .I1(n6970), .I2(n6971), .O(n6972));
  LUT3 #(.INIT(8'hE8)) lut_n6973 (.I0(x2376), .I1(x2377), .I2(x2378), .O(n6973));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6974 (.I0(x2367), .I1(x2368), .I2(x2369), .I3(n6966), .I4(n6967), .O(n6974));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6975 (.I0(x2373), .I1(x2374), .I2(x2375), .I3(n6973), .I4(n6974), .O(n6975));
  LUT3 #(.INIT(8'hE8)) lut_n6976 (.I0(x2382), .I1(x2383), .I2(x2384), .O(n6976));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6977 (.I0(x2373), .I1(x2374), .I2(x2375), .I3(n6973), .I4(n6974), .O(n6977));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6978 (.I0(x2379), .I1(x2380), .I2(x2381), .I3(n6976), .I4(n6977), .O(n6978));
  LUT3 #(.INIT(8'h96)) lut_n6979 (.I0(n6965), .I1(n6968), .I2(n6969), .O(n6979));
  LUT3 #(.INIT(8'hE8)) lut_n6980 (.I0(n6975), .I1(n6978), .I2(n6979), .O(n6980));
  LUT3 #(.INIT(8'hE8)) lut_n6981 (.I0(x2388), .I1(x2389), .I2(x2390), .O(n6981));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6982 (.I0(x2379), .I1(x2380), .I2(x2381), .I3(n6976), .I4(n6977), .O(n6982));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6983 (.I0(x2385), .I1(x2386), .I2(x2387), .I3(n6981), .I4(n6982), .O(n6983));
  LUT3 #(.INIT(8'hE8)) lut_n6984 (.I0(x2394), .I1(x2395), .I2(x2396), .O(n6984));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6985 (.I0(x2385), .I1(x2386), .I2(x2387), .I3(n6981), .I4(n6982), .O(n6985));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6986 (.I0(x2391), .I1(x2392), .I2(x2393), .I3(n6984), .I4(n6985), .O(n6986));
  LUT3 #(.INIT(8'h96)) lut_n6987 (.I0(n6975), .I1(n6978), .I2(n6979), .O(n6987));
  LUT3 #(.INIT(8'hE8)) lut_n6988 (.I0(n6983), .I1(n6986), .I2(n6987), .O(n6988));
  LUT3 #(.INIT(8'h96)) lut_n6989 (.I0(n6962), .I1(n6970), .I2(n6971), .O(n6989));
  LUT3 #(.INIT(8'hE8)) lut_n6990 (.I0(n6980), .I1(n6988), .I2(n6989), .O(n6990));
  LUT3 #(.INIT(8'h96)) lut_n6991 (.I0(n6934), .I1(n6952), .I2(n6953), .O(n6991));
  LUT3 #(.INIT(8'hE8)) lut_n6992 (.I0(n6972), .I1(n6990), .I2(n6991), .O(n6992));
  LUT3 #(.INIT(8'h96)) lut_n6993 (.I0(n6870), .I1(n6908), .I2(n6909), .O(n6993));
  LUT3 #(.INIT(8'hE8)) lut_n6994 (.I0(n6954), .I1(n6992), .I2(n6993), .O(n6994));
  LUT3 #(.INIT(8'hE8)) lut_n6995 (.I0(x2400), .I1(x2401), .I2(x2402), .O(n6995));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6996 (.I0(x2391), .I1(x2392), .I2(x2393), .I3(n6984), .I4(n6985), .O(n6996));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n6997 (.I0(x2397), .I1(x2398), .I2(x2399), .I3(n6995), .I4(n6996), .O(n6997));
  LUT3 #(.INIT(8'hE8)) lut_n6998 (.I0(x2406), .I1(x2407), .I2(x2408), .O(n6998));
  LUT5 #(.INIT(32'hE81717E8)) lut_n6999 (.I0(x2397), .I1(x2398), .I2(x2399), .I3(n6995), .I4(n6996), .O(n6999));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7000 (.I0(x2403), .I1(x2404), .I2(x2405), .I3(n6998), .I4(n6999), .O(n7000));
  LUT3 #(.INIT(8'h96)) lut_n7001 (.I0(n6983), .I1(n6986), .I2(n6987), .O(n7001));
  LUT3 #(.INIT(8'hE8)) lut_n7002 (.I0(n6997), .I1(n7000), .I2(n7001), .O(n7002));
  LUT3 #(.INIT(8'hE8)) lut_n7003 (.I0(x2412), .I1(x2413), .I2(x2414), .O(n7003));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7004 (.I0(x2403), .I1(x2404), .I2(x2405), .I3(n6998), .I4(n6999), .O(n7004));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7005 (.I0(x2409), .I1(x2410), .I2(x2411), .I3(n7003), .I4(n7004), .O(n7005));
  LUT3 #(.INIT(8'hE8)) lut_n7006 (.I0(x2418), .I1(x2419), .I2(x2420), .O(n7006));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7007 (.I0(x2409), .I1(x2410), .I2(x2411), .I3(n7003), .I4(n7004), .O(n7007));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7008 (.I0(x2415), .I1(x2416), .I2(x2417), .I3(n7006), .I4(n7007), .O(n7008));
  LUT3 #(.INIT(8'h96)) lut_n7009 (.I0(n6997), .I1(n7000), .I2(n7001), .O(n7009));
  LUT3 #(.INIT(8'hE8)) lut_n7010 (.I0(n7005), .I1(n7008), .I2(n7009), .O(n7010));
  LUT3 #(.INIT(8'h96)) lut_n7011 (.I0(n6980), .I1(n6988), .I2(n6989), .O(n7011));
  LUT3 #(.INIT(8'hE8)) lut_n7012 (.I0(n7002), .I1(n7010), .I2(n7011), .O(n7012));
  LUT3 #(.INIT(8'hE8)) lut_n7013 (.I0(x2424), .I1(x2425), .I2(x2426), .O(n7013));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7014 (.I0(x2415), .I1(x2416), .I2(x2417), .I3(n7006), .I4(n7007), .O(n7014));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7015 (.I0(x2421), .I1(x2422), .I2(x2423), .I3(n7013), .I4(n7014), .O(n7015));
  LUT3 #(.INIT(8'hE8)) lut_n7016 (.I0(x2430), .I1(x2431), .I2(x2432), .O(n7016));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7017 (.I0(x2421), .I1(x2422), .I2(x2423), .I3(n7013), .I4(n7014), .O(n7017));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7018 (.I0(x2427), .I1(x2428), .I2(x2429), .I3(n7016), .I4(n7017), .O(n7018));
  LUT3 #(.INIT(8'h96)) lut_n7019 (.I0(n7005), .I1(n7008), .I2(n7009), .O(n7019));
  LUT3 #(.INIT(8'hE8)) lut_n7020 (.I0(n7015), .I1(n7018), .I2(n7019), .O(n7020));
  LUT3 #(.INIT(8'hE8)) lut_n7021 (.I0(x2436), .I1(x2437), .I2(x2438), .O(n7021));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7022 (.I0(x2427), .I1(x2428), .I2(x2429), .I3(n7016), .I4(n7017), .O(n7022));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7023 (.I0(x2433), .I1(x2434), .I2(x2435), .I3(n7021), .I4(n7022), .O(n7023));
  LUT3 #(.INIT(8'hE8)) lut_n7024 (.I0(x2442), .I1(x2443), .I2(x2444), .O(n7024));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7025 (.I0(x2433), .I1(x2434), .I2(x2435), .I3(n7021), .I4(n7022), .O(n7025));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7026 (.I0(x2439), .I1(x2440), .I2(x2441), .I3(n7024), .I4(n7025), .O(n7026));
  LUT3 #(.INIT(8'h96)) lut_n7027 (.I0(n7015), .I1(n7018), .I2(n7019), .O(n7027));
  LUT3 #(.INIT(8'hE8)) lut_n7028 (.I0(n7023), .I1(n7026), .I2(n7027), .O(n7028));
  LUT3 #(.INIT(8'h96)) lut_n7029 (.I0(n7002), .I1(n7010), .I2(n7011), .O(n7029));
  LUT3 #(.INIT(8'hE8)) lut_n7030 (.I0(n7020), .I1(n7028), .I2(n7029), .O(n7030));
  LUT3 #(.INIT(8'h96)) lut_n7031 (.I0(n6972), .I1(n6990), .I2(n6991), .O(n7031));
  LUT3 #(.INIT(8'hE8)) lut_n7032 (.I0(n7012), .I1(n7030), .I2(n7031), .O(n7032));
  LUT3 #(.INIT(8'hE8)) lut_n7033 (.I0(x2448), .I1(x2449), .I2(x2450), .O(n7033));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7034 (.I0(x2439), .I1(x2440), .I2(x2441), .I3(n7024), .I4(n7025), .O(n7034));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7035 (.I0(x2445), .I1(x2446), .I2(x2447), .I3(n7033), .I4(n7034), .O(n7035));
  LUT3 #(.INIT(8'hE8)) lut_n7036 (.I0(x2454), .I1(x2455), .I2(x2456), .O(n7036));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7037 (.I0(x2445), .I1(x2446), .I2(x2447), .I3(n7033), .I4(n7034), .O(n7037));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7038 (.I0(x2451), .I1(x2452), .I2(x2453), .I3(n7036), .I4(n7037), .O(n7038));
  LUT3 #(.INIT(8'h96)) lut_n7039 (.I0(n7023), .I1(n7026), .I2(n7027), .O(n7039));
  LUT3 #(.INIT(8'hE8)) lut_n7040 (.I0(n7035), .I1(n7038), .I2(n7039), .O(n7040));
  LUT3 #(.INIT(8'hE8)) lut_n7041 (.I0(x2460), .I1(x2461), .I2(x2462), .O(n7041));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7042 (.I0(x2451), .I1(x2452), .I2(x2453), .I3(n7036), .I4(n7037), .O(n7042));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7043 (.I0(x2457), .I1(x2458), .I2(x2459), .I3(n7041), .I4(n7042), .O(n7043));
  LUT3 #(.INIT(8'hE8)) lut_n7044 (.I0(x2466), .I1(x2467), .I2(x2468), .O(n7044));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7045 (.I0(x2457), .I1(x2458), .I2(x2459), .I3(n7041), .I4(n7042), .O(n7045));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7046 (.I0(x2463), .I1(x2464), .I2(x2465), .I3(n7044), .I4(n7045), .O(n7046));
  LUT3 #(.INIT(8'h96)) lut_n7047 (.I0(n7035), .I1(n7038), .I2(n7039), .O(n7047));
  LUT3 #(.INIT(8'hE8)) lut_n7048 (.I0(n7043), .I1(n7046), .I2(n7047), .O(n7048));
  LUT3 #(.INIT(8'h96)) lut_n7049 (.I0(n7020), .I1(n7028), .I2(n7029), .O(n7049));
  LUT3 #(.INIT(8'hE8)) lut_n7050 (.I0(n7040), .I1(n7048), .I2(n7049), .O(n7050));
  LUT3 #(.INIT(8'hE8)) lut_n7051 (.I0(x2472), .I1(x2473), .I2(x2474), .O(n7051));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7052 (.I0(x2463), .I1(x2464), .I2(x2465), .I3(n7044), .I4(n7045), .O(n7052));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7053 (.I0(x2469), .I1(x2470), .I2(x2471), .I3(n7051), .I4(n7052), .O(n7053));
  LUT3 #(.INIT(8'hE8)) lut_n7054 (.I0(x2478), .I1(x2479), .I2(x2480), .O(n7054));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7055 (.I0(x2469), .I1(x2470), .I2(x2471), .I3(n7051), .I4(n7052), .O(n7055));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7056 (.I0(x2475), .I1(x2476), .I2(x2477), .I3(n7054), .I4(n7055), .O(n7056));
  LUT3 #(.INIT(8'h96)) lut_n7057 (.I0(n7043), .I1(n7046), .I2(n7047), .O(n7057));
  LUT3 #(.INIT(8'hE8)) lut_n7058 (.I0(n7053), .I1(n7056), .I2(n7057), .O(n7058));
  LUT3 #(.INIT(8'hE8)) lut_n7059 (.I0(x2484), .I1(x2485), .I2(x2486), .O(n7059));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7060 (.I0(x2475), .I1(x2476), .I2(x2477), .I3(n7054), .I4(n7055), .O(n7060));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7061 (.I0(x2481), .I1(x2482), .I2(x2483), .I3(n7059), .I4(n7060), .O(n7061));
  LUT3 #(.INIT(8'hE8)) lut_n7062 (.I0(x2490), .I1(x2491), .I2(x2492), .O(n7062));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7063 (.I0(x2481), .I1(x2482), .I2(x2483), .I3(n7059), .I4(n7060), .O(n7063));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7064 (.I0(x2487), .I1(x2488), .I2(x2489), .I3(n7062), .I4(n7063), .O(n7064));
  LUT3 #(.INIT(8'h96)) lut_n7065 (.I0(n7053), .I1(n7056), .I2(n7057), .O(n7065));
  LUT3 #(.INIT(8'hE8)) lut_n7066 (.I0(n7061), .I1(n7064), .I2(n7065), .O(n7066));
  LUT3 #(.INIT(8'h96)) lut_n7067 (.I0(n7040), .I1(n7048), .I2(n7049), .O(n7067));
  LUT3 #(.INIT(8'hE8)) lut_n7068 (.I0(n7058), .I1(n7066), .I2(n7067), .O(n7068));
  LUT3 #(.INIT(8'h96)) lut_n7069 (.I0(n7012), .I1(n7030), .I2(n7031), .O(n7069));
  LUT3 #(.INIT(8'hE8)) lut_n7070 (.I0(n7050), .I1(n7068), .I2(n7069), .O(n7070));
  LUT3 #(.INIT(8'h96)) lut_n7071 (.I0(n6954), .I1(n6992), .I2(n6993), .O(n7071));
  LUT3 #(.INIT(8'hE8)) lut_n7072 (.I0(n7032), .I1(n7070), .I2(n7071), .O(n7072));
  LUT3 #(.INIT(8'h96)) lut_n7073 (.I0(n6832), .I1(n6910), .I2(n6911), .O(n7073));
  LUT3 #(.INIT(8'hE8)) lut_n7074 (.I0(n6994), .I1(n7072), .I2(n7073), .O(n7074));
  LUT3 #(.INIT(8'hE8)) lut_n7075 (.I0(x2496), .I1(x2497), .I2(x2498), .O(n7075));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7076 (.I0(x2487), .I1(x2488), .I2(x2489), .I3(n7062), .I4(n7063), .O(n7076));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7077 (.I0(x2493), .I1(x2494), .I2(x2495), .I3(n7075), .I4(n7076), .O(n7077));
  LUT3 #(.INIT(8'hE8)) lut_n7078 (.I0(x2502), .I1(x2503), .I2(x2504), .O(n7078));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7079 (.I0(x2493), .I1(x2494), .I2(x2495), .I3(n7075), .I4(n7076), .O(n7079));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7080 (.I0(x2499), .I1(x2500), .I2(x2501), .I3(n7078), .I4(n7079), .O(n7080));
  LUT3 #(.INIT(8'h96)) lut_n7081 (.I0(n7061), .I1(n7064), .I2(n7065), .O(n7081));
  LUT3 #(.INIT(8'hE8)) lut_n7082 (.I0(n7077), .I1(n7080), .I2(n7081), .O(n7082));
  LUT3 #(.INIT(8'hE8)) lut_n7083 (.I0(x2508), .I1(x2509), .I2(x2510), .O(n7083));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7084 (.I0(x2499), .I1(x2500), .I2(x2501), .I3(n7078), .I4(n7079), .O(n7084));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7085 (.I0(x2505), .I1(x2506), .I2(x2507), .I3(n7083), .I4(n7084), .O(n7085));
  LUT3 #(.INIT(8'hE8)) lut_n7086 (.I0(x2514), .I1(x2515), .I2(x2516), .O(n7086));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7087 (.I0(x2505), .I1(x2506), .I2(x2507), .I3(n7083), .I4(n7084), .O(n7087));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7088 (.I0(x2511), .I1(x2512), .I2(x2513), .I3(n7086), .I4(n7087), .O(n7088));
  LUT3 #(.INIT(8'h96)) lut_n7089 (.I0(n7077), .I1(n7080), .I2(n7081), .O(n7089));
  LUT3 #(.INIT(8'hE8)) lut_n7090 (.I0(n7085), .I1(n7088), .I2(n7089), .O(n7090));
  LUT3 #(.INIT(8'h96)) lut_n7091 (.I0(n7058), .I1(n7066), .I2(n7067), .O(n7091));
  LUT3 #(.INIT(8'hE8)) lut_n7092 (.I0(n7082), .I1(n7090), .I2(n7091), .O(n7092));
  LUT3 #(.INIT(8'hE8)) lut_n7093 (.I0(x2520), .I1(x2521), .I2(x2522), .O(n7093));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7094 (.I0(x2511), .I1(x2512), .I2(x2513), .I3(n7086), .I4(n7087), .O(n7094));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7095 (.I0(x2517), .I1(x2518), .I2(x2519), .I3(n7093), .I4(n7094), .O(n7095));
  LUT3 #(.INIT(8'hE8)) lut_n7096 (.I0(x2526), .I1(x2527), .I2(x2528), .O(n7096));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7097 (.I0(x2517), .I1(x2518), .I2(x2519), .I3(n7093), .I4(n7094), .O(n7097));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7098 (.I0(x2523), .I1(x2524), .I2(x2525), .I3(n7096), .I4(n7097), .O(n7098));
  LUT3 #(.INIT(8'h96)) lut_n7099 (.I0(n7085), .I1(n7088), .I2(n7089), .O(n7099));
  LUT3 #(.INIT(8'hE8)) lut_n7100 (.I0(n7095), .I1(n7098), .I2(n7099), .O(n7100));
  LUT3 #(.INIT(8'hE8)) lut_n7101 (.I0(x2532), .I1(x2533), .I2(x2534), .O(n7101));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7102 (.I0(x2523), .I1(x2524), .I2(x2525), .I3(n7096), .I4(n7097), .O(n7102));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7103 (.I0(x2529), .I1(x2530), .I2(x2531), .I3(n7101), .I4(n7102), .O(n7103));
  LUT3 #(.INIT(8'hE8)) lut_n7104 (.I0(x2538), .I1(x2539), .I2(x2540), .O(n7104));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7105 (.I0(x2529), .I1(x2530), .I2(x2531), .I3(n7101), .I4(n7102), .O(n7105));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7106 (.I0(x2535), .I1(x2536), .I2(x2537), .I3(n7104), .I4(n7105), .O(n7106));
  LUT3 #(.INIT(8'h96)) lut_n7107 (.I0(n7095), .I1(n7098), .I2(n7099), .O(n7107));
  LUT3 #(.INIT(8'hE8)) lut_n7108 (.I0(n7103), .I1(n7106), .I2(n7107), .O(n7108));
  LUT3 #(.INIT(8'h96)) lut_n7109 (.I0(n7082), .I1(n7090), .I2(n7091), .O(n7109));
  LUT3 #(.INIT(8'hE8)) lut_n7110 (.I0(n7100), .I1(n7108), .I2(n7109), .O(n7110));
  LUT3 #(.INIT(8'h96)) lut_n7111 (.I0(n7050), .I1(n7068), .I2(n7069), .O(n7111));
  LUT3 #(.INIT(8'hE8)) lut_n7112 (.I0(n7092), .I1(n7110), .I2(n7111), .O(n7112));
  LUT3 #(.INIT(8'hE8)) lut_n7113 (.I0(x2544), .I1(x2545), .I2(x2546), .O(n7113));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7114 (.I0(x2535), .I1(x2536), .I2(x2537), .I3(n7104), .I4(n7105), .O(n7114));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7115 (.I0(x2541), .I1(x2542), .I2(x2543), .I3(n7113), .I4(n7114), .O(n7115));
  LUT3 #(.INIT(8'hE8)) lut_n7116 (.I0(x2550), .I1(x2551), .I2(x2552), .O(n7116));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7117 (.I0(x2541), .I1(x2542), .I2(x2543), .I3(n7113), .I4(n7114), .O(n7117));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7118 (.I0(x2547), .I1(x2548), .I2(x2549), .I3(n7116), .I4(n7117), .O(n7118));
  LUT3 #(.INIT(8'h96)) lut_n7119 (.I0(n7103), .I1(n7106), .I2(n7107), .O(n7119));
  LUT3 #(.INIT(8'hE8)) lut_n7120 (.I0(n7115), .I1(n7118), .I2(n7119), .O(n7120));
  LUT3 #(.INIT(8'hE8)) lut_n7121 (.I0(x2556), .I1(x2557), .I2(x2558), .O(n7121));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7122 (.I0(x2547), .I1(x2548), .I2(x2549), .I3(n7116), .I4(n7117), .O(n7122));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7123 (.I0(x2553), .I1(x2554), .I2(x2555), .I3(n7121), .I4(n7122), .O(n7123));
  LUT3 #(.INIT(8'hE8)) lut_n7124 (.I0(x2562), .I1(x2563), .I2(x2564), .O(n7124));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7125 (.I0(x2553), .I1(x2554), .I2(x2555), .I3(n7121), .I4(n7122), .O(n7125));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7126 (.I0(x2559), .I1(x2560), .I2(x2561), .I3(n7124), .I4(n7125), .O(n7126));
  LUT3 #(.INIT(8'h96)) lut_n7127 (.I0(n7115), .I1(n7118), .I2(n7119), .O(n7127));
  LUT3 #(.INIT(8'hE8)) lut_n7128 (.I0(n7123), .I1(n7126), .I2(n7127), .O(n7128));
  LUT3 #(.INIT(8'h96)) lut_n7129 (.I0(n7100), .I1(n7108), .I2(n7109), .O(n7129));
  LUT3 #(.INIT(8'hE8)) lut_n7130 (.I0(n7120), .I1(n7128), .I2(n7129), .O(n7130));
  LUT3 #(.INIT(8'hE8)) lut_n7131 (.I0(x2568), .I1(x2569), .I2(x2570), .O(n7131));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7132 (.I0(x2559), .I1(x2560), .I2(x2561), .I3(n7124), .I4(n7125), .O(n7132));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7133 (.I0(x2565), .I1(x2566), .I2(x2567), .I3(n7131), .I4(n7132), .O(n7133));
  LUT3 #(.INIT(8'hE8)) lut_n7134 (.I0(x2574), .I1(x2575), .I2(x2576), .O(n7134));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7135 (.I0(x2565), .I1(x2566), .I2(x2567), .I3(n7131), .I4(n7132), .O(n7135));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7136 (.I0(x2571), .I1(x2572), .I2(x2573), .I3(n7134), .I4(n7135), .O(n7136));
  LUT3 #(.INIT(8'h96)) lut_n7137 (.I0(n7123), .I1(n7126), .I2(n7127), .O(n7137));
  LUT3 #(.INIT(8'hE8)) lut_n7138 (.I0(n7133), .I1(n7136), .I2(n7137), .O(n7138));
  LUT3 #(.INIT(8'hE8)) lut_n7139 (.I0(x2580), .I1(x2581), .I2(x2582), .O(n7139));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7140 (.I0(x2571), .I1(x2572), .I2(x2573), .I3(n7134), .I4(n7135), .O(n7140));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7141 (.I0(x2577), .I1(x2578), .I2(x2579), .I3(n7139), .I4(n7140), .O(n7141));
  LUT3 #(.INIT(8'hE8)) lut_n7142 (.I0(x2586), .I1(x2587), .I2(x2588), .O(n7142));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7143 (.I0(x2577), .I1(x2578), .I2(x2579), .I3(n7139), .I4(n7140), .O(n7143));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7144 (.I0(x2583), .I1(x2584), .I2(x2585), .I3(n7142), .I4(n7143), .O(n7144));
  LUT3 #(.INIT(8'h96)) lut_n7145 (.I0(n7133), .I1(n7136), .I2(n7137), .O(n7145));
  LUT3 #(.INIT(8'hE8)) lut_n7146 (.I0(n7141), .I1(n7144), .I2(n7145), .O(n7146));
  LUT3 #(.INIT(8'h96)) lut_n7147 (.I0(n7120), .I1(n7128), .I2(n7129), .O(n7147));
  LUT3 #(.INIT(8'hE8)) lut_n7148 (.I0(n7138), .I1(n7146), .I2(n7147), .O(n7148));
  LUT3 #(.INIT(8'h96)) lut_n7149 (.I0(n7092), .I1(n7110), .I2(n7111), .O(n7149));
  LUT3 #(.INIT(8'hE8)) lut_n7150 (.I0(n7130), .I1(n7148), .I2(n7149), .O(n7150));
  LUT3 #(.INIT(8'h96)) lut_n7151 (.I0(n7032), .I1(n7070), .I2(n7071), .O(n7151));
  LUT3 #(.INIT(8'hE8)) lut_n7152 (.I0(n7112), .I1(n7150), .I2(n7151), .O(n7152));
  LUT3 #(.INIT(8'hE8)) lut_n7153 (.I0(x2592), .I1(x2593), .I2(x2594), .O(n7153));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7154 (.I0(x2583), .I1(x2584), .I2(x2585), .I3(n7142), .I4(n7143), .O(n7154));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7155 (.I0(x2589), .I1(x2590), .I2(x2591), .I3(n7153), .I4(n7154), .O(n7155));
  LUT3 #(.INIT(8'hE8)) lut_n7156 (.I0(x2598), .I1(x2599), .I2(x2600), .O(n7156));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7157 (.I0(x2589), .I1(x2590), .I2(x2591), .I3(n7153), .I4(n7154), .O(n7157));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7158 (.I0(x2595), .I1(x2596), .I2(x2597), .I3(n7156), .I4(n7157), .O(n7158));
  LUT3 #(.INIT(8'h96)) lut_n7159 (.I0(n7141), .I1(n7144), .I2(n7145), .O(n7159));
  LUT3 #(.INIT(8'hE8)) lut_n7160 (.I0(n7155), .I1(n7158), .I2(n7159), .O(n7160));
  LUT3 #(.INIT(8'hE8)) lut_n7161 (.I0(x2604), .I1(x2605), .I2(x2606), .O(n7161));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7162 (.I0(x2595), .I1(x2596), .I2(x2597), .I3(n7156), .I4(n7157), .O(n7162));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7163 (.I0(x2601), .I1(x2602), .I2(x2603), .I3(n7161), .I4(n7162), .O(n7163));
  LUT3 #(.INIT(8'hE8)) lut_n7164 (.I0(x2610), .I1(x2611), .I2(x2612), .O(n7164));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7165 (.I0(x2601), .I1(x2602), .I2(x2603), .I3(n7161), .I4(n7162), .O(n7165));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7166 (.I0(x2607), .I1(x2608), .I2(x2609), .I3(n7164), .I4(n7165), .O(n7166));
  LUT3 #(.INIT(8'h96)) lut_n7167 (.I0(n7155), .I1(n7158), .I2(n7159), .O(n7167));
  LUT3 #(.INIT(8'hE8)) lut_n7168 (.I0(n7163), .I1(n7166), .I2(n7167), .O(n7168));
  LUT3 #(.INIT(8'h96)) lut_n7169 (.I0(n7138), .I1(n7146), .I2(n7147), .O(n7169));
  LUT3 #(.INIT(8'hE8)) lut_n7170 (.I0(n7160), .I1(n7168), .I2(n7169), .O(n7170));
  LUT3 #(.INIT(8'hE8)) lut_n7171 (.I0(x2616), .I1(x2617), .I2(x2618), .O(n7171));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7172 (.I0(x2607), .I1(x2608), .I2(x2609), .I3(n7164), .I4(n7165), .O(n7172));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7173 (.I0(x2613), .I1(x2614), .I2(x2615), .I3(n7171), .I4(n7172), .O(n7173));
  LUT3 #(.INIT(8'hE8)) lut_n7174 (.I0(x2622), .I1(x2623), .I2(x2624), .O(n7174));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7175 (.I0(x2613), .I1(x2614), .I2(x2615), .I3(n7171), .I4(n7172), .O(n7175));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7176 (.I0(x2619), .I1(x2620), .I2(x2621), .I3(n7174), .I4(n7175), .O(n7176));
  LUT3 #(.INIT(8'h96)) lut_n7177 (.I0(n7163), .I1(n7166), .I2(n7167), .O(n7177));
  LUT3 #(.INIT(8'hE8)) lut_n7178 (.I0(n7173), .I1(n7176), .I2(n7177), .O(n7178));
  LUT3 #(.INIT(8'hE8)) lut_n7179 (.I0(x2628), .I1(x2629), .I2(x2630), .O(n7179));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7180 (.I0(x2619), .I1(x2620), .I2(x2621), .I3(n7174), .I4(n7175), .O(n7180));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7181 (.I0(x2625), .I1(x2626), .I2(x2627), .I3(n7179), .I4(n7180), .O(n7181));
  LUT3 #(.INIT(8'hE8)) lut_n7182 (.I0(x2634), .I1(x2635), .I2(x2636), .O(n7182));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7183 (.I0(x2625), .I1(x2626), .I2(x2627), .I3(n7179), .I4(n7180), .O(n7183));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7184 (.I0(x2631), .I1(x2632), .I2(x2633), .I3(n7182), .I4(n7183), .O(n7184));
  LUT3 #(.INIT(8'h96)) lut_n7185 (.I0(n7173), .I1(n7176), .I2(n7177), .O(n7185));
  LUT3 #(.INIT(8'hE8)) lut_n7186 (.I0(n7181), .I1(n7184), .I2(n7185), .O(n7186));
  LUT3 #(.INIT(8'h96)) lut_n7187 (.I0(n7160), .I1(n7168), .I2(n7169), .O(n7187));
  LUT3 #(.INIT(8'hE8)) lut_n7188 (.I0(n7178), .I1(n7186), .I2(n7187), .O(n7188));
  LUT3 #(.INIT(8'h96)) lut_n7189 (.I0(n7130), .I1(n7148), .I2(n7149), .O(n7189));
  LUT3 #(.INIT(8'hE8)) lut_n7190 (.I0(n7170), .I1(n7188), .I2(n7189), .O(n7190));
  LUT3 #(.INIT(8'hE8)) lut_n7191 (.I0(x2640), .I1(x2641), .I2(x2642), .O(n7191));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7192 (.I0(x2631), .I1(x2632), .I2(x2633), .I3(n7182), .I4(n7183), .O(n7192));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7193 (.I0(x2637), .I1(x2638), .I2(x2639), .I3(n7191), .I4(n7192), .O(n7193));
  LUT3 #(.INIT(8'hE8)) lut_n7194 (.I0(x2646), .I1(x2647), .I2(x2648), .O(n7194));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7195 (.I0(x2637), .I1(x2638), .I2(x2639), .I3(n7191), .I4(n7192), .O(n7195));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7196 (.I0(x2643), .I1(x2644), .I2(x2645), .I3(n7194), .I4(n7195), .O(n7196));
  LUT3 #(.INIT(8'h96)) lut_n7197 (.I0(n7181), .I1(n7184), .I2(n7185), .O(n7197));
  LUT3 #(.INIT(8'hE8)) lut_n7198 (.I0(n7193), .I1(n7196), .I2(n7197), .O(n7198));
  LUT3 #(.INIT(8'hE8)) lut_n7199 (.I0(x2652), .I1(x2653), .I2(x2654), .O(n7199));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7200 (.I0(x2643), .I1(x2644), .I2(x2645), .I3(n7194), .I4(n7195), .O(n7200));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7201 (.I0(x2649), .I1(x2650), .I2(x2651), .I3(n7199), .I4(n7200), .O(n7201));
  LUT3 #(.INIT(8'hE8)) lut_n7202 (.I0(x2658), .I1(x2659), .I2(x2660), .O(n7202));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7203 (.I0(x2649), .I1(x2650), .I2(x2651), .I3(n7199), .I4(n7200), .O(n7203));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7204 (.I0(x2655), .I1(x2656), .I2(x2657), .I3(n7202), .I4(n7203), .O(n7204));
  LUT3 #(.INIT(8'h96)) lut_n7205 (.I0(n7193), .I1(n7196), .I2(n7197), .O(n7205));
  LUT3 #(.INIT(8'hE8)) lut_n7206 (.I0(n7201), .I1(n7204), .I2(n7205), .O(n7206));
  LUT3 #(.INIT(8'h96)) lut_n7207 (.I0(n7178), .I1(n7186), .I2(n7187), .O(n7207));
  LUT3 #(.INIT(8'hE8)) lut_n7208 (.I0(n7198), .I1(n7206), .I2(n7207), .O(n7208));
  LUT3 #(.INIT(8'hE8)) lut_n7209 (.I0(x2664), .I1(x2665), .I2(x2666), .O(n7209));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7210 (.I0(x2655), .I1(x2656), .I2(x2657), .I3(n7202), .I4(n7203), .O(n7210));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7211 (.I0(x2661), .I1(x2662), .I2(x2663), .I3(n7209), .I4(n7210), .O(n7211));
  LUT3 #(.INIT(8'hE8)) lut_n7212 (.I0(x2670), .I1(x2671), .I2(x2672), .O(n7212));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7213 (.I0(x2661), .I1(x2662), .I2(x2663), .I3(n7209), .I4(n7210), .O(n7213));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7214 (.I0(x2667), .I1(x2668), .I2(x2669), .I3(n7212), .I4(n7213), .O(n7214));
  LUT3 #(.INIT(8'h96)) lut_n7215 (.I0(n7201), .I1(n7204), .I2(n7205), .O(n7215));
  LUT3 #(.INIT(8'hE8)) lut_n7216 (.I0(n7211), .I1(n7214), .I2(n7215), .O(n7216));
  LUT3 #(.INIT(8'hE8)) lut_n7217 (.I0(x2676), .I1(x2677), .I2(x2678), .O(n7217));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7218 (.I0(x2667), .I1(x2668), .I2(x2669), .I3(n7212), .I4(n7213), .O(n7218));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7219 (.I0(x2673), .I1(x2674), .I2(x2675), .I3(n7217), .I4(n7218), .O(n7219));
  LUT3 #(.INIT(8'hE8)) lut_n7220 (.I0(x2682), .I1(x2683), .I2(x2684), .O(n7220));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7221 (.I0(x2673), .I1(x2674), .I2(x2675), .I3(n7217), .I4(n7218), .O(n7221));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7222 (.I0(x2679), .I1(x2680), .I2(x2681), .I3(n7220), .I4(n7221), .O(n7222));
  LUT3 #(.INIT(8'h96)) lut_n7223 (.I0(n7211), .I1(n7214), .I2(n7215), .O(n7223));
  LUT3 #(.INIT(8'hE8)) lut_n7224 (.I0(n7219), .I1(n7222), .I2(n7223), .O(n7224));
  LUT3 #(.INIT(8'h96)) lut_n7225 (.I0(n7198), .I1(n7206), .I2(n7207), .O(n7225));
  LUT3 #(.INIT(8'hE8)) lut_n7226 (.I0(n7216), .I1(n7224), .I2(n7225), .O(n7226));
  LUT3 #(.INIT(8'h96)) lut_n7227 (.I0(n7170), .I1(n7188), .I2(n7189), .O(n7227));
  LUT3 #(.INIT(8'hE8)) lut_n7228 (.I0(n7208), .I1(n7226), .I2(n7227), .O(n7228));
  LUT3 #(.INIT(8'h96)) lut_n7229 (.I0(n7112), .I1(n7150), .I2(n7151), .O(n7229));
  LUT3 #(.INIT(8'hE8)) lut_n7230 (.I0(n7190), .I1(n7228), .I2(n7229), .O(n7230));
  LUT3 #(.INIT(8'h96)) lut_n7231 (.I0(n6994), .I1(n7072), .I2(n7073), .O(n7231));
  LUT3 #(.INIT(8'hE8)) lut_n7232 (.I0(n7152), .I1(n7230), .I2(n7231), .O(n7232));
  LUT3 #(.INIT(8'h96)) lut_n7233 (.I0(n6754), .I1(n6912), .I2(n6913), .O(n7233));
  LUT3 #(.INIT(8'hE8)) lut_n7234 (.I0(n7074), .I1(n7232), .I2(n7233), .O(n7234));
  LUT3 #(.INIT(8'hE8)) lut_n7235 (.I0(x2688), .I1(x2689), .I2(x2690), .O(n7235));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7236 (.I0(x2679), .I1(x2680), .I2(x2681), .I3(n7220), .I4(n7221), .O(n7236));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7237 (.I0(x2685), .I1(x2686), .I2(x2687), .I3(n7235), .I4(n7236), .O(n7237));
  LUT3 #(.INIT(8'hE8)) lut_n7238 (.I0(x2694), .I1(x2695), .I2(x2696), .O(n7238));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7239 (.I0(x2685), .I1(x2686), .I2(x2687), .I3(n7235), .I4(n7236), .O(n7239));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7240 (.I0(x2691), .I1(x2692), .I2(x2693), .I3(n7238), .I4(n7239), .O(n7240));
  LUT3 #(.INIT(8'h96)) lut_n7241 (.I0(n7219), .I1(n7222), .I2(n7223), .O(n7241));
  LUT3 #(.INIT(8'hE8)) lut_n7242 (.I0(n7237), .I1(n7240), .I2(n7241), .O(n7242));
  LUT3 #(.INIT(8'hE8)) lut_n7243 (.I0(x2700), .I1(x2701), .I2(x2702), .O(n7243));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7244 (.I0(x2691), .I1(x2692), .I2(x2693), .I3(n7238), .I4(n7239), .O(n7244));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7245 (.I0(x2697), .I1(x2698), .I2(x2699), .I3(n7243), .I4(n7244), .O(n7245));
  LUT3 #(.INIT(8'hE8)) lut_n7246 (.I0(x2706), .I1(x2707), .I2(x2708), .O(n7246));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7247 (.I0(x2697), .I1(x2698), .I2(x2699), .I3(n7243), .I4(n7244), .O(n7247));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7248 (.I0(x2703), .I1(x2704), .I2(x2705), .I3(n7246), .I4(n7247), .O(n7248));
  LUT3 #(.INIT(8'h96)) lut_n7249 (.I0(n7237), .I1(n7240), .I2(n7241), .O(n7249));
  LUT3 #(.INIT(8'hE8)) lut_n7250 (.I0(n7245), .I1(n7248), .I2(n7249), .O(n7250));
  LUT3 #(.INIT(8'h96)) lut_n7251 (.I0(n7216), .I1(n7224), .I2(n7225), .O(n7251));
  LUT3 #(.INIT(8'hE8)) lut_n7252 (.I0(n7242), .I1(n7250), .I2(n7251), .O(n7252));
  LUT3 #(.INIT(8'hE8)) lut_n7253 (.I0(x2712), .I1(x2713), .I2(x2714), .O(n7253));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7254 (.I0(x2703), .I1(x2704), .I2(x2705), .I3(n7246), .I4(n7247), .O(n7254));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7255 (.I0(x2709), .I1(x2710), .I2(x2711), .I3(n7253), .I4(n7254), .O(n7255));
  LUT3 #(.INIT(8'hE8)) lut_n7256 (.I0(x2718), .I1(x2719), .I2(x2720), .O(n7256));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7257 (.I0(x2709), .I1(x2710), .I2(x2711), .I3(n7253), .I4(n7254), .O(n7257));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7258 (.I0(x2715), .I1(x2716), .I2(x2717), .I3(n7256), .I4(n7257), .O(n7258));
  LUT3 #(.INIT(8'h96)) lut_n7259 (.I0(n7245), .I1(n7248), .I2(n7249), .O(n7259));
  LUT3 #(.INIT(8'hE8)) lut_n7260 (.I0(n7255), .I1(n7258), .I2(n7259), .O(n7260));
  LUT3 #(.INIT(8'hE8)) lut_n7261 (.I0(x2724), .I1(x2725), .I2(x2726), .O(n7261));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7262 (.I0(x2715), .I1(x2716), .I2(x2717), .I3(n7256), .I4(n7257), .O(n7262));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7263 (.I0(x2721), .I1(x2722), .I2(x2723), .I3(n7261), .I4(n7262), .O(n7263));
  LUT3 #(.INIT(8'hE8)) lut_n7264 (.I0(x2730), .I1(x2731), .I2(x2732), .O(n7264));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7265 (.I0(x2721), .I1(x2722), .I2(x2723), .I3(n7261), .I4(n7262), .O(n7265));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7266 (.I0(x2727), .I1(x2728), .I2(x2729), .I3(n7264), .I4(n7265), .O(n7266));
  LUT3 #(.INIT(8'h96)) lut_n7267 (.I0(n7255), .I1(n7258), .I2(n7259), .O(n7267));
  LUT3 #(.INIT(8'hE8)) lut_n7268 (.I0(n7263), .I1(n7266), .I2(n7267), .O(n7268));
  LUT3 #(.INIT(8'h96)) lut_n7269 (.I0(n7242), .I1(n7250), .I2(n7251), .O(n7269));
  LUT3 #(.INIT(8'hE8)) lut_n7270 (.I0(n7260), .I1(n7268), .I2(n7269), .O(n7270));
  LUT3 #(.INIT(8'h96)) lut_n7271 (.I0(n7208), .I1(n7226), .I2(n7227), .O(n7271));
  LUT3 #(.INIT(8'hE8)) lut_n7272 (.I0(n7252), .I1(n7270), .I2(n7271), .O(n7272));
  LUT3 #(.INIT(8'hE8)) lut_n7273 (.I0(x2736), .I1(x2737), .I2(x2738), .O(n7273));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7274 (.I0(x2727), .I1(x2728), .I2(x2729), .I3(n7264), .I4(n7265), .O(n7274));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7275 (.I0(x2733), .I1(x2734), .I2(x2735), .I3(n7273), .I4(n7274), .O(n7275));
  LUT3 #(.INIT(8'hE8)) lut_n7276 (.I0(x2742), .I1(x2743), .I2(x2744), .O(n7276));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7277 (.I0(x2733), .I1(x2734), .I2(x2735), .I3(n7273), .I4(n7274), .O(n7277));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7278 (.I0(x2739), .I1(x2740), .I2(x2741), .I3(n7276), .I4(n7277), .O(n7278));
  LUT3 #(.INIT(8'h96)) lut_n7279 (.I0(n7263), .I1(n7266), .I2(n7267), .O(n7279));
  LUT3 #(.INIT(8'hE8)) lut_n7280 (.I0(n7275), .I1(n7278), .I2(n7279), .O(n7280));
  LUT3 #(.INIT(8'hE8)) lut_n7281 (.I0(x2748), .I1(x2749), .I2(x2750), .O(n7281));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7282 (.I0(x2739), .I1(x2740), .I2(x2741), .I3(n7276), .I4(n7277), .O(n7282));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7283 (.I0(x2745), .I1(x2746), .I2(x2747), .I3(n7281), .I4(n7282), .O(n7283));
  LUT3 #(.INIT(8'hE8)) lut_n7284 (.I0(x2754), .I1(x2755), .I2(x2756), .O(n7284));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7285 (.I0(x2745), .I1(x2746), .I2(x2747), .I3(n7281), .I4(n7282), .O(n7285));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7286 (.I0(x2751), .I1(x2752), .I2(x2753), .I3(n7284), .I4(n7285), .O(n7286));
  LUT3 #(.INIT(8'h96)) lut_n7287 (.I0(n7275), .I1(n7278), .I2(n7279), .O(n7287));
  LUT3 #(.INIT(8'hE8)) lut_n7288 (.I0(n7283), .I1(n7286), .I2(n7287), .O(n7288));
  LUT3 #(.INIT(8'h96)) lut_n7289 (.I0(n7260), .I1(n7268), .I2(n7269), .O(n7289));
  LUT3 #(.INIT(8'hE8)) lut_n7290 (.I0(n7280), .I1(n7288), .I2(n7289), .O(n7290));
  LUT3 #(.INIT(8'hE8)) lut_n7291 (.I0(x2760), .I1(x2761), .I2(x2762), .O(n7291));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7292 (.I0(x2751), .I1(x2752), .I2(x2753), .I3(n7284), .I4(n7285), .O(n7292));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7293 (.I0(x2757), .I1(x2758), .I2(x2759), .I3(n7291), .I4(n7292), .O(n7293));
  LUT3 #(.INIT(8'hE8)) lut_n7294 (.I0(x2766), .I1(x2767), .I2(x2768), .O(n7294));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7295 (.I0(x2757), .I1(x2758), .I2(x2759), .I3(n7291), .I4(n7292), .O(n7295));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7296 (.I0(x2763), .I1(x2764), .I2(x2765), .I3(n7294), .I4(n7295), .O(n7296));
  LUT3 #(.INIT(8'h96)) lut_n7297 (.I0(n7283), .I1(n7286), .I2(n7287), .O(n7297));
  LUT3 #(.INIT(8'hE8)) lut_n7298 (.I0(n7293), .I1(n7296), .I2(n7297), .O(n7298));
  LUT3 #(.INIT(8'hE8)) lut_n7299 (.I0(x2772), .I1(x2773), .I2(x2774), .O(n7299));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7300 (.I0(x2763), .I1(x2764), .I2(x2765), .I3(n7294), .I4(n7295), .O(n7300));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7301 (.I0(x2769), .I1(x2770), .I2(x2771), .I3(n7299), .I4(n7300), .O(n7301));
  LUT3 #(.INIT(8'hE8)) lut_n7302 (.I0(x2778), .I1(x2779), .I2(x2780), .O(n7302));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7303 (.I0(x2769), .I1(x2770), .I2(x2771), .I3(n7299), .I4(n7300), .O(n7303));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7304 (.I0(x2775), .I1(x2776), .I2(x2777), .I3(n7302), .I4(n7303), .O(n7304));
  LUT3 #(.INIT(8'h96)) lut_n7305 (.I0(n7293), .I1(n7296), .I2(n7297), .O(n7305));
  LUT3 #(.INIT(8'hE8)) lut_n7306 (.I0(n7301), .I1(n7304), .I2(n7305), .O(n7306));
  LUT3 #(.INIT(8'h96)) lut_n7307 (.I0(n7280), .I1(n7288), .I2(n7289), .O(n7307));
  LUT3 #(.INIT(8'hE8)) lut_n7308 (.I0(n7298), .I1(n7306), .I2(n7307), .O(n7308));
  LUT3 #(.INIT(8'h96)) lut_n7309 (.I0(n7252), .I1(n7270), .I2(n7271), .O(n7309));
  LUT3 #(.INIT(8'hE8)) lut_n7310 (.I0(n7290), .I1(n7308), .I2(n7309), .O(n7310));
  LUT3 #(.INIT(8'h96)) lut_n7311 (.I0(n7190), .I1(n7228), .I2(n7229), .O(n7311));
  LUT3 #(.INIT(8'hE8)) lut_n7312 (.I0(n7272), .I1(n7310), .I2(n7311), .O(n7312));
  LUT3 #(.INIT(8'hE8)) lut_n7313 (.I0(x2784), .I1(x2785), .I2(x2786), .O(n7313));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7314 (.I0(x2775), .I1(x2776), .I2(x2777), .I3(n7302), .I4(n7303), .O(n7314));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7315 (.I0(x2781), .I1(x2782), .I2(x2783), .I3(n7313), .I4(n7314), .O(n7315));
  LUT3 #(.INIT(8'hE8)) lut_n7316 (.I0(x2790), .I1(x2791), .I2(x2792), .O(n7316));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7317 (.I0(x2781), .I1(x2782), .I2(x2783), .I3(n7313), .I4(n7314), .O(n7317));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7318 (.I0(x2787), .I1(x2788), .I2(x2789), .I3(n7316), .I4(n7317), .O(n7318));
  LUT3 #(.INIT(8'h96)) lut_n7319 (.I0(n7301), .I1(n7304), .I2(n7305), .O(n7319));
  LUT3 #(.INIT(8'hE8)) lut_n7320 (.I0(n7315), .I1(n7318), .I2(n7319), .O(n7320));
  LUT3 #(.INIT(8'hE8)) lut_n7321 (.I0(x2796), .I1(x2797), .I2(x2798), .O(n7321));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7322 (.I0(x2787), .I1(x2788), .I2(x2789), .I3(n7316), .I4(n7317), .O(n7322));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7323 (.I0(x2793), .I1(x2794), .I2(x2795), .I3(n7321), .I4(n7322), .O(n7323));
  LUT3 #(.INIT(8'hE8)) lut_n7324 (.I0(x2802), .I1(x2803), .I2(x2804), .O(n7324));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7325 (.I0(x2793), .I1(x2794), .I2(x2795), .I3(n7321), .I4(n7322), .O(n7325));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7326 (.I0(x2799), .I1(x2800), .I2(x2801), .I3(n7324), .I4(n7325), .O(n7326));
  LUT3 #(.INIT(8'h96)) lut_n7327 (.I0(n7315), .I1(n7318), .I2(n7319), .O(n7327));
  LUT3 #(.INIT(8'hE8)) lut_n7328 (.I0(n7323), .I1(n7326), .I2(n7327), .O(n7328));
  LUT3 #(.INIT(8'h96)) lut_n7329 (.I0(n7298), .I1(n7306), .I2(n7307), .O(n7329));
  LUT3 #(.INIT(8'hE8)) lut_n7330 (.I0(n7320), .I1(n7328), .I2(n7329), .O(n7330));
  LUT3 #(.INIT(8'hE8)) lut_n7331 (.I0(x2808), .I1(x2809), .I2(x2810), .O(n7331));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7332 (.I0(x2799), .I1(x2800), .I2(x2801), .I3(n7324), .I4(n7325), .O(n7332));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7333 (.I0(x2805), .I1(x2806), .I2(x2807), .I3(n7331), .I4(n7332), .O(n7333));
  LUT3 #(.INIT(8'hE8)) lut_n7334 (.I0(x2814), .I1(x2815), .I2(x2816), .O(n7334));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7335 (.I0(x2805), .I1(x2806), .I2(x2807), .I3(n7331), .I4(n7332), .O(n7335));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7336 (.I0(x2811), .I1(x2812), .I2(x2813), .I3(n7334), .I4(n7335), .O(n7336));
  LUT3 #(.INIT(8'h96)) lut_n7337 (.I0(n7323), .I1(n7326), .I2(n7327), .O(n7337));
  LUT3 #(.INIT(8'hE8)) lut_n7338 (.I0(n7333), .I1(n7336), .I2(n7337), .O(n7338));
  LUT3 #(.INIT(8'hE8)) lut_n7339 (.I0(x2820), .I1(x2821), .I2(x2822), .O(n7339));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7340 (.I0(x2811), .I1(x2812), .I2(x2813), .I3(n7334), .I4(n7335), .O(n7340));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7341 (.I0(x2817), .I1(x2818), .I2(x2819), .I3(n7339), .I4(n7340), .O(n7341));
  LUT3 #(.INIT(8'hE8)) lut_n7342 (.I0(x2826), .I1(x2827), .I2(x2828), .O(n7342));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7343 (.I0(x2817), .I1(x2818), .I2(x2819), .I3(n7339), .I4(n7340), .O(n7343));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7344 (.I0(x2823), .I1(x2824), .I2(x2825), .I3(n7342), .I4(n7343), .O(n7344));
  LUT3 #(.INIT(8'h96)) lut_n7345 (.I0(n7333), .I1(n7336), .I2(n7337), .O(n7345));
  LUT3 #(.INIT(8'hE8)) lut_n7346 (.I0(n7341), .I1(n7344), .I2(n7345), .O(n7346));
  LUT3 #(.INIT(8'h96)) lut_n7347 (.I0(n7320), .I1(n7328), .I2(n7329), .O(n7347));
  LUT3 #(.INIT(8'hE8)) lut_n7348 (.I0(n7338), .I1(n7346), .I2(n7347), .O(n7348));
  LUT3 #(.INIT(8'h96)) lut_n7349 (.I0(n7290), .I1(n7308), .I2(n7309), .O(n7349));
  LUT3 #(.INIT(8'hE8)) lut_n7350 (.I0(n7330), .I1(n7348), .I2(n7349), .O(n7350));
  LUT3 #(.INIT(8'hE8)) lut_n7351 (.I0(x2832), .I1(x2833), .I2(x2834), .O(n7351));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7352 (.I0(x2823), .I1(x2824), .I2(x2825), .I3(n7342), .I4(n7343), .O(n7352));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7353 (.I0(x2829), .I1(x2830), .I2(x2831), .I3(n7351), .I4(n7352), .O(n7353));
  LUT3 #(.INIT(8'hE8)) lut_n7354 (.I0(x2838), .I1(x2839), .I2(x2840), .O(n7354));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7355 (.I0(x2829), .I1(x2830), .I2(x2831), .I3(n7351), .I4(n7352), .O(n7355));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7356 (.I0(x2835), .I1(x2836), .I2(x2837), .I3(n7354), .I4(n7355), .O(n7356));
  LUT3 #(.INIT(8'h96)) lut_n7357 (.I0(n7341), .I1(n7344), .I2(n7345), .O(n7357));
  LUT3 #(.INIT(8'hE8)) lut_n7358 (.I0(n7353), .I1(n7356), .I2(n7357), .O(n7358));
  LUT3 #(.INIT(8'hE8)) lut_n7359 (.I0(x2844), .I1(x2845), .I2(x2846), .O(n7359));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7360 (.I0(x2835), .I1(x2836), .I2(x2837), .I3(n7354), .I4(n7355), .O(n7360));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7361 (.I0(x2841), .I1(x2842), .I2(x2843), .I3(n7359), .I4(n7360), .O(n7361));
  LUT3 #(.INIT(8'hE8)) lut_n7362 (.I0(x2850), .I1(x2851), .I2(x2852), .O(n7362));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7363 (.I0(x2841), .I1(x2842), .I2(x2843), .I3(n7359), .I4(n7360), .O(n7363));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7364 (.I0(x2847), .I1(x2848), .I2(x2849), .I3(n7362), .I4(n7363), .O(n7364));
  LUT3 #(.INIT(8'h96)) lut_n7365 (.I0(n7353), .I1(n7356), .I2(n7357), .O(n7365));
  LUT3 #(.INIT(8'hE8)) lut_n7366 (.I0(n7361), .I1(n7364), .I2(n7365), .O(n7366));
  LUT3 #(.INIT(8'h96)) lut_n7367 (.I0(n7338), .I1(n7346), .I2(n7347), .O(n7367));
  LUT3 #(.INIT(8'hE8)) lut_n7368 (.I0(n7358), .I1(n7366), .I2(n7367), .O(n7368));
  LUT3 #(.INIT(8'hE8)) lut_n7369 (.I0(x2856), .I1(x2857), .I2(x2858), .O(n7369));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7370 (.I0(x2847), .I1(x2848), .I2(x2849), .I3(n7362), .I4(n7363), .O(n7370));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7371 (.I0(x2853), .I1(x2854), .I2(x2855), .I3(n7369), .I4(n7370), .O(n7371));
  LUT3 #(.INIT(8'hE8)) lut_n7372 (.I0(x2862), .I1(x2863), .I2(x2864), .O(n7372));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7373 (.I0(x2853), .I1(x2854), .I2(x2855), .I3(n7369), .I4(n7370), .O(n7373));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7374 (.I0(x2859), .I1(x2860), .I2(x2861), .I3(n7372), .I4(n7373), .O(n7374));
  LUT3 #(.INIT(8'h96)) lut_n7375 (.I0(n7361), .I1(n7364), .I2(n7365), .O(n7375));
  LUT3 #(.INIT(8'hE8)) lut_n7376 (.I0(n7371), .I1(n7374), .I2(n7375), .O(n7376));
  LUT3 #(.INIT(8'hE8)) lut_n7377 (.I0(x2868), .I1(x2869), .I2(x2870), .O(n7377));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7378 (.I0(x2859), .I1(x2860), .I2(x2861), .I3(n7372), .I4(n7373), .O(n7378));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7379 (.I0(x2865), .I1(x2866), .I2(x2867), .I3(n7377), .I4(n7378), .O(n7379));
  LUT3 #(.INIT(8'hE8)) lut_n7380 (.I0(x2874), .I1(x2875), .I2(x2876), .O(n7380));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7381 (.I0(x2865), .I1(x2866), .I2(x2867), .I3(n7377), .I4(n7378), .O(n7381));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7382 (.I0(x2871), .I1(x2872), .I2(x2873), .I3(n7380), .I4(n7381), .O(n7382));
  LUT3 #(.INIT(8'h96)) lut_n7383 (.I0(n7371), .I1(n7374), .I2(n7375), .O(n7383));
  LUT3 #(.INIT(8'hE8)) lut_n7384 (.I0(n7379), .I1(n7382), .I2(n7383), .O(n7384));
  LUT3 #(.INIT(8'h96)) lut_n7385 (.I0(n7358), .I1(n7366), .I2(n7367), .O(n7385));
  LUT3 #(.INIT(8'hE8)) lut_n7386 (.I0(n7376), .I1(n7384), .I2(n7385), .O(n7386));
  LUT3 #(.INIT(8'h96)) lut_n7387 (.I0(n7330), .I1(n7348), .I2(n7349), .O(n7387));
  LUT3 #(.INIT(8'hE8)) lut_n7388 (.I0(n7368), .I1(n7386), .I2(n7387), .O(n7388));
  LUT3 #(.INIT(8'h96)) lut_n7389 (.I0(n7272), .I1(n7310), .I2(n7311), .O(n7389));
  LUT3 #(.INIT(8'hE8)) lut_n7390 (.I0(n7350), .I1(n7388), .I2(n7389), .O(n7390));
  LUT3 #(.INIT(8'h96)) lut_n7391 (.I0(n7152), .I1(n7230), .I2(n7231), .O(n7391));
  LUT3 #(.INIT(8'hE8)) lut_n7392 (.I0(n7312), .I1(n7390), .I2(n7391), .O(n7392));
  LUT3 #(.INIT(8'hE8)) lut_n7393 (.I0(x2880), .I1(x2881), .I2(x2882), .O(n7393));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7394 (.I0(x2871), .I1(x2872), .I2(x2873), .I3(n7380), .I4(n7381), .O(n7394));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7395 (.I0(x2877), .I1(x2878), .I2(x2879), .I3(n7393), .I4(n7394), .O(n7395));
  LUT3 #(.INIT(8'hE8)) lut_n7396 (.I0(x2886), .I1(x2887), .I2(x2888), .O(n7396));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7397 (.I0(x2877), .I1(x2878), .I2(x2879), .I3(n7393), .I4(n7394), .O(n7397));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7398 (.I0(x2883), .I1(x2884), .I2(x2885), .I3(n7396), .I4(n7397), .O(n7398));
  LUT3 #(.INIT(8'h96)) lut_n7399 (.I0(n7379), .I1(n7382), .I2(n7383), .O(n7399));
  LUT3 #(.INIT(8'hE8)) lut_n7400 (.I0(n7395), .I1(n7398), .I2(n7399), .O(n7400));
  LUT3 #(.INIT(8'hE8)) lut_n7401 (.I0(x2892), .I1(x2893), .I2(x2894), .O(n7401));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7402 (.I0(x2883), .I1(x2884), .I2(x2885), .I3(n7396), .I4(n7397), .O(n7402));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7403 (.I0(x2889), .I1(x2890), .I2(x2891), .I3(n7401), .I4(n7402), .O(n7403));
  LUT3 #(.INIT(8'hE8)) lut_n7404 (.I0(x2898), .I1(x2899), .I2(x2900), .O(n7404));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7405 (.I0(x2889), .I1(x2890), .I2(x2891), .I3(n7401), .I4(n7402), .O(n7405));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7406 (.I0(x2895), .I1(x2896), .I2(x2897), .I3(n7404), .I4(n7405), .O(n7406));
  LUT3 #(.INIT(8'h96)) lut_n7407 (.I0(n7395), .I1(n7398), .I2(n7399), .O(n7407));
  LUT3 #(.INIT(8'hE8)) lut_n7408 (.I0(n7403), .I1(n7406), .I2(n7407), .O(n7408));
  LUT3 #(.INIT(8'h96)) lut_n7409 (.I0(n7376), .I1(n7384), .I2(n7385), .O(n7409));
  LUT3 #(.INIT(8'hE8)) lut_n7410 (.I0(n7400), .I1(n7408), .I2(n7409), .O(n7410));
  LUT3 #(.INIT(8'hE8)) lut_n7411 (.I0(x2904), .I1(x2905), .I2(x2906), .O(n7411));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7412 (.I0(x2895), .I1(x2896), .I2(x2897), .I3(n7404), .I4(n7405), .O(n7412));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7413 (.I0(x2901), .I1(x2902), .I2(x2903), .I3(n7411), .I4(n7412), .O(n7413));
  LUT3 #(.INIT(8'hE8)) lut_n7414 (.I0(x2910), .I1(x2911), .I2(x2912), .O(n7414));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7415 (.I0(x2901), .I1(x2902), .I2(x2903), .I3(n7411), .I4(n7412), .O(n7415));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7416 (.I0(x2907), .I1(x2908), .I2(x2909), .I3(n7414), .I4(n7415), .O(n7416));
  LUT3 #(.INIT(8'h96)) lut_n7417 (.I0(n7403), .I1(n7406), .I2(n7407), .O(n7417));
  LUT3 #(.INIT(8'hE8)) lut_n7418 (.I0(n7413), .I1(n7416), .I2(n7417), .O(n7418));
  LUT3 #(.INIT(8'hE8)) lut_n7419 (.I0(x2916), .I1(x2917), .I2(x2918), .O(n7419));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7420 (.I0(x2907), .I1(x2908), .I2(x2909), .I3(n7414), .I4(n7415), .O(n7420));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7421 (.I0(x2913), .I1(x2914), .I2(x2915), .I3(n7419), .I4(n7420), .O(n7421));
  LUT3 #(.INIT(8'hE8)) lut_n7422 (.I0(x2922), .I1(x2923), .I2(x2924), .O(n7422));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7423 (.I0(x2913), .I1(x2914), .I2(x2915), .I3(n7419), .I4(n7420), .O(n7423));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7424 (.I0(x2919), .I1(x2920), .I2(x2921), .I3(n7422), .I4(n7423), .O(n7424));
  LUT3 #(.INIT(8'h96)) lut_n7425 (.I0(n7413), .I1(n7416), .I2(n7417), .O(n7425));
  LUT3 #(.INIT(8'hE8)) lut_n7426 (.I0(n7421), .I1(n7424), .I2(n7425), .O(n7426));
  LUT3 #(.INIT(8'h96)) lut_n7427 (.I0(n7400), .I1(n7408), .I2(n7409), .O(n7427));
  LUT3 #(.INIT(8'hE8)) lut_n7428 (.I0(n7418), .I1(n7426), .I2(n7427), .O(n7428));
  LUT3 #(.INIT(8'h96)) lut_n7429 (.I0(n7368), .I1(n7386), .I2(n7387), .O(n7429));
  LUT3 #(.INIT(8'hE8)) lut_n7430 (.I0(n7410), .I1(n7428), .I2(n7429), .O(n7430));
  LUT3 #(.INIT(8'hE8)) lut_n7431 (.I0(x2928), .I1(x2929), .I2(x2930), .O(n7431));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7432 (.I0(x2919), .I1(x2920), .I2(x2921), .I3(n7422), .I4(n7423), .O(n7432));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7433 (.I0(x2925), .I1(x2926), .I2(x2927), .I3(n7431), .I4(n7432), .O(n7433));
  LUT3 #(.INIT(8'hE8)) lut_n7434 (.I0(x2934), .I1(x2935), .I2(x2936), .O(n7434));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7435 (.I0(x2925), .I1(x2926), .I2(x2927), .I3(n7431), .I4(n7432), .O(n7435));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7436 (.I0(x2931), .I1(x2932), .I2(x2933), .I3(n7434), .I4(n7435), .O(n7436));
  LUT3 #(.INIT(8'h96)) lut_n7437 (.I0(n7421), .I1(n7424), .I2(n7425), .O(n7437));
  LUT3 #(.INIT(8'hE8)) lut_n7438 (.I0(n7433), .I1(n7436), .I2(n7437), .O(n7438));
  LUT3 #(.INIT(8'hE8)) lut_n7439 (.I0(x2940), .I1(x2941), .I2(x2942), .O(n7439));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7440 (.I0(x2931), .I1(x2932), .I2(x2933), .I3(n7434), .I4(n7435), .O(n7440));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7441 (.I0(x2937), .I1(x2938), .I2(x2939), .I3(n7439), .I4(n7440), .O(n7441));
  LUT3 #(.INIT(8'hE8)) lut_n7442 (.I0(x2946), .I1(x2947), .I2(x2948), .O(n7442));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7443 (.I0(x2937), .I1(x2938), .I2(x2939), .I3(n7439), .I4(n7440), .O(n7443));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7444 (.I0(x2943), .I1(x2944), .I2(x2945), .I3(n7442), .I4(n7443), .O(n7444));
  LUT3 #(.INIT(8'h96)) lut_n7445 (.I0(n7433), .I1(n7436), .I2(n7437), .O(n7445));
  LUT3 #(.INIT(8'hE8)) lut_n7446 (.I0(n7441), .I1(n7444), .I2(n7445), .O(n7446));
  LUT3 #(.INIT(8'h96)) lut_n7447 (.I0(n7418), .I1(n7426), .I2(n7427), .O(n7447));
  LUT3 #(.INIT(8'hE8)) lut_n7448 (.I0(n7438), .I1(n7446), .I2(n7447), .O(n7448));
  LUT3 #(.INIT(8'hE8)) lut_n7449 (.I0(x2952), .I1(x2953), .I2(x2954), .O(n7449));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7450 (.I0(x2943), .I1(x2944), .I2(x2945), .I3(n7442), .I4(n7443), .O(n7450));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7451 (.I0(x2949), .I1(x2950), .I2(x2951), .I3(n7449), .I4(n7450), .O(n7451));
  LUT3 #(.INIT(8'hE8)) lut_n7452 (.I0(x2958), .I1(x2959), .I2(x2960), .O(n7452));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7453 (.I0(x2949), .I1(x2950), .I2(x2951), .I3(n7449), .I4(n7450), .O(n7453));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7454 (.I0(x2955), .I1(x2956), .I2(x2957), .I3(n7452), .I4(n7453), .O(n7454));
  LUT3 #(.INIT(8'h96)) lut_n7455 (.I0(n7441), .I1(n7444), .I2(n7445), .O(n7455));
  LUT3 #(.INIT(8'hE8)) lut_n7456 (.I0(n7451), .I1(n7454), .I2(n7455), .O(n7456));
  LUT3 #(.INIT(8'hE8)) lut_n7457 (.I0(x2964), .I1(x2965), .I2(x2966), .O(n7457));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7458 (.I0(x2955), .I1(x2956), .I2(x2957), .I3(n7452), .I4(n7453), .O(n7458));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7459 (.I0(x2961), .I1(x2962), .I2(x2963), .I3(n7457), .I4(n7458), .O(n7459));
  LUT3 #(.INIT(8'hE8)) lut_n7460 (.I0(x2970), .I1(x2971), .I2(x2972), .O(n7460));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7461 (.I0(x2961), .I1(x2962), .I2(x2963), .I3(n7457), .I4(n7458), .O(n7461));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7462 (.I0(x2967), .I1(x2968), .I2(x2969), .I3(n7460), .I4(n7461), .O(n7462));
  LUT3 #(.INIT(8'h96)) lut_n7463 (.I0(n7451), .I1(n7454), .I2(n7455), .O(n7463));
  LUT3 #(.INIT(8'hE8)) lut_n7464 (.I0(n7459), .I1(n7462), .I2(n7463), .O(n7464));
  LUT3 #(.INIT(8'h96)) lut_n7465 (.I0(n7438), .I1(n7446), .I2(n7447), .O(n7465));
  LUT3 #(.INIT(8'hE8)) lut_n7466 (.I0(n7456), .I1(n7464), .I2(n7465), .O(n7466));
  LUT3 #(.INIT(8'h96)) lut_n7467 (.I0(n7410), .I1(n7428), .I2(n7429), .O(n7467));
  LUT3 #(.INIT(8'hE8)) lut_n7468 (.I0(n7448), .I1(n7466), .I2(n7467), .O(n7468));
  LUT3 #(.INIT(8'h96)) lut_n7469 (.I0(n7350), .I1(n7388), .I2(n7389), .O(n7469));
  LUT3 #(.INIT(8'hE8)) lut_n7470 (.I0(n7430), .I1(n7468), .I2(n7469), .O(n7470));
  LUT3 #(.INIT(8'hE8)) lut_n7471 (.I0(x2976), .I1(x2977), .I2(x2978), .O(n7471));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7472 (.I0(x2967), .I1(x2968), .I2(x2969), .I3(n7460), .I4(n7461), .O(n7472));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7473 (.I0(x2973), .I1(x2974), .I2(x2975), .I3(n7471), .I4(n7472), .O(n7473));
  LUT3 #(.INIT(8'hE8)) lut_n7474 (.I0(x2982), .I1(x2983), .I2(x2984), .O(n7474));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7475 (.I0(x2973), .I1(x2974), .I2(x2975), .I3(n7471), .I4(n7472), .O(n7475));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7476 (.I0(x2979), .I1(x2980), .I2(x2981), .I3(n7474), .I4(n7475), .O(n7476));
  LUT3 #(.INIT(8'h96)) lut_n7477 (.I0(n7459), .I1(n7462), .I2(n7463), .O(n7477));
  LUT3 #(.INIT(8'hE8)) lut_n7478 (.I0(n7473), .I1(n7476), .I2(n7477), .O(n7478));
  LUT3 #(.INIT(8'hE8)) lut_n7479 (.I0(x2988), .I1(x2989), .I2(x2990), .O(n7479));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7480 (.I0(x2979), .I1(x2980), .I2(x2981), .I3(n7474), .I4(n7475), .O(n7480));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7481 (.I0(x2985), .I1(x2986), .I2(x2987), .I3(n7479), .I4(n7480), .O(n7481));
  LUT3 #(.INIT(8'hE8)) lut_n7482 (.I0(x2994), .I1(x2995), .I2(x2996), .O(n7482));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7483 (.I0(x2985), .I1(x2986), .I2(x2987), .I3(n7479), .I4(n7480), .O(n7483));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7484 (.I0(x2991), .I1(x2992), .I2(x2993), .I3(n7482), .I4(n7483), .O(n7484));
  LUT3 #(.INIT(8'h96)) lut_n7485 (.I0(n7473), .I1(n7476), .I2(n7477), .O(n7485));
  LUT3 #(.INIT(8'hE8)) lut_n7486 (.I0(n7481), .I1(n7484), .I2(n7485), .O(n7486));
  LUT3 #(.INIT(8'h96)) lut_n7487 (.I0(n7456), .I1(n7464), .I2(n7465), .O(n7487));
  LUT3 #(.INIT(8'hE8)) lut_n7488 (.I0(n7478), .I1(n7486), .I2(n7487), .O(n7488));
  LUT3 #(.INIT(8'hE8)) lut_n7489 (.I0(x2997), .I1(x2998), .I2(x2999), .O(n7489));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7490 (.I0(x2991), .I1(x2992), .I2(x2993), .I3(n7482), .I4(n7483), .O(n7490));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7491 (.I0(x3000), .I1(x3001), .I2(x3002), .I3(n7489), .I4(n7490), .O(n7491));
  LUT3 #(.INIT(8'hE8)) lut_n7492 (.I0(x3006), .I1(x3007), .I2(x3008), .O(n7492));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7493 (.I0(x3000), .I1(x3001), .I2(x3002), .I3(n7489), .I4(n7490), .O(n7493));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7494 (.I0(x3003), .I1(x3004), .I2(x3005), .I3(n7492), .I4(n7493), .O(n7494));
  LUT3 #(.INIT(8'h96)) lut_n7495 (.I0(n7481), .I1(n7484), .I2(n7485), .O(n7495));
  LUT3 #(.INIT(8'hE8)) lut_n7496 (.I0(n7491), .I1(n7494), .I2(n7495), .O(n7496));
  LUT3 #(.INIT(8'hE8)) lut_n7497 (.I0(x3012), .I1(x3013), .I2(x3014), .O(n7497));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7498 (.I0(x3003), .I1(x3004), .I2(x3005), .I3(n7492), .I4(n7493), .O(n7498));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7499 (.I0(x3009), .I1(x3010), .I2(x3011), .I3(n7497), .I4(n7498), .O(n7499));
  LUT3 #(.INIT(8'hE8)) lut_n7500 (.I0(x3018), .I1(x3019), .I2(x3020), .O(n7500));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7501 (.I0(x3009), .I1(x3010), .I2(x3011), .I3(n7497), .I4(n7498), .O(n7501));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7502 (.I0(x3015), .I1(x3016), .I2(x3017), .I3(n7500), .I4(n7501), .O(n7502));
  LUT3 #(.INIT(8'h96)) lut_n7503 (.I0(n7491), .I1(n7494), .I2(n7495), .O(n7503));
  LUT3 #(.INIT(8'hE8)) lut_n7504 (.I0(n7499), .I1(n7502), .I2(n7503), .O(n7504));
  LUT3 #(.INIT(8'h96)) lut_n7505 (.I0(n7478), .I1(n7486), .I2(n7487), .O(n7505));
  LUT3 #(.INIT(8'hE8)) lut_n7506 (.I0(n7496), .I1(n7504), .I2(n7505), .O(n7506));
  LUT3 #(.INIT(8'h96)) lut_n7507 (.I0(n7448), .I1(n7466), .I2(n7467), .O(n7507));
  LUT3 #(.INIT(8'hE8)) lut_n7508 (.I0(n7488), .I1(n7506), .I2(n7507), .O(n7508));
  LUT3 #(.INIT(8'hE8)) lut_n7509 (.I0(x3024), .I1(x3025), .I2(x3026), .O(n7509));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7510 (.I0(x3015), .I1(x3016), .I2(x3017), .I3(n7500), .I4(n7501), .O(n7510));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7511 (.I0(x3021), .I1(x3022), .I2(x3023), .I3(n7509), .I4(n7510), .O(n7511));
  LUT3 #(.INIT(8'hE8)) lut_n7512 (.I0(x3030), .I1(x3031), .I2(x3032), .O(n7512));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7513 (.I0(x3021), .I1(x3022), .I2(x3023), .I3(n7509), .I4(n7510), .O(n7513));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7514 (.I0(x3027), .I1(x3028), .I2(x3029), .I3(n7512), .I4(n7513), .O(n7514));
  LUT3 #(.INIT(8'h96)) lut_n7515 (.I0(n7499), .I1(n7502), .I2(n7503), .O(n7515));
  LUT3 #(.INIT(8'hE8)) lut_n7516 (.I0(n7511), .I1(n7514), .I2(n7515), .O(n7516));
  LUT3 #(.INIT(8'hE8)) lut_n7517 (.I0(x3036), .I1(x3037), .I2(x3038), .O(n7517));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7518 (.I0(x3027), .I1(x3028), .I2(x3029), .I3(n7512), .I4(n7513), .O(n7518));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7519 (.I0(x3033), .I1(x3034), .I2(x3035), .I3(n7517), .I4(n7518), .O(n7519));
  LUT3 #(.INIT(8'hE8)) lut_n7520 (.I0(x3042), .I1(x3043), .I2(x3044), .O(n7520));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7521 (.I0(x3033), .I1(x3034), .I2(x3035), .I3(n7517), .I4(n7518), .O(n7521));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7522 (.I0(x3039), .I1(x3040), .I2(x3041), .I3(n7520), .I4(n7521), .O(n7522));
  LUT3 #(.INIT(8'h96)) lut_n7523 (.I0(n7511), .I1(n7514), .I2(n7515), .O(n7523));
  LUT3 #(.INIT(8'hE8)) lut_n7524 (.I0(n7519), .I1(n7522), .I2(n7523), .O(n7524));
  LUT3 #(.INIT(8'h96)) lut_n7525 (.I0(n7496), .I1(n7504), .I2(n7505), .O(n7525));
  LUT3 #(.INIT(8'hE8)) lut_n7526 (.I0(n7516), .I1(n7524), .I2(n7525), .O(n7526));
  LUT3 #(.INIT(8'hE8)) lut_n7527 (.I0(x3048), .I1(x3049), .I2(x3050), .O(n7527));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7528 (.I0(x3039), .I1(x3040), .I2(x3041), .I3(n7520), .I4(n7521), .O(n7528));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7529 (.I0(x3045), .I1(x3046), .I2(x3047), .I3(n7527), .I4(n7528), .O(n7529));
  LUT3 #(.INIT(8'hE8)) lut_n7530 (.I0(x3054), .I1(x3055), .I2(x3056), .O(n7530));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7531 (.I0(x3045), .I1(x3046), .I2(x3047), .I3(n7527), .I4(n7528), .O(n7531));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7532 (.I0(x3051), .I1(x3052), .I2(x3053), .I3(n7530), .I4(n7531), .O(n7532));
  LUT3 #(.INIT(8'h96)) lut_n7533 (.I0(n7519), .I1(n7522), .I2(n7523), .O(n7533));
  LUT3 #(.INIT(8'hE8)) lut_n7534 (.I0(n7529), .I1(n7532), .I2(n7533), .O(n7534));
  LUT3 #(.INIT(8'hE8)) lut_n7535 (.I0(x3060), .I1(x3061), .I2(x3062), .O(n7535));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7536 (.I0(x3051), .I1(x3052), .I2(x3053), .I3(n7530), .I4(n7531), .O(n7536));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7537 (.I0(x3057), .I1(x3058), .I2(x3059), .I3(n7535), .I4(n7536), .O(n7537));
  LUT3 #(.INIT(8'hE8)) lut_n7538 (.I0(x3066), .I1(x3067), .I2(x3068), .O(n7538));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7539 (.I0(x3057), .I1(x3058), .I2(x3059), .I3(n7535), .I4(n7536), .O(n7539));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7540 (.I0(x3063), .I1(x3064), .I2(x3065), .I3(n7538), .I4(n7539), .O(n7540));
  LUT3 #(.INIT(8'h96)) lut_n7541 (.I0(n7529), .I1(n7532), .I2(n7533), .O(n7541));
  LUT3 #(.INIT(8'hE8)) lut_n7542 (.I0(n7537), .I1(n7540), .I2(n7541), .O(n7542));
  LUT3 #(.INIT(8'h96)) lut_n7543 (.I0(n7516), .I1(n7524), .I2(n7525), .O(n7543));
  LUT3 #(.INIT(8'hE8)) lut_n7544 (.I0(n7534), .I1(n7542), .I2(n7543), .O(n7544));
  LUT3 #(.INIT(8'h96)) lut_n7545 (.I0(n7488), .I1(n7506), .I2(n7507), .O(n7545));
  LUT3 #(.INIT(8'hE8)) lut_n7546 (.I0(n7526), .I1(n7544), .I2(n7545), .O(n7546));
  LUT3 #(.INIT(8'h96)) lut_n7547 (.I0(n7430), .I1(n7468), .I2(n7469), .O(n7547));
  LUT3 #(.INIT(8'hE8)) lut_n7548 (.I0(n7508), .I1(n7546), .I2(n7547), .O(n7548));
  LUT3 #(.INIT(8'h96)) lut_n7549 (.I0(n7312), .I1(n7390), .I2(n7391), .O(n7549));
  LUT3 #(.INIT(8'hE8)) lut_n7550 (.I0(n7470), .I1(n7548), .I2(n7549), .O(n7550));
  LUT3 #(.INIT(8'h96)) lut_n7551 (.I0(n7074), .I1(n7232), .I2(n7233), .O(n7551));
  LUT3 #(.INIT(8'hE8)) lut_n7552 (.I0(n7392), .I1(n7550), .I2(n7551), .O(n7552));
  LUT3 #(.INIT(8'h96)) lut_n7553 (.I0(n6596), .I1(n6914), .I2(n6915), .O(n7553));
  LUT3 #(.INIT(8'hE8)) lut_n7554 (.I0(n7234), .I1(n7552), .I2(n7553), .O(n7554));
  LUT3 #(.INIT(8'hE8)) lut_n7555 (.I0(n6278), .I1(n6916), .I2(n7554), .O(n7555));
  LUT3 #(.INIT(8'hE8)) lut_n7556 (.I0(x3072), .I1(x3073), .I2(x3074), .O(n7556));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7557 (.I0(x3063), .I1(x3064), .I2(x3065), .I3(n7538), .I4(n7539), .O(n7557));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7558 (.I0(x3069), .I1(x3070), .I2(x3071), .I3(n7556), .I4(n7557), .O(n7558));
  LUT3 #(.INIT(8'hE8)) lut_n7559 (.I0(x3078), .I1(x3079), .I2(x3080), .O(n7559));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7560 (.I0(x3069), .I1(x3070), .I2(x3071), .I3(n7556), .I4(n7557), .O(n7560));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7561 (.I0(x3075), .I1(x3076), .I2(x3077), .I3(n7559), .I4(n7560), .O(n7561));
  LUT3 #(.INIT(8'h96)) lut_n7562 (.I0(n7537), .I1(n7540), .I2(n7541), .O(n7562));
  LUT3 #(.INIT(8'hE8)) lut_n7563 (.I0(n7558), .I1(n7561), .I2(n7562), .O(n7563));
  LUT3 #(.INIT(8'hE8)) lut_n7564 (.I0(x3084), .I1(x3085), .I2(x3086), .O(n7564));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7565 (.I0(x3075), .I1(x3076), .I2(x3077), .I3(n7559), .I4(n7560), .O(n7565));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7566 (.I0(x3081), .I1(x3082), .I2(x3083), .I3(n7564), .I4(n7565), .O(n7566));
  LUT3 #(.INIT(8'hE8)) lut_n7567 (.I0(x3090), .I1(x3091), .I2(x3092), .O(n7567));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7568 (.I0(x3081), .I1(x3082), .I2(x3083), .I3(n7564), .I4(n7565), .O(n7568));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7569 (.I0(x3087), .I1(x3088), .I2(x3089), .I3(n7567), .I4(n7568), .O(n7569));
  LUT3 #(.INIT(8'h96)) lut_n7570 (.I0(n7558), .I1(n7561), .I2(n7562), .O(n7570));
  LUT3 #(.INIT(8'hE8)) lut_n7571 (.I0(n7566), .I1(n7569), .I2(n7570), .O(n7571));
  LUT3 #(.INIT(8'h96)) lut_n7572 (.I0(n7534), .I1(n7542), .I2(n7543), .O(n7572));
  LUT3 #(.INIT(8'hE8)) lut_n7573 (.I0(n7563), .I1(n7571), .I2(n7572), .O(n7573));
  LUT3 #(.INIT(8'hE8)) lut_n7574 (.I0(x3096), .I1(x3097), .I2(x3098), .O(n7574));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7575 (.I0(x3087), .I1(x3088), .I2(x3089), .I3(n7567), .I4(n7568), .O(n7575));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7576 (.I0(x3093), .I1(x3094), .I2(x3095), .I3(n7574), .I4(n7575), .O(n7576));
  LUT3 #(.INIT(8'hE8)) lut_n7577 (.I0(x3102), .I1(x3103), .I2(x3104), .O(n7577));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7578 (.I0(x3093), .I1(x3094), .I2(x3095), .I3(n7574), .I4(n7575), .O(n7578));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7579 (.I0(x3099), .I1(x3100), .I2(x3101), .I3(n7577), .I4(n7578), .O(n7579));
  LUT3 #(.INIT(8'h96)) lut_n7580 (.I0(n7566), .I1(n7569), .I2(n7570), .O(n7580));
  LUT3 #(.INIT(8'hE8)) lut_n7581 (.I0(n7576), .I1(n7579), .I2(n7580), .O(n7581));
  LUT3 #(.INIT(8'hE8)) lut_n7582 (.I0(x3108), .I1(x3109), .I2(x3110), .O(n7582));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7583 (.I0(x3099), .I1(x3100), .I2(x3101), .I3(n7577), .I4(n7578), .O(n7583));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7584 (.I0(x3105), .I1(x3106), .I2(x3107), .I3(n7582), .I4(n7583), .O(n7584));
  LUT3 #(.INIT(8'hE8)) lut_n7585 (.I0(x3114), .I1(x3115), .I2(x3116), .O(n7585));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7586 (.I0(x3105), .I1(x3106), .I2(x3107), .I3(n7582), .I4(n7583), .O(n7586));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7587 (.I0(x3111), .I1(x3112), .I2(x3113), .I3(n7585), .I4(n7586), .O(n7587));
  LUT3 #(.INIT(8'h96)) lut_n7588 (.I0(n7576), .I1(n7579), .I2(n7580), .O(n7588));
  LUT3 #(.INIT(8'hE8)) lut_n7589 (.I0(n7584), .I1(n7587), .I2(n7588), .O(n7589));
  LUT3 #(.INIT(8'h96)) lut_n7590 (.I0(n7563), .I1(n7571), .I2(n7572), .O(n7590));
  LUT3 #(.INIT(8'hE8)) lut_n7591 (.I0(n7581), .I1(n7589), .I2(n7590), .O(n7591));
  LUT3 #(.INIT(8'h96)) lut_n7592 (.I0(n7526), .I1(n7544), .I2(n7545), .O(n7592));
  LUT3 #(.INIT(8'hE8)) lut_n7593 (.I0(n7573), .I1(n7591), .I2(n7592), .O(n7593));
  LUT3 #(.INIT(8'hE8)) lut_n7594 (.I0(x3120), .I1(x3121), .I2(x3122), .O(n7594));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7595 (.I0(x3111), .I1(x3112), .I2(x3113), .I3(n7585), .I4(n7586), .O(n7595));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7596 (.I0(x3117), .I1(x3118), .I2(x3119), .I3(n7594), .I4(n7595), .O(n7596));
  LUT3 #(.INIT(8'hE8)) lut_n7597 (.I0(x3126), .I1(x3127), .I2(x3128), .O(n7597));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7598 (.I0(x3117), .I1(x3118), .I2(x3119), .I3(n7594), .I4(n7595), .O(n7598));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7599 (.I0(x3123), .I1(x3124), .I2(x3125), .I3(n7597), .I4(n7598), .O(n7599));
  LUT3 #(.INIT(8'h96)) lut_n7600 (.I0(n7584), .I1(n7587), .I2(n7588), .O(n7600));
  LUT3 #(.INIT(8'hE8)) lut_n7601 (.I0(n7596), .I1(n7599), .I2(n7600), .O(n7601));
  LUT3 #(.INIT(8'hE8)) lut_n7602 (.I0(x3132), .I1(x3133), .I2(x3134), .O(n7602));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7603 (.I0(x3123), .I1(x3124), .I2(x3125), .I3(n7597), .I4(n7598), .O(n7603));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7604 (.I0(x3129), .I1(x3130), .I2(x3131), .I3(n7602), .I4(n7603), .O(n7604));
  LUT3 #(.INIT(8'hE8)) lut_n7605 (.I0(x3138), .I1(x3139), .I2(x3140), .O(n7605));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7606 (.I0(x3129), .I1(x3130), .I2(x3131), .I3(n7602), .I4(n7603), .O(n7606));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7607 (.I0(x3135), .I1(x3136), .I2(x3137), .I3(n7605), .I4(n7606), .O(n7607));
  LUT3 #(.INIT(8'h96)) lut_n7608 (.I0(n7596), .I1(n7599), .I2(n7600), .O(n7608));
  LUT3 #(.INIT(8'hE8)) lut_n7609 (.I0(n7604), .I1(n7607), .I2(n7608), .O(n7609));
  LUT3 #(.INIT(8'h96)) lut_n7610 (.I0(n7581), .I1(n7589), .I2(n7590), .O(n7610));
  LUT3 #(.INIT(8'hE8)) lut_n7611 (.I0(n7601), .I1(n7609), .I2(n7610), .O(n7611));
  LUT3 #(.INIT(8'hE8)) lut_n7612 (.I0(x3144), .I1(x3145), .I2(x3146), .O(n7612));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7613 (.I0(x3135), .I1(x3136), .I2(x3137), .I3(n7605), .I4(n7606), .O(n7613));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7614 (.I0(x3141), .I1(x3142), .I2(x3143), .I3(n7612), .I4(n7613), .O(n7614));
  LUT3 #(.INIT(8'hE8)) lut_n7615 (.I0(x3150), .I1(x3151), .I2(x3152), .O(n7615));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7616 (.I0(x3141), .I1(x3142), .I2(x3143), .I3(n7612), .I4(n7613), .O(n7616));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7617 (.I0(x3147), .I1(x3148), .I2(x3149), .I3(n7615), .I4(n7616), .O(n7617));
  LUT3 #(.INIT(8'h96)) lut_n7618 (.I0(n7604), .I1(n7607), .I2(n7608), .O(n7618));
  LUT3 #(.INIT(8'hE8)) lut_n7619 (.I0(n7614), .I1(n7617), .I2(n7618), .O(n7619));
  LUT3 #(.INIT(8'hE8)) lut_n7620 (.I0(x3156), .I1(x3157), .I2(x3158), .O(n7620));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7621 (.I0(x3147), .I1(x3148), .I2(x3149), .I3(n7615), .I4(n7616), .O(n7621));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7622 (.I0(x3153), .I1(x3154), .I2(x3155), .I3(n7620), .I4(n7621), .O(n7622));
  LUT3 #(.INIT(8'hE8)) lut_n7623 (.I0(x3162), .I1(x3163), .I2(x3164), .O(n7623));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7624 (.I0(x3153), .I1(x3154), .I2(x3155), .I3(n7620), .I4(n7621), .O(n7624));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7625 (.I0(x3159), .I1(x3160), .I2(x3161), .I3(n7623), .I4(n7624), .O(n7625));
  LUT3 #(.INIT(8'h96)) lut_n7626 (.I0(n7614), .I1(n7617), .I2(n7618), .O(n7626));
  LUT3 #(.INIT(8'hE8)) lut_n7627 (.I0(n7622), .I1(n7625), .I2(n7626), .O(n7627));
  LUT3 #(.INIT(8'h96)) lut_n7628 (.I0(n7601), .I1(n7609), .I2(n7610), .O(n7628));
  LUT3 #(.INIT(8'hE8)) lut_n7629 (.I0(n7619), .I1(n7627), .I2(n7628), .O(n7629));
  LUT3 #(.INIT(8'h96)) lut_n7630 (.I0(n7573), .I1(n7591), .I2(n7592), .O(n7630));
  LUT3 #(.INIT(8'hE8)) lut_n7631 (.I0(n7611), .I1(n7629), .I2(n7630), .O(n7631));
  LUT3 #(.INIT(8'h96)) lut_n7632 (.I0(n7508), .I1(n7546), .I2(n7547), .O(n7632));
  LUT3 #(.INIT(8'hE8)) lut_n7633 (.I0(n7593), .I1(n7631), .I2(n7632), .O(n7633));
  LUT3 #(.INIT(8'hE8)) lut_n7634 (.I0(x3168), .I1(x3169), .I2(x3170), .O(n7634));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7635 (.I0(x3159), .I1(x3160), .I2(x3161), .I3(n7623), .I4(n7624), .O(n7635));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7636 (.I0(x3165), .I1(x3166), .I2(x3167), .I3(n7634), .I4(n7635), .O(n7636));
  LUT3 #(.INIT(8'hE8)) lut_n7637 (.I0(x3174), .I1(x3175), .I2(x3176), .O(n7637));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7638 (.I0(x3165), .I1(x3166), .I2(x3167), .I3(n7634), .I4(n7635), .O(n7638));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7639 (.I0(x3171), .I1(x3172), .I2(x3173), .I3(n7637), .I4(n7638), .O(n7639));
  LUT3 #(.INIT(8'h96)) lut_n7640 (.I0(n7622), .I1(n7625), .I2(n7626), .O(n7640));
  LUT3 #(.INIT(8'hE8)) lut_n7641 (.I0(n7636), .I1(n7639), .I2(n7640), .O(n7641));
  LUT3 #(.INIT(8'hE8)) lut_n7642 (.I0(x3180), .I1(x3181), .I2(x3182), .O(n7642));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7643 (.I0(x3171), .I1(x3172), .I2(x3173), .I3(n7637), .I4(n7638), .O(n7643));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7644 (.I0(x3177), .I1(x3178), .I2(x3179), .I3(n7642), .I4(n7643), .O(n7644));
  LUT3 #(.INIT(8'hE8)) lut_n7645 (.I0(x3186), .I1(x3187), .I2(x3188), .O(n7645));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7646 (.I0(x3177), .I1(x3178), .I2(x3179), .I3(n7642), .I4(n7643), .O(n7646));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7647 (.I0(x3183), .I1(x3184), .I2(x3185), .I3(n7645), .I4(n7646), .O(n7647));
  LUT3 #(.INIT(8'h96)) lut_n7648 (.I0(n7636), .I1(n7639), .I2(n7640), .O(n7648));
  LUT3 #(.INIT(8'hE8)) lut_n7649 (.I0(n7644), .I1(n7647), .I2(n7648), .O(n7649));
  LUT3 #(.INIT(8'h96)) lut_n7650 (.I0(n7619), .I1(n7627), .I2(n7628), .O(n7650));
  LUT3 #(.INIT(8'hE8)) lut_n7651 (.I0(n7641), .I1(n7649), .I2(n7650), .O(n7651));
  LUT3 #(.INIT(8'hE8)) lut_n7652 (.I0(x3192), .I1(x3193), .I2(x3194), .O(n7652));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7653 (.I0(x3183), .I1(x3184), .I2(x3185), .I3(n7645), .I4(n7646), .O(n7653));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7654 (.I0(x3189), .I1(x3190), .I2(x3191), .I3(n7652), .I4(n7653), .O(n7654));
  LUT3 #(.INIT(8'hE8)) lut_n7655 (.I0(x3198), .I1(x3199), .I2(x3200), .O(n7655));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7656 (.I0(x3189), .I1(x3190), .I2(x3191), .I3(n7652), .I4(n7653), .O(n7656));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7657 (.I0(x3195), .I1(x3196), .I2(x3197), .I3(n7655), .I4(n7656), .O(n7657));
  LUT3 #(.INIT(8'h96)) lut_n7658 (.I0(n7644), .I1(n7647), .I2(n7648), .O(n7658));
  LUT3 #(.INIT(8'hE8)) lut_n7659 (.I0(n7654), .I1(n7657), .I2(n7658), .O(n7659));
  LUT3 #(.INIT(8'hE8)) lut_n7660 (.I0(x3204), .I1(x3205), .I2(x3206), .O(n7660));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7661 (.I0(x3195), .I1(x3196), .I2(x3197), .I3(n7655), .I4(n7656), .O(n7661));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7662 (.I0(x3201), .I1(x3202), .I2(x3203), .I3(n7660), .I4(n7661), .O(n7662));
  LUT3 #(.INIT(8'hE8)) lut_n7663 (.I0(x3210), .I1(x3211), .I2(x3212), .O(n7663));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7664 (.I0(x3201), .I1(x3202), .I2(x3203), .I3(n7660), .I4(n7661), .O(n7664));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7665 (.I0(x3207), .I1(x3208), .I2(x3209), .I3(n7663), .I4(n7664), .O(n7665));
  LUT3 #(.INIT(8'h96)) lut_n7666 (.I0(n7654), .I1(n7657), .I2(n7658), .O(n7666));
  LUT3 #(.INIT(8'hE8)) lut_n7667 (.I0(n7662), .I1(n7665), .I2(n7666), .O(n7667));
  LUT3 #(.INIT(8'h96)) lut_n7668 (.I0(n7641), .I1(n7649), .I2(n7650), .O(n7668));
  LUT3 #(.INIT(8'hE8)) lut_n7669 (.I0(n7659), .I1(n7667), .I2(n7668), .O(n7669));
  LUT3 #(.INIT(8'h96)) lut_n7670 (.I0(n7611), .I1(n7629), .I2(n7630), .O(n7670));
  LUT3 #(.INIT(8'hE8)) lut_n7671 (.I0(n7651), .I1(n7669), .I2(n7670), .O(n7671));
  LUT3 #(.INIT(8'hE8)) lut_n7672 (.I0(x3216), .I1(x3217), .I2(x3218), .O(n7672));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7673 (.I0(x3207), .I1(x3208), .I2(x3209), .I3(n7663), .I4(n7664), .O(n7673));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7674 (.I0(x3213), .I1(x3214), .I2(x3215), .I3(n7672), .I4(n7673), .O(n7674));
  LUT3 #(.INIT(8'hE8)) lut_n7675 (.I0(x3222), .I1(x3223), .I2(x3224), .O(n7675));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7676 (.I0(x3213), .I1(x3214), .I2(x3215), .I3(n7672), .I4(n7673), .O(n7676));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7677 (.I0(x3219), .I1(x3220), .I2(x3221), .I3(n7675), .I4(n7676), .O(n7677));
  LUT3 #(.INIT(8'h96)) lut_n7678 (.I0(n7662), .I1(n7665), .I2(n7666), .O(n7678));
  LUT3 #(.INIT(8'hE8)) lut_n7679 (.I0(n7674), .I1(n7677), .I2(n7678), .O(n7679));
  LUT3 #(.INIT(8'hE8)) lut_n7680 (.I0(x3228), .I1(x3229), .I2(x3230), .O(n7680));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7681 (.I0(x3219), .I1(x3220), .I2(x3221), .I3(n7675), .I4(n7676), .O(n7681));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7682 (.I0(x3225), .I1(x3226), .I2(x3227), .I3(n7680), .I4(n7681), .O(n7682));
  LUT3 #(.INIT(8'hE8)) lut_n7683 (.I0(x3234), .I1(x3235), .I2(x3236), .O(n7683));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7684 (.I0(x3225), .I1(x3226), .I2(x3227), .I3(n7680), .I4(n7681), .O(n7684));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7685 (.I0(x3231), .I1(x3232), .I2(x3233), .I3(n7683), .I4(n7684), .O(n7685));
  LUT3 #(.INIT(8'h96)) lut_n7686 (.I0(n7674), .I1(n7677), .I2(n7678), .O(n7686));
  LUT3 #(.INIT(8'hE8)) lut_n7687 (.I0(n7682), .I1(n7685), .I2(n7686), .O(n7687));
  LUT3 #(.INIT(8'h96)) lut_n7688 (.I0(n7659), .I1(n7667), .I2(n7668), .O(n7688));
  LUT3 #(.INIT(8'hE8)) lut_n7689 (.I0(n7679), .I1(n7687), .I2(n7688), .O(n7689));
  LUT3 #(.INIT(8'hE8)) lut_n7690 (.I0(x3240), .I1(x3241), .I2(x3242), .O(n7690));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7691 (.I0(x3231), .I1(x3232), .I2(x3233), .I3(n7683), .I4(n7684), .O(n7691));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7692 (.I0(x3237), .I1(x3238), .I2(x3239), .I3(n7690), .I4(n7691), .O(n7692));
  LUT3 #(.INIT(8'hE8)) lut_n7693 (.I0(x3246), .I1(x3247), .I2(x3248), .O(n7693));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7694 (.I0(x3237), .I1(x3238), .I2(x3239), .I3(n7690), .I4(n7691), .O(n7694));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7695 (.I0(x3243), .I1(x3244), .I2(x3245), .I3(n7693), .I4(n7694), .O(n7695));
  LUT3 #(.INIT(8'h96)) lut_n7696 (.I0(n7682), .I1(n7685), .I2(n7686), .O(n7696));
  LUT3 #(.INIT(8'hE8)) lut_n7697 (.I0(n7692), .I1(n7695), .I2(n7696), .O(n7697));
  LUT3 #(.INIT(8'hE8)) lut_n7698 (.I0(x3252), .I1(x3253), .I2(x3254), .O(n7698));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7699 (.I0(x3243), .I1(x3244), .I2(x3245), .I3(n7693), .I4(n7694), .O(n7699));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7700 (.I0(x3249), .I1(x3250), .I2(x3251), .I3(n7698), .I4(n7699), .O(n7700));
  LUT3 #(.INIT(8'hE8)) lut_n7701 (.I0(x3258), .I1(x3259), .I2(x3260), .O(n7701));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7702 (.I0(x3249), .I1(x3250), .I2(x3251), .I3(n7698), .I4(n7699), .O(n7702));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7703 (.I0(x3255), .I1(x3256), .I2(x3257), .I3(n7701), .I4(n7702), .O(n7703));
  LUT3 #(.INIT(8'h96)) lut_n7704 (.I0(n7692), .I1(n7695), .I2(n7696), .O(n7704));
  LUT3 #(.INIT(8'hE8)) lut_n7705 (.I0(n7700), .I1(n7703), .I2(n7704), .O(n7705));
  LUT3 #(.INIT(8'h96)) lut_n7706 (.I0(n7679), .I1(n7687), .I2(n7688), .O(n7706));
  LUT3 #(.INIT(8'hE8)) lut_n7707 (.I0(n7697), .I1(n7705), .I2(n7706), .O(n7707));
  LUT3 #(.INIT(8'h96)) lut_n7708 (.I0(n7651), .I1(n7669), .I2(n7670), .O(n7708));
  LUT3 #(.INIT(8'hE8)) lut_n7709 (.I0(n7689), .I1(n7707), .I2(n7708), .O(n7709));
  LUT3 #(.INIT(8'h96)) lut_n7710 (.I0(n7593), .I1(n7631), .I2(n7632), .O(n7710));
  LUT3 #(.INIT(8'hE8)) lut_n7711 (.I0(n7671), .I1(n7709), .I2(n7710), .O(n7711));
  LUT3 #(.INIT(8'h96)) lut_n7712 (.I0(n7470), .I1(n7548), .I2(n7549), .O(n7712));
  LUT3 #(.INIT(8'hE8)) lut_n7713 (.I0(n7633), .I1(n7711), .I2(n7712), .O(n7713));
  LUT3 #(.INIT(8'hE8)) lut_n7714 (.I0(x3264), .I1(x3265), .I2(x3266), .O(n7714));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7715 (.I0(x3255), .I1(x3256), .I2(x3257), .I3(n7701), .I4(n7702), .O(n7715));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7716 (.I0(x3261), .I1(x3262), .I2(x3263), .I3(n7714), .I4(n7715), .O(n7716));
  LUT3 #(.INIT(8'hE8)) lut_n7717 (.I0(x3270), .I1(x3271), .I2(x3272), .O(n7717));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7718 (.I0(x3261), .I1(x3262), .I2(x3263), .I3(n7714), .I4(n7715), .O(n7718));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7719 (.I0(x3267), .I1(x3268), .I2(x3269), .I3(n7717), .I4(n7718), .O(n7719));
  LUT3 #(.INIT(8'h96)) lut_n7720 (.I0(n7700), .I1(n7703), .I2(n7704), .O(n7720));
  LUT3 #(.INIT(8'hE8)) lut_n7721 (.I0(n7716), .I1(n7719), .I2(n7720), .O(n7721));
  LUT3 #(.INIT(8'hE8)) lut_n7722 (.I0(x3276), .I1(x3277), .I2(x3278), .O(n7722));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7723 (.I0(x3267), .I1(x3268), .I2(x3269), .I3(n7717), .I4(n7718), .O(n7723));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7724 (.I0(x3273), .I1(x3274), .I2(x3275), .I3(n7722), .I4(n7723), .O(n7724));
  LUT3 #(.INIT(8'hE8)) lut_n7725 (.I0(x3282), .I1(x3283), .I2(x3284), .O(n7725));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7726 (.I0(x3273), .I1(x3274), .I2(x3275), .I3(n7722), .I4(n7723), .O(n7726));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7727 (.I0(x3279), .I1(x3280), .I2(x3281), .I3(n7725), .I4(n7726), .O(n7727));
  LUT3 #(.INIT(8'h96)) lut_n7728 (.I0(n7716), .I1(n7719), .I2(n7720), .O(n7728));
  LUT3 #(.INIT(8'hE8)) lut_n7729 (.I0(n7724), .I1(n7727), .I2(n7728), .O(n7729));
  LUT3 #(.INIT(8'h96)) lut_n7730 (.I0(n7697), .I1(n7705), .I2(n7706), .O(n7730));
  LUT3 #(.INIT(8'hE8)) lut_n7731 (.I0(n7721), .I1(n7729), .I2(n7730), .O(n7731));
  LUT3 #(.INIT(8'hE8)) lut_n7732 (.I0(x3288), .I1(x3289), .I2(x3290), .O(n7732));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7733 (.I0(x3279), .I1(x3280), .I2(x3281), .I3(n7725), .I4(n7726), .O(n7733));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7734 (.I0(x3285), .I1(x3286), .I2(x3287), .I3(n7732), .I4(n7733), .O(n7734));
  LUT3 #(.INIT(8'hE8)) lut_n7735 (.I0(x3294), .I1(x3295), .I2(x3296), .O(n7735));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7736 (.I0(x3285), .I1(x3286), .I2(x3287), .I3(n7732), .I4(n7733), .O(n7736));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7737 (.I0(x3291), .I1(x3292), .I2(x3293), .I3(n7735), .I4(n7736), .O(n7737));
  LUT3 #(.INIT(8'h96)) lut_n7738 (.I0(n7724), .I1(n7727), .I2(n7728), .O(n7738));
  LUT3 #(.INIT(8'hE8)) lut_n7739 (.I0(n7734), .I1(n7737), .I2(n7738), .O(n7739));
  LUT3 #(.INIT(8'hE8)) lut_n7740 (.I0(x3300), .I1(x3301), .I2(x3302), .O(n7740));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7741 (.I0(x3291), .I1(x3292), .I2(x3293), .I3(n7735), .I4(n7736), .O(n7741));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7742 (.I0(x3297), .I1(x3298), .I2(x3299), .I3(n7740), .I4(n7741), .O(n7742));
  LUT3 #(.INIT(8'hE8)) lut_n7743 (.I0(x3306), .I1(x3307), .I2(x3308), .O(n7743));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7744 (.I0(x3297), .I1(x3298), .I2(x3299), .I3(n7740), .I4(n7741), .O(n7744));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7745 (.I0(x3303), .I1(x3304), .I2(x3305), .I3(n7743), .I4(n7744), .O(n7745));
  LUT3 #(.INIT(8'h96)) lut_n7746 (.I0(n7734), .I1(n7737), .I2(n7738), .O(n7746));
  LUT3 #(.INIT(8'hE8)) lut_n7747 (.I0(n7742), .I1(n7745), .I2(n7746), .O(n7747));
  LUT3 #(.INIT(8'h96)) lut_n7748 (.I0(n7721), .I1(n7729), .I2(n7730), .O(n7748));
  LUT3 #(.INIT(8'hE8)) lut_n7749 (.I0(n7739), .I1(n7747), .I2(n7748), .O(n7749));
  LUT3 #(.INIT(8'h96)) lut_n7750 (.I0(n7689), .I1(n7707), .I2(n7708), .O(n7750));
  LUT3 #(.INIT(8'hE8)) lut_n7751 (.I0(n7731), .I1(n7749), .I2(n7750), .O(n7751));
  LUT3 #(.INIT(8'hE8)) lut_n7752 (.I0(x3312), .I1(x3313), .I2(x3314), .O(n7752));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7753 (.I0(x3303), .I1(x3304), .I2(x3305), .I3(n7743), .I4(n7744), .O(n7753));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7754 (.I0(x3309), .I1(x3310), .I2(x3311), .I3(n7752), .I4(n7753), .O(n7754));
  LUT3 #(.INIT(8'hE8)) lut_n7755 (.I0(x3318), .I1(x3319), .I2(x3320), .O(n7755));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7756 (.I0(x3309), .I1(x3310), .I2(x3311), .I3(n7752), .I4(n7753), .O(n7756));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7757 (.I0(x3315), .I1(x3316), .I2(x3317), .I3(n7755), .I4(n7756), .O(n7757));
  LUT3 #(.INIT(8'h96)) lut_n7758 (.I0(n7742), .I1(n7745), .I2(n7746), .O(n7758));
  LUT3 #(.INIT(8'hE8)) lut_n7759 (.I0(n7754), .I1(n7757), .I2(n7758), .O(n7759));
  LUT3 #(.INIT(8'hE8)) lut_n7760 (.I0(x3324), .I1(x3325), .I2(x3326), .O(n7760));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7761 (.I0(x3315), .I1(x3316), .I2(x3317), .I3(n7755), .I4(n7756), .O(n7761));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7762 (.I0(x3321), .I1(x3322), .I2(x3323), .I3(n7760), .I4(n7761), .O(n7762));
  LUT3 #(.INIT(8'hE8)) lut_n7763 (.I0(x3330), .I1(x3331), .I2(x3332), .O(n7763));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7764 (.I0(x3321), .I1(x3322), .I2(x3323), .I3(n7760), .I4(n7761), .O(n7764));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7765 (.I0(x3327), .I1(x3328), .I2(x3329), .I3(n7763), .I4(n7764), .O(n7765));
  LUT3 #(.INIT(8'h96)) lut_n7766 (.I0(n7754), .I1(n7757), .I2(n7758), .O(n7766));
  LUT3 #(.INIT(8'hE8)) lut_n7767 (.I0(n7762), .I1(n7765), .I2(n7766), .O(n7767));
  LUT3 #(.INIT(8'h96)) lut_n7768 (.I0(n7739), .I1(n7747), .I2(n7748), .O(n7768));
  LUT3 #(.INIT(8'hE8)) lut_n7769 (.I0(n7759), .I1(n7767), .I2(n7768), .O(n7769));
  LUT3 #(.INIT(8'hE8)) lut_n7770 (.I0(x3336), .I1(x3337), .I2(x3338), .O(n7770));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7771 (.I0(x3327), .I1(x3328), .I2(x3329), .I3(n7763), .I4(n7764), .O(n7771));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7772 (.I0(x3333), .I1(x3334), .I2(x3335), .I3(n7770), .I4(n7771), .O(n7772));
  LUT3 #(.INIT(8'hE8)) lut_n7773 (.I0(x3342), .I1(x3343), .I2(x3344), .O(n7773));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7774 (.I0(x3333), .I1(x3334), .I2(x3335), .I3(n7770), .I4(n7771), .O(n7774));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7775 (.I0(x3339), .I1(x3340), .I2(x3341), .I3(n7773), .I4(n7774), .O(n7775));
  LUT3 #(.INIT(8'h96)) lut_n7776 (.I0(n7762), .I1(n7765), .I2(n7766), .O(n7776));
  LUT3 #(.INIT(8'hE8)) lut_n7777 (.I0(n7772), .I1(n7775), .I2(n7776), .O(n7777));
  LUT3 #(.INIT(8'hE8)) lut_n7778 (.I0(x3348), .I1(x3349), .I2(x3350), .O(n7778));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7779 (.I0(x3339), .I1(x3340), .I2(x3341), .I3(n7773), .I4(n7774), .O(n7779));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7780 (.I0(x3345), .I1(x3346), .I2(x3347), .I3(n7778), .I4(n7779), .O(n7780));
  LUT3 #(.INIT(8'hE8)) lut_n7781 (.I0(x3354), .I1(x3355), .I2(x3356), .O(n7781));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7782 (.I0(x3345), .I1(x3346), .I2(x3347), .I3(n7778), .I4(n7779), .O(n7782));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7783 (.I0(x3351), .I1(x3352), .I2(x3353), .I3(n7781), .I4(n7782), .O(n7783));
  LUT3 #(.INIT(8'h96)) lut_n7784 (.I0(n7772), .I1(n7775), .I2(n7776), .O(n7784));
  LUT3 #(.INIT(8'hE8)) lut_n7785 (.I0(n7780), .I1(n7783), .I2(n7784), .O(n7785));
  LUT3 #(.INIT(8'h96)) lut_n7786 (.I0(n7759), .I1(n7767), .I2(n7768), .O(n7786));
  LUT3 #(.INIT(8'hE8)) lut_n7787 (.I0(n7777), .I1(n7785), .I2(n7786), .O(n7787));
  LUT3 #(.INIT(8'h96)) lut_n7788 (.I0(n7731), .I1(n7749), .I2(n7750), .O(n7788));
  LUT3 #(.INIT(8'hE8)) lut_n7789 (.I0(n7769), .I1(n7787), .I2(n7788), .O(n7789));
  LUT3 #(.INIT(8'h96)) lut_n7790 (.I0(n7671), .I1(n7709), .I2(n7710), .O(n7790));
  LUT3 #(.INIT(8'hE8)) lut_n7791 (.I0(n7751), .I1(n7789), .I2(n7790), .O(n7791));
  LUT3 #(.INIT(8'hE8)) lut_n7792 (.I0(x3360), .I1(x3361), .I2(x3362), .O(n7792));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7793 (.I0(x3351), .I1(x3352), .I2(x3353), .I3(n7781), .I4(n7782), .O(n7793));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7794 (.I0(x3357), .I1(x3358), .I2(x3359), .I3(n7792), .I4(n7793), .O(n7794));
  LUT3 #(.INIT(8'hE8)) lut_n7795 (.I0(x3366), .I1(x3367), .I2(x3368), .O(n7795));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7796 (.I0(x3357), .I1(x3358), .I2(x3359), .I3(n7792), .I4(n7793), .O(n7796));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7797 (.I0(x3363), .I1(x3364), .I2(x3365), .I3(n7795), .I4(n7796), .O(n7797));
  LUT3 #(.INIT(8'h96)) lut_n7798 (.I0(n7780), .I1(n7783), .I2(n7784), .O(n7798));
  LUT3 #(.INIT(8'hE8)) lut_n7799 (.I0(n7794), .I1(n7797), .I2(n7798), .O(n7799));
  LUT3 #(.INIT(8'hE8)) lut_n7800 (.I0(x3372), .I1(x3373), .I2(x3374), .O(n7800));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7801 (.I0(x3363), .I1(x3364), .I2(x3365), .I3(n7795), .I4(n7796), .O(n7801));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7802 (.I0(x3369), .I1(x3370), .I2(x3371), .I3(n7800), .I4(n7801), .O(n7802));
  LUT3 #(.INIT(8'hE8)) lut_n7803 (.I0(x3378), .I1(x3379), .I2(x3380), .O(n7803));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7804 (.I0(x3369), .I1(x3370), .I2(x3371), .I3(n7800), .I4(n7801), .O(n7804));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7805 (.I0(x3375), .I1(x3376), .I2(x3377), .I3(n7803), .I4(n7804), .O(n7805));
  LUT3 #(.INIT(8'h96)) lut_n7806 (.I0(n7794), .I1(n7797), .I2(n7798), .O(n7806));
  LUT3 #(.INIT(8'hE8)) lut_n7807 (.I0(n7802), .I1(n7805), .I2(n7806), .O(n7807));
  LUT3 #(.INIT(8'h96)) lut_n7808 (.I0(n7777), .I1(n7785), .I2(n7786), .O(n7808));
  LUT3 #(.INIT(8'hE8)) lut_n7809 (.I0(n7799), .I1(n7807), .I2(n7808), .O(n7809));
  LUT3 #(.INIT(8'hE8)) lut_n7810 (.I0(x3384), .I1(x3385), .I2(x3386), .O(n7810));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7811 (.I0(x3375), .I1(x3376), .I2(x3377), .I3(n7803), .I4(n7804), .O(n7811));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7812 (.I0(x3381), .I1(x3382), .I2(x3383), .I3(n7810), .I4(n7811), .O(n7812));
  LUT3 #(.INIT(8'hE8)) lut_n7813 (.I0(x3390), .I1(x3391), .I2(x3392), .O(n7813));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7814 (.I0(x3381), .I1(x3382), .I2(x3383), .I3(n7810), .I4(n7811), .O(n7814));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7815 (.I0(x3387), .I1(x3388), .I2(x3389), .I3(n7813), .I4(n7814), .O(n7815));
  LUT3 #(.INIT(8'h96)) lut_n7816 (.I0(n7802), .I1(n7805), .I2(n7806), .O(n7816));
  LUT3 #(.INIT(8'hE8)) lut_n7817 (.I0(n7812), .I1(n7815), .I2(n7816), .O(n7817));
  LUT3 #(.INIT(8'hE8)) lut_n7818 (.I0(x3396), .I1(x3397), .I2(x3398), .O(n7818));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7819 (.I0(x3387), .I1(x3388), .I2(x3389), .I3(n7813), .I4(n7814), .O(n7819));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7820 (.I0(x3393), .I1(x3394), .I2(x3395), .I3(n7818), .I4(n7819), .O(n7820));
  LUT3 #(.INIT(8'hE8)) lut_n7821 (.I0(x3402), .I1(x3403), .I2(x3404), .O(n7821));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7822 (.I0(x3393), .I1(x3394), .I2(x3395), .I3(n7818), .I4(n7819), .O(n7822));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7823 (.I0(x3399), .I1(x3400), .I2(x3401), .I3(n7821), .I4(n7822), .O(n7823));
  LUT3 #(.INIT(8'h96)) lut_n7824 (.I0(n7812), .I1(n7815), .I2(n7816), .O(n7824));
  LUT3 #(.INIT(8'hE8)) lut_n7825 (.I0(n7820), .I1(n7823), .I2(n7824), .O(n7825));
  LUT3 #(.INIT(8'h96)) lut_n7826 (.I0(n7799), .I1(n7807), .I2(n7808), .O(n7826));
  LUT3 #(.INIT(8'hE8)) lut_n7827 (.I0(n7817), .I1(n7825), .I2(n7826), .O(n7827));
  LUT3 #(.INIT(8'h96)) lut_n7828 (.I0(n7769), .I1(n7787), .I2(n7788), .O(n7828));
  LUT3 #(.INIT(8'hE8)) lut_n7829 (.I0(n7809), .I1(n7827), .I2(n7828), .O(n7829));
  LUT3 #(.INIT(8'hE8)) lut_n7830 (.I0(x3408), .I1(x3409), .I2(x3410), .O(n7830));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7831 (.I0(x3399), .I1(x3400), .I2(x3401), .I3(n7821), .I4(n7822), .O(n7831));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7832 (.I0(x3405), .I1(x3406), .I2(x3407), .I3(n7830), .I4(n7831), .O(n7832));
  LUT3 #(.INIT(8'hE8)) lut_n7833 (.I0(x3414), .I1(x3415), .I2(x3416), .O(n7833));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7834 (.I0(x3405), .I1(x3406), .I2(x3407), .I3(n7830), .I4(n7831), .O(n7834));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7835 (.I0(x3411), .I1(x3412), .I2(x3413), .I3(n7833), .I4(n7834), .O(n7835));
  LUT3 #(.INIT(8'h96)) lut_n7836 (.I0(n7820), .I1(n7823), .I2(n7824), .O(n7836));
  LUT3 #(.INIT(8'hE8)) lut_n7837 (.I0(n7832), .I1(n7835), .I2(n7836), .O(n7837));
  LUT3 #(.INIT(8'hE8)) lut_n7838 (.I0(x3420), .I1(x3421), .I2(x3422), .O(n7838));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7839 (.I0(x3411), .I1(x3412), .I2(x3413), .I3(n7833), .I4(n7834), .O(n7839));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7840 (.I0(x3417), .I1(x3418), .I2(x3419), .I3(n7838), .I4(n7839), .O(n7840));
  LUT3 #(.INIT(8'hE8)) lut_n7841 (.I0(x3426), .I1(x3427), .I2(x3428), .O(n7841));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7842 (.I0(x3417), .I1(x3418), .I2(x3419), .I3(n7838), .I4(n7839), .O(n7842));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7843 (.I0(x3423), .I1(x3424), .I2(x3425), .I3(n7841), .I4(n7842), .O(n7843));
  LUT3 #(.INIT(8'h96)) lut_n7844 (.I0(n7832), .I1(n7835), .I2(n7836), .O(n7844));
  LUT3 #(.INIT(8'hE8)) lut_n7845 (.I0(n7840), .I1(n7843), .I2(n7844), .O(n7845));
  LUT3 #(.INIT(8'h96)) lut_n7846 (.I0(n7817), .I1(n7825), .I2(n7826), .O(n7846));
  LUT3 #(.INIT(8'hE8)) lut_n7847 (.I0(n7837), .I1(n7845), .I2(n7846), .O(n7847));
  LUT3 #(.INIT(8'hE8)) lut_n7848 (.I0(x3432), .I1(x3433), .I2(x3434), .O(n7848));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7849 (.I0(x3423), .I1(x3424), .I2(x3425), .I3(n7841), .I4(n7842), .O(n7849));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7850 (.I0(x3429), .I1(x3430), .I2(x3431), .I3(n7848), .I4(n7849), .O(n7850));
  LUT3 #(.INIT(8'hE8)) lut_n7851 (.I0(x3438), .I1(x3439), .I2(x3440), .O(n7851));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7852 (.I0(x3429), .I1(x3430), .I2(x3431), .I3(n7848), .I4(n7849), .O(n7852));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7853 (.I0(x3435), .I1(x3436), .I2(x3437), .I3(n7851), .I4(n7852), .O(n7853));
  LUT3 #(.INIT(8'h96)) lut_n7854 (.I0(n7840), .I1(n7843), .I2(n7844), .O(n7854));
  LUT3 #(.INIT(8'hE8)) lut_n7855 (.I0(n7850), .I1(n7853), .I2(n7854), .O(n7855));
  LUT3 #(.INIT(8'hE8)) lut_n7856 (.I0(x3444), .I1(x3445), .I2(x3446), .O(n7856));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7857 (.I0(x3435), .I1(x3436), .I2(x3437), .I3(n7851), .I4(n7852), .O(n7857));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7858 (.I0(x3441), .I1(x3442), .I2(x3443), .I3(n7856), .I4(n7857), .O(n7858));
  LUT3 #(.INIT(8'hE8)) lut_n7859 (.I0(x3450), .I1(x3451), .I2(x3452), .O(n7859));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7860 (.I0(x3441), .I1(x3442), .I2(x3443), .I3(n7856), .I4(n7857), .O(n7860));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7861 (.I0(x3447), .I1(x3448), .I2(x3449), .I3(n7859), .I4(n7860), .O(n7861));
  LUT3 #(.INIT(8'h96)) lut_n7862 (.I0(n7850), .I1(n7853), .I2(n7854), .O(n7862));
  LUT3 #(.INIT(8'hE8)) lut_n7863 (.I0(n7858), .I1(n7861), .I2(n7862), .O(n7863));
  LUT3 #(.INIT(8'h96)) lut_n7864 (.I0(n7837), .I1(n7845), .I2(n7846), .O(n7864));
  LUT3 #(.INIT(8'hE8)) lut_n7865 (.I0(n7855), .I1(n7863), .I2(n7864), .O(n7865));
  LUT3 #(.INIT(8'h96)) lut_n7866 (.I0(n7809), .I1(n7827), .I2(n7828), .O(n7866));
  LUT3 #(.INIT(8'hE8)) lut_n7867 (.I0(n7847), .I1(n7865), .I2(n7866), .O(n7867));
  LUT3 #(.INIT(8'h96)) lut_n7868 (.I0(n7751), .I1(n7789), .I2(n7790), .O(n7868));
  LUT3 #(.INIT(8'hE8)) lut_n7869 (.I0(n7829), .I1(n7867), .I2(n7868), .O(n7869));
  LUT3 #(.INIT(8'h96)) lut_n7870 (.I0(n7633), .I1(n7711), .I2(n7712), .O(n7870));
  LUT3 #(.INIT(8'hE8)) lut_n7871 (.I0(n7791), .I1(n7869), .I2(n7870), .O(n7871));
  LUT3 #(.INIT(8'h96)) lut_n7872 (.I0(n7392), .I1(n7550), .I2(n7551), .O(n7872));
  LUT3 #(.INIT(8'hE8)) lut_n7873 (.I0(n7713), .I1(n7871), .I2(n7872), .O(n7873));
  LUT3 #(.INIT(8'hE8)) lut_n7874 (.I0(x3456), .I1(x3457), .I2(x3458), .O(n7874));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7875 (.I0(x3447), .I1(x3448), .I2(x3449), .I3(n7859), .I4(n7860), .O(n7875));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7876 (.I0(x3453), .I1(x3454), .I2(x3455), .I3(n7874), .I4(n7875), .O(n7876));
  LUT3 #(.INIT(8'hE8)) lut_n7877 (.I0(x3462), .I1(x3463), .I2(x3464), .O(n7877));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7878 (.I0(x3453), .I1(x3454), .I2(x3455), .I3(n7874), .I4(n7875), .O(n7878));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7879 (.I0(x3459), .I1(x3460), .I2(x3461), .I3(n7877), .I4(n7878), .O(n7879));
  LUT3 #(.INIT(8'h96)) lut_n7880 (.I0(n7858), .I1(n7861), .I2(n7862), .O(n7880));
  LUT3 #(.INIT(8'hE8)) lut_n7881 (.I0(n7876), .I1(n7879), .I2(n7880), .O(n7881));
  LUT3 #(.INIT(8'hE8)) lut_n7882 (.I0(x3468), .I1(x3469), .I2(x3470), .O(n7882));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7883 (.I0(x3459), .I1(x3460), .I2(x3461), .I3(n7877), .I4(n7878), .O(n7883));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7884 (.I0(x3465), .I1(x3466), .I2(x3467), .I3(n7882), .I4(n7883), .O(n7884));
  LUT3 #(.INIT(8'hE8)) lut_n7885 (.I0(x3474), .I1(x3475), .I2(x3476), .O(n7885));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7886 (.I0(x3465), .I1(x3466), .I2(x3467), .I3(n7882), .I4(n7883), .O(n7886));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7887 (.I0(x3471), .I1(x3472), .I2(x3473), .I3(n7885), .I4(n7886), .O(n7887));
  LUT3 #(.INIT(8'h96)) lut_n7888 (.I0(n7876), .I1(n7879), .I2(n7880), .O(n7888));
  LUT3 #(.INIT(8'hE8)) lut_n7889 (.I0(n7884), .I1(n7887), .I2(n7888), .O(n7889));
  LUT3 #(.INIT(8'h96)) lut_n7890 (.I0(n7855), .I1(n7863), .I2(n7864), .O(n7890));
  LUT3 #(.INIT(8'hE8)) lut_n7891 (.I0(n7881), .I1(n7889), .I2(n7890), .O(n7891));
  LUT3 #(.INIT(8'hE8)) lut_n7892 (.I0(x3480), .I1(x3481), .I2(x3482), .O(n7892));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7893 (.I0(x3471), .I1(x3472), .I2(x3473), .I3(n7885), .I4(n7886), .O(n7893));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7894 (.I0(x3477), .I1(x3478), .I2(x3479), .I3(n7892), .I4(n7893), .O(n7894));
  LUT3 #(.INIT(8'hE8)) lut_n7895 (.I0(x3486), .I1(x3487), .I2(x3488), .O(n7895));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7896 (.I0(x3477), .I1(x3478), .I2(x3479), .I3(n7892), .I4(n7893), .O(n7896));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7897 (.I0(x3483), .I1(x3484), .I2(x3485), .I3(n7895), .I4(n7896), .O(n7897));
  LUT3 #(.INIT(8'h96)) lut_n7898 (.I0(n7884), .I1(n7887), .I2(n7888), .O(n7898));
  LUT3 #(.INIT(8'hE8)) lut_n7899 (.I0(n7894), .I1(n7897), .I2(n7898), .O(n7899));
  LUT3 #(.INIT(8'hE8)) lut_n7900 (.I0(x3492), .I1(x3493), .I2(x3494), .O(n7900));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7901 (.I0(x3483), .I1(x3484), .I2(x3485), .I3(n7895), .I4(n7896), .O(n7901));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7902 (.I0(x3489), .I1(x3490), .I2(x3491), .I3(n7900), .I4(n7901), .O(n7902));
  LUT3 #(.INIT(8'hE8)) lut_n7903 (.I0(x3498), .I1(x3499), .I2(x3500), .O(n7903));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7904 (.I0(x3489), .I1(x3490), .I2(x3491), .I3(n7900), .I4(n7901), .O(n7904));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7905 (.I0(x3495), .I1(x3496), .I2(x3497), .I3(n7903), .I4(n7904), .O(n7905));
  LUT3 #(.INIT(8'h96)) lut_n7906 (.I0(n7894), .I1(n7897), .I2(n7898), .O(n7906));
  LUT3 #(.INIT(8'hE8)) lut_n7907 (.I0(n7902), .I1(n7905), .I2(n7906), .O(n7907));
  LUT3 #(.INIT(8'h96)) lut_n7908 (.I0(n7881), .I1(n7889), .I2(n7890), .O(n7908));
  LUT3 #(.INIT(8'hE8)) lut_n7909 (.I0(n7899), .I1(n7907), .I2(n7908), .O(n7909));
  LUT3 #(.INIT(8'h96)) lut_n7910 (.I0(n7847), .I1(n7865), .I2(n7866), .O(n7910));
  LUT3 #(.INIT(8'hE8)) lut_n7911 (.I0(n7891), .I1(n7909), .I2(n7910), .O(n7911));
  LUT3 #(.INIT(8'hE8)) lut_n7912 (.I0(x3504), .I1(x3505), .I2(x3506), .O(n7912));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7913 (.I0(x3495), .I1(x3496), .I2(x3497), .I3(n7903), .I4(n7904), .O(n7913));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7914 (.I0(x3501), .I1(x3502), .I2(x3503), .I3(n7912), .I4(n7913), .O(n7914));
  LUT3 #(.INIT(8'hE8)) lut_n7915 (.I0(x3510), .I1(x3511), .I2(x3512), .O(n7915));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7916 (.I0(x3501), .I1(x3502), .I2(x3503), .I3(n7912), .I4(n7913), .O(n7916));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7917 (.I0(x3507), .I1(x3508), .I2(x3509), .I3(n7915), .I4(n7916), .O(n7917));
  LUT3 #(.INIT(8'h96)) lut_n7918 (.I0(n7902), .I1(n7905), .I2(n7906), .O(n7918));
  LUT3 #(.INIT(8'hE8)) lut_n7919 (.I0(n7914), .I1(n7917), .I2(n7918), .O(n7919));
  LUT3 #(.INIT(8'hE8)) lut_n7920 (.I0(x3516), .I1(x3517), .I2(x3518), .O(n7920));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7921 (.I0(x3507), .I1(x3508), .I2(x3509), .I3(n7915), .I4(n7916), .O(n7921));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7922 (.I0(x3513), .I1(x3514), .I2(x3515), .I3(n7920), .I4(n7921), .O(n7922));
  LUT3 #(.INIT(8'hE8)) lut_n7923 (.I0(x3522), .I1(x3523), .I2(x3524), .O(n7923));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7924 (.I0(x3513), .I1(x3514), .I2(x3515), .I3(n7920), .I4(n7921), .O(n7924));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7925 (.I0(x3519), .I1(x3520), .I2(x3521), .I3(n7923), .I4(n7924), .O(n7925));
  LUT3 #(.INIT(8'h96)) lut_n7926 (.I0(n7914), .I1(n7917), .I2(n7918), .O(n7926));
  LUT3 #(.INIT(8'hE8)) lut_n7927 (.I0(n7922), .I1(n7925), .I2(n7926), .O(n7927));
  LUT3 #(.INIT(8'h96)) lut_n7928 (.I0(n7899), .I1(n7907), .I2(n7908), .O(n7928));
  LUT3 #(.INIT(8'hE8)) lut_n7929 (.I0(n7919), .I1(n7927), .I2(n7928), .O(n7929));
  LUT3 #(.INIT(8'hE8)) lut_n7930 (.I0(x3528), .I1(x3529), .I2(x3530), .O(n7930));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7931 (.I0(x3519), .I1(x3520), .I2(x3521), .I3(n7923), .I4(n7924), .O(n7931));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7932 (.I0(x3525), .I1(x3526), .I2(x3527), .I3(n7930), .I4(n7931), .O(n7932));
  LUT3 #(.INIT(8'hE8)) lut_n7933 (.I0(x3534), .I1(x3535), .I2(x3536), .O(n7933));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7934 (.I0(x3525), .I1(x3526), .I2(x3527), .I3(n7930), .I4(n7931), .O(n7934));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7935 (.I0(x3531), .I1(x3532), .I2(x3533), .I3(n7933), .I4(n7934), .O(n7935));
  LUT3 #(.INIT(8'h96)) lut_n7936 (.I0(n7922), .I1(n7925), .I2(n7926), .O(n7936));
  LUT3 #(.INIT(8'hE8)) lut_n7937 (.I0(n7932), .I1(n7935), .I2(n7936), .O(n7937));
  LUT3 #(.INIT(8'hE8)) lut_n7938 (.I0(x3540), .I1(x3541), .I2(x3542), .O(n7938));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7939 (.I0(x3531), .I1(x3532), .I2(x3533), .I3(n7933), .I4(n7934), .O(n7939));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7940 (.I0(x3537), .I1(x3538), .I2(x3539), .I3(n7938), .I4(n7939), .O(n7940));
  LUT3 #(.INIT(8'hE8)) lut_n7941 (.I0(x3546), .I1(x3547), .I2(x3548), .O(n7941));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7942 (.I0(x3537), .I1(x3538), .I2(x3539), .I3(n7938), .I4(n7939), .O(n7942));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7943 (.I0(x3543), .I1(x3544), .I2(x3545), .I3(n7941), .I4(n7942), .O(n7943));
  LUT3 #(.INIT(8'h96)) lut_n7944 (.I0(n7932), .I1(n7935), .I2(n7936), .O(n7944));
  LUT3 #(.INIT(8'hE8)) lut_n7945 (.I0(n7940), .I1(n7943), .I2(n7944), .O(n7945));
  LUT3 #(.INIT(8'h96)) lut_n7946 (.I0(n7919), .I1(n7927), .I2(n7928), .O(n7946));
  LUT3 #(.INIT(8'hE8)) lut_n7947 (.I0(n7937), .I1(n7945), .I2(n7946), .O(n7947));
  LUT3 #(.INIT(8'h96)) lut_n7948 (.I0(n7891), .I1(n7909), .I2(n7910), .O(n7948));
  LUT3 #(.INIT(8'hE8)) lut_n7949 (.I0(n7929), .I1(n7947), .I2(n7948), .O(n7949));
  LUT3 #(.INIT(8'h96)) lut_n7950 (.I0(n7829), .I1(n7867), .I2(n7868), .O(n7950));
  LUT3 #(.INIT(8'hE8)) lut_n7951 (.I0(n7911), .I1(n7949), .I2(n7950), .O(n7951));
  LUT3 #(.INIT(8'hE8)) lut_n7952 (.I0(x3552), .I1(x3553), .I2(x3554), .O(n7952));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7953 (.I0(x3543), .I1(x3544), .I2(x3545), .I3(n7941), .I4(n7942), .O(n7953));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7954 (.I0(x3549), .I1(x3550), .I2(x3551), .I3(n7952), .I4(n7953), .O(n7954));
  LUT3 #(.INIT(8'hE8)) lut_n7955 (.I0(x3558), .I1(x3559), .I2(x3560), .O(n7955));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7956 (.I0(x3549), .I1(x3550), .I2(x3551), .I3(n7952), .I4(n7953), .O(n7956));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7957 (.I0(x3555), .I1(x3556), .I2(x3557), .I3(n7955), .I4(n7956), .O(n7957));
  LUT3 #(.INIT(8'h96)) lut_n7958 (.I0(n7940), .I1(n7943), .I2(n7944), .O(n7958));
  LUT3 #(.INIT(8'hE8)) lut_n7959 (.I0(n7954), .I1(n7957), .I2(n7958), .O(n7959));
  LUT3 #(.INIT(8'hE8)) lut_n7960 (.I0(x3564), .I1(x3565), .I2(x3566), .O(n7960));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7961 (.I0(x3555), .I1(x3556), .I2(x3557), .I3(n7955), .I4(n7956), .O(n7961));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7962 (.I0(x3561), .I1(x3562), .I2(x3563), .I3(n7960), .I4(n7961), .O(n7962));
  LUT3 #(.INIT(8'hE8)) lut_n7963 (.I0(x3570), .I1(x3571), .I2(x3572), .O(n7963));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7964 (.I0(x3561), .I1(x3562), .I2(x3563), .I3(n7960), .I4(n7961), .O(n7964));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7965 (.I0(x3567), .I1(x3568), .I2(x3569), .I3(n7963), .I4(n7964), .O(n7965));
  LUT3 #(.INIT(8'h96)) lut_n7966 (.I0(n7954), .I1(n7957), .I2(n7958), .O(n7966));
  LUT3 #(.INIT(8'hE8)) lut_n7967 (.I0(n7962), .I1(n7965), .I2(n7966), .O(n7967));
  LUT3 #(.INIT(8'h96)) lut_n7968 (.I0(n7937), .I1(n7945), .I2(n7946), .O(n7968));
  LUT3 #(.INIT(8'hE8)) lut_n7969 (.I0(n7959), .I1(n7967), .I2(n7968), .O(n7969));
  LUT3 #(.INIT(8'hE8)) lut_n7970 (.I0(x3576), .I1(x3577), .I2(x3578), .O(n7970));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7971 (.I0(x3567), .I1(x3568), .I2(x3569), .I3(n7963), .I4(n7964), .O(n7971));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7972 (.I0(x3573), .I1(x3574), .I2(x3575), .I3(n7970), .I4(n7971), .O(n7972));
  LUT3 #(.INIT(8'hE8)) lut_n7973 (.I0(x3582), .I1(x3583), .I2(x3584), .O(n7973));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7974 (.I0(x3573), .I1(x3574), .I2(x3575), .I3(n7970), .I4(n7971), .O(n7974));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7975 (.I0(x3579), .I1(x3580), .I2(x3581), .I3(n7973), .I4(n7974), .O(n7975));
  LUT3 #(.INIT(8'h96)) lut_n7976 (.I0(n7962), .I1(n7965), .I2(n7966), .O(n7976));
  LUT3 #(.INIT(8'hE8)) lut_n7977 (.I0(n7972), .I1(n7975), .I2(n7976), .O(n7977));
  LUT3 #(.INIT(8'hE8)) lut_n7978 (.I0(x3588), .I1(x3589), .I2(x3590), .O(n7978));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7979 (.I0(x3579), .I1(x3580), .I2(x3581), .I3(n7973), .I4(n7974), .O(n7979));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7980 (.I0(x3585), .I1(x3586), .I2(x3587), .I3(n7978), .I4(n7979), .O(n7980));
  LUT3 #(.INIT(8'hE8)) lut_n7981 (.I0(x3594), .I1(x3595), .I2(x3596), .O(n7981));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7982 (.I0(x3585), .I1(x3586), .I2(x3587), .I3(n7978), .I4(n7979), .O(n7982));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7983 (.I0(x3591), .I1(x3592), .I2(x3593), .I3(n7981), .I4(n7982), .O(n7983));
  LUT3 #(.INIT(8'h96)) lut_n7984 (.I0(n7972), .I1(n7975), .I2(n7976), .O(n7984));
  LUT3 #(.INIT(8'hE8)) lut_n7985 (.I0(n7980), .I1(n7983), .I2(n7984), .O(n7985));
  LUT3 #(.INIT(8'h96)) lut_n7986 (.I0(n7959), .I1(n7967), .I2(n7968), .O(n7986));
  LUT3 #(.INIT(8'hE8)) lut_n7987 (.I0(n7977), .I1(n7985), .I2(n7986), .O(n7987));
  LUT3 #(.INIT(8'h96)) lut_n7988 (.I0(n7929), .I1(n7947), .I2(n7948), .O(n7988));
  LUT3 #(.INIT(8'hE8)) lut_n7989 (.I0(n7969), .I1(n7987), .I2(n7988), .O(n7989));
  LUT3 #(.INIT(8'hE8)) lut_n7990 (.I0(x3600), .I1(x3601), .I2(x3602), .O(n7990));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7991 (.I0(x3591), .I1(x3592), .I2(x3593), .I3(n7981), .I4(n7982), .O(n7991));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7992 (.I0(x3597), .I1(x3598), .I2(x3599), .I3(n7990), .I4(n7991), .O(n7992));
  LUT3 #(.INIT(8'hE8)) lut_n7993 (.I0(x3606), .I1(x3607), .I2(x3608), .O(n7993));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7994 (.I0(x3597), .I1(x3598), .I2(x3599), .I3(n7990), .I4(n7991), .O(n7994));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n7995 (.I0(x3603), .I1(x3604), .I2(x3605), .I3(n7993), .I4(n7994), .O(n7995));
  LUT3 #(.INIT(8'h96)) lut_n7996 (.I0(n7980), .I1(n7983), .I2(n7984), .O(n7996));
  LUT3 #(.INIT(8'hE8)) lut_n7997 (.I0(n7992), .I1(n7995), .I2(n7996), .O(n7997));
  LUT3 #(.INIT(8'hE8)) lut_n7998 (.I0(x3612), .I1(x3613), .I2(x3614), .O(n7998));
  LUT5 #(.INIT(32'hE81717E8)) lut_n7999 (.I0(x3603), .I1(x3604), .I2(x3605), .I3(n7993), .I4(n7994), .O(n7999));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8000 (.I0(x3609), .I1(x3610), .I2(x3611), .I3(n7998), .I4(n7999), .O(n8000));
  LUT3 #(.INIT(8'hE8)) lut_n8001 (.I0(x3618), .I1(x3619), .I2(x3620), .O(n8001));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8002 (.I0(x3609), .I1(x3610), .I2(x3611), .I3(n7998), .I4(n7999), .O(n8002));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8003 (.I0(x3615), .I1(x3616), .I2(x3617), .I3(n8001), .I4(n8002), .O(n8003));
  LUT3 #(.INIT(8'h96)) lut_n8004 (.I0(n7992), .I1(n7995), .I2(n7996), .O(n8004));
  LUT3 #(.INIT(8'hE8)) lut_n8005 (.I0(n8000), .I1(n8003), .I2(n8004), .O(n8005));
  LUT3 #(.INIT(8'h96)) lut_n8006 (.I0(n7977), .I1(n7985), .I2(n7986), .O(n8006));
  LUT3 #(.INIT(8'hE8)) lut_n8007 (.I0(n7997), .I1(n8005), .I2(n8006), .O(n8007));
  LUT3 #(.INIT(8'hE8)) lut_n8008 (.I0(x3624), .I1(x3625), .I2(x3626), .O(n8008));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8009 (.I0(x3615), .I1(x3616), .I2(x3617), .I3(n8001), .I4(n8002), .O(n8009));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8010 (.I0(x3621), .I1(x3622), .I2(x3623), .I3(n8008), .I4(n8009), .O(n8010));
  LUT3 #(.INIT(8'hE8)) lut_n8011 (.I0(x3630), .I1(x3631), .I2(x3632), .O(n8011));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8012 (.I0(x3621), .I1(x3622), .I2(x3623), .I3(n8008), .I4(n8009), .O(n8012));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8013 (.I0(x3627), .I1(x3628), .I2(x3629), .I3(n8011), .I4(n8012), .O(n8013));
  LUT3 #(.INIT(8'h96)) lut_n8014 (.I0(n8000), .I1(n8003), .I2(n8004), .O(n8014));
  LUT3 #(.INIT(8'hE8)) lut_n8015 (.I0(n8010), .I1(n8013), .I2(n8014), .O(n8015));
  LUT3 #(.INIT(8'hE8)) lut_n8016 (.I0(x3636), .I1(x3637), .I2(x3638), .O(n8016));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8017 (.I0(x3627), .I1(x3628), .I2(x3629), .I3(n8011), .I4(n8012), .O(n8017));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8018 (.I0(x3633), .I1(x3634), .I2(x3635), .I3(n8016), .I4(n8017), .O(n8018));
  LUT3 #(.INIT(8'hE8)) lut_n8019 (.I0(x3642), .I1(x3643), .I2(x3644), .O(n8019));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8020 (.I0(x3633), .I1(x3634), .I2(x3635), .I3(n8016), .I4(n8017), .O(n8020));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8021 (.I0(x3639), .I1(x3640), .I2(x3641), .I3(n8019), .I4(n8020), .O(n8021));
  LUT3 #(.INIT(8'h96)) lut_n8022 (.I0(n8010), .I1(n8013), .I2(n8014), .O(n8022));
  LUT3 #(.INIT(8'hE8)) lut_n8023 (.I0(n8018), .I1(n8021), .I2(n8022), .O(n8023));
  LUT3 #(.INIT(8'h96)) lut_n8024 (.I0(n7997), .I1(n8005), .I2(n8006), .O(n8024));
  LUT3 #(.INIT(8'hE8)) lut_n8025 (.I0(n8015), .I1(n8023), .I2(n8024), .O(n8025));
  LUT3 #(.INIT(8'h96)) lut_n8026 (.I0(n7969), .I1(n7987), .I2(n7988), .O(n8026));
  LUT3 #(.INIT(8'hE8)) lut_n8027 (.I0(n8007), .I1(n8025), .I2(n8026), .O(n8027));
  LUT3 #(.INIT(8'h96)) lut_n8028 (.I0(n7911), .I1(n7949), .I2(n7950), .O(n8028));
  LUT3 #(.INIT(8'hE8)) lut_n8029 (.I0(n7989), .I1(n8027), .I2(n8028), .O(n8029));
  LUT3 #(.INIT(8'h96)) lut_n8030 (.I0(n7791), .I1(n7869), .I2(n7870), .O(n8030));
  LUT3 #(.INIT(8'hE8)) lut_n8031 (.I0(n7951), .I1(n8029), .I2(n8030), .O(n8031));
  LUT3 #(.INIT(8'hE8)) lut_n8032 (.I0(x3648), .I1(x3649), .I2(x3650), .O(n8032));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8033 (.I0(x3639), .I1(x3640), .I2(x3641), .I3(n8019), .I4(n8020), .O(n8033));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8034 (.I0(x3645), .I1(x3646), .I2(x3647), .I3(n8032), .I4(n8033), .O(n8034));
  LUT3 #(.INIT(8'hE8)) lut_n8035 (.I0(x3654), .I1(x3655), .I2(x3656), .O(n8035));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8036 (.I0(x3645), .I1(x3646), .I2(x3647), .I3(n8032), .I4(n8033), .O(n8036));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8037 (.I0(x3651), .I1(x3652), .I2(x3653), .I3(n8035), .I4(n8036), .O(n8037));
  LUT3 #(.INIT(8'h96)) lut_n8038 (.I0(n8018), .I1(n8021), .I2(n8022), .O(n8038));
  LUT3 #(.INIT(8'hE8)) lut_n8039 (.I0(n8034), .I1(n8037), .I2(n8038), .O(n8039));
  LUT3 #(.INIT(8'hE8)) lut_n8040 (.I0(x3660), .I1(x3661), .I2(x3662), .O(n8040));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8041 (.I0(x3651), .I1(x3652), .I2(x3653), .I3(n8035), .I4(n8036), .O(n8041));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8042 (.I0(x3657), .I1(x3658), .I2(x3659), .I3(n8040), .I4(n8041), .O(n8042));
  LUT3 #(.INIT(8'hE8)) lut_n8043 (.I0(x3666), .I1(x3667), .I2(x3668), .O(n8043));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8044 (.I0(x3657), .I1(x3658), .I2(x3659), .I3(n8040), .I4(n8041), .O(n8044));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8045 (.I0(x3663), .I1(x3664), .I2(x3665), .I3(n8043), .I4(n8044), .O(n8045));
  LUT3 #(.INIT(8'h96)) lut_n8046 (.I0(n8034), .I1(n8037), .I2(n8038), .O(n8046));
  LUT3 #(.INIT(8'hE8)) lut_n8047 (.I0(n8042), .I1(n8045), .I2(n8046), .O(n8047));
  LUT3 #(.INIT(8'h96)) lut_n8048 (.I0(n8015), .I1(n8023), .I2(n8024), .O(n8048));
  LUT3 #(.INIT(8'hE8)) lut_n8049 (.I0(n8039), .I1(n8047), .I2(n8048), .O(n8049));
  LUT3 #(.INIT(8'hE8)) lut_n8050 (.I0(x3672), .I1(x3673), .I2(x3674), .O(n8050));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8051 (.I0(x3663), .I1(x3664), .I2(x3665), .I3(n8043), .I4(n8044), .O(n8051));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8052 (.I0(x3669), .I1(x3670), .I2(x3671), .I3(n8050), .I4(n8051), .O(n8052));
  LUT3 #(.INIT(8'hE8)) lut_n8053 (.I0(x3678), .I1(x3679), .I2(x3680), .O(n8053));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8054 (.I0(x3669), .I1(x3670), .I2(x3671), .I3(n8050), .I4(n8051), .O(n8054));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8055 (.I0(x3675), .I1(x3676), .I2(x3677), .I3(n8053), .I4(n8054), .O(n8055));
  LUT3 #(.INIT(8'h96)) lut_n8056 (.I0(n8042), .I1(n8045), .I2(n8046), .O(n8056));
  LUT3 #(.INIT(8'hE8)) lut_n8057 (.I0(n8052), .I1(n8055), .I2(n8056), .O(n8057));
  LUT3 #(.INIT(8'hE8)) lut_n8058 (.I0(x3684), .I1(x3685), .I2(x3686), .O(n8058));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8059 (.I0(x3675), .I1(x3676), .I2(x3677), .I3(n8053), .I4(n8054), .O(n8059));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8060 (.I0(x3681), .I1(x3682), .I2(x3683), .I3(n8058), .I4(n8059), .O(n8060));
  LUT3 #(.INIT(8'hE8)) lut_n8061 (.I0(x3690), .I1(x3691), .I2(x3692), .O(n8061));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8062 (.I0(x3681), .I1(x3682), .I2(x3683), .I3(n8058), .I4(n8059), .O(n8062));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8063 (.I0(x3687), .I1(x3688), .I2(x3689), .I3(n8061), .I4(n8062), .O(n8063));
  LUT3 #(.INIT(8'h96)) lut_n8064 (.I0(n8052), .I1(n8055), .I2(n8056), .O(n8064));
  LUT3 #(.INIT(8'hE8)) lut_n8065 (.I0(n8060), .I1(n8063), .I2(n8064), .O(n8065));
  LUT3 #(.INIT(8'h96)) lut_n8066 (.I0(n8039), .I1(n8047), .I2(n8048), .O(n8066));
  LUT3 #(.INIT(8'hE8)) lut_n8067 (.I0(n8057), .I1(n8065), .I2(n8066), .O(n8067));
  LUT3 #(.INIT(8'h96)) lut_n8068 (.I0(n8007), .I1(n8025), .I2(n8026), .O(n8068));
  LUT3 #(.INIT(8'hE8)) lut_n8069 (.I0(n8049), .I1(n8067), .I2(n8068), .O(n8069));
  LUT3 #(.INIT(8'hE8)) lut_n8070 (.I0(x3696), .I1(x3697), .I2(x3698), .O(n8070));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8071 (.I0(x3687), .I1(x3688), .I2(x3689), .I3(n8061), .I4(n8062), .O(n8071));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8072 (.I0(x3693), .I1(x3694), .I2(x3695), .I3(n8070), .I4(n8071), .O(n8072));
  LUT3 #(.INIT(8'hE8)) lut_n8073 (.I0(x3702), .I1(x3703), .I2(x3704), .O(n8073));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8074 (.I0(x3693), .I1(x3694), .I2(x3695), .I3(n8070), .I4(n8071), .O(n8074));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8075 (.I0(x3699), .I1(x3700), .I2(x3701), .I3(n8073), .I4(n8074), .O(n8075));
  LUT3 #(.INIT(8'h96)) lut_n8076 (.I0(n8060), .I1(n8063), .I2(n8064), .O(n8076));
  LUT3 #(.INIT(8'hE8)) lut_n8077 (.I0(n8072), .I1(n8075), .I2(n8076), .O(n8077));
  LUT3 #(.INIT(8'hE8)) lut_n8078 (.I0(x3708), .I1(x3709), .I2(x3710), .O(n8078));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8079 (.I0(x3699), .I1(x3700), .I2(x3701), .I3(n8073), .I4(n8074), .O(n8079));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8080 (.I0(x3705), .I1(x3706), .I2(x3707), .I3(n8078), .I4(n8079), .O(n8080));
  LUT3 #(.INIT(8'hE8)) lut_n8081 (.I0(x3714), .I1(x3715), .I2(x3716), .O(n8081));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8082 (.I0(x3705), .I1(x3706), .I2(x3707), .I3(n8078), .I4(n8079), .O(n8082));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8083 (.I0(x3711), .I1(x3712), .I2(x3713), .I3(n8081), .I4(n8082), .O(n8083));
  LUT3 #(.INIT(8'h96)) lut_n8084 (.I0(n8072), .I1(n8075), .I2(n8076), .O(n8084));
  LUT3 #(.INIT(8'hE8)) lut_n8085 (.I0(n8080), .I1(n8083), .I2(n8084), .O(n8085));
  LUT3 #(.INIT(8'h96)) lut_n8086 (.I0(n8057), .I1(n8065), .I2(n8066), .O(n8086));
  LUT3 #(.INIT(8'hE8)) lut_n8087 (.I0(n8077), .I1(n8085), .I2(n8086), .O(n8087));
  LUT3 #(.INIT(8'hE8)) lut_n8088 (.I0(x3720), .I1(x3721), .I2(x3722), .O(n8088));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8089 (.I0(x3711), .I1(x3712), .I2(x3713), .I3(n8081), .I4(n8082), .O(n8089));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8090 (.I0(x3717), .I1(x3718), .I2(x3719), .I3(n8088), .I4(n8089), .O(n8090));
  LUT3 #(.INIT(8'hE8)) lut_n8091 (.I0(x3726), .I1(x3727), .I2(x3728), .O(n8091));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8092 (.I0(x3717), .I1(x3718), .I2(x3719), .I3(n8088), .I4(n8089), .O(n8092));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8093 (.I0(x3723), .I1(x3724), .I2(x3725), .I3(n8091), .I4(n8092), .O(n8093));
  LUT3 #(.INIT(8'h96)) lut_n8094 (.I0(n8080), .I1(n8083), .I2(n8084), .O(n8094));
  LUT3 #(.INIT(8'hE8)) lut_n8095 (.I0(n8090), .I1(n8093), .I2(n8094), .O(n8095));
  LUT3 #(.INIT(8'hE8)) lut_n8096 (.I0(x3732), .I1(x3733), .I2(x3734), .O(n8096));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8097 (.I0(x3723), .I1(x3724), .I2(x3725), .I3(n8091), .I4(n8092), .O(n8097));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8098 (.I0(x3729), .I1(x3730), .I2(x3731), .I3(n8096), .I4(n8097), .O(n8098));
  LUT3 #(.INIT(8'hE8)) lut_n8099 (.I0(x3738), .I1(x3739), .I2(x3740), .O(n8099));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8100 (.I0(x3729), .I1(x3730), .I2(x3731), .I3(n8096), .I4(n8097), .O(n8100));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8101 (.I0(x3735), .I1(x3736), .I2(x3737), .I3(n8099), .I4(n8100), .O(n8101));
  LUT3 #(.INIT(8'h96)) lut_n8102 (.I0(n8090), .I1(n8093), .I2(n8094), .O(n8102));
  LUT3 #(.INIT(8'hE8)) lut_n8103 (.I0(n8098), .I1(n8101), .I2(n8102), .O(n8103));
  LUT3 #(.INIT(8'h96)) lut_n8104 (.I0(n8077), .I1(n8085), .I2(n8086), .O(n8104));
  LUT3 #(.INIT(8'hE8)) lut_n8105 (.I0(n8095), .I1(n8103), .I2(n8104), .O(n8105));
  LUT3 #(.INIT(8'h96)) lut_n8106 (.I0(n8049), .I1(n8067), .I2(n8068), .O(n8106));
  LUT3 #(.INIT(8'hE8)) lut_n8107 (.I0(n8087), .I1(n8105), .I2(n8106), .O(n8107));
  LUT3 #(.INIT(8'h96)) lut_n8108 (.I0(n7989), .I1(n8027), .I2(n8028), .O(n8108));
  LUT3 #(.INIT(8'hE8)) lut_n8109 (.I0(n8069), .I1(n8107), .I2(n8108), .O(n8109));
  LUT3 #(.INIT(8'hE8)) lut_n8110 (.I0(x3744), .I1(x3745), .I2(x3746), .O(n8110));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8111 (.I0(x3735), .I1(x3736), .I2(x3737), .I3(n8099), .I4(n8100), .O(n8111));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8112 (.I0(x3741), .I1(x3742), .I2(x3743), .I3(n8110), .I4(n8111), .O(n8112));
  LUT3 #(.INIT(8'hE8)) lut_n8113 (.I0(x3750), .I1(x3751), .I2(x3752), .O(n8113));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8114 (.I0(x3741), .I1(x3742), .I2(x3743), .I3(n8110), .I4(n8111), .O(n8114));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8115 (.I0(x3747), .I1(x3748), .I2(x3749), .I3(n8113), .I4(n8114), .O(n8115));
  LUT3 #(.INIT(8'h96)) lut_n8116 (.I0(n8098), .I1(n8101), .I2(n8102), .O(n8116));
  LUT3 #(.INIT(8'hE8)) lut_n8117 (.I0(n8112), .I1(n8115), .I2(n8116), .O(n8117));
  LUT3 #(.INIT(8'hE8)) lut_n8118 (.I0(x3756), .I1(x3757), .I2(x3758), .O(n8118));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8119 (.I0(x3747), .I1(x3748), .I2(x3749), .I3(n8113), .I4(n8114), .O(n8119));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8120 (.I0(x3753), .I1(x3754), .I2(x3755), .I3(n8118), .I4(n8119), .O(n8120));
  LUT3 #(.INIT(8'hE8)) lut_n8121 (.I0(x3762), .I1(x3763), .I2(x3764), .O(n8121));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8122 (.I0(x3753), .I1(x3754), .I2(x3755), .I3(n8118), .I4(n8119), .O(n8122));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8123 (.I0(x3759), .I1(x3760), .I2(x3761), .I3(n8121), .I4(n8122), .O(n8123));
  LUT3 #(.INIT(8'h96)) lut_n8124 (.I0(n8112), .I1(n8115), .I2(n8116), .O(n8124));
  LUT3 #(.INIT(8'hE8)) lut_n8125 (.I0(n8120), .I1(n8123), .I2(n8124), .O(n8125));
  LUT3 #(.INIT(8'h96)) lut_n8126 (.I0(n8095), .I1(n8103), .I2(n8104), .O(n8126));
  LUT3 #(.INIT(8'hE8)) lut_n8127 (.I0(n8117), .I1(n8125), .I2(n8126), .O(n8127));
  LUT3 #(.INIT(8'hE8)) lut_n8128 (.I0(x3768), .I1(x3769), .I2(x3770), .O(n8128));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8129 (.I0(x3759), .I1(x3760), .I2(x3761), .I3(n8121), .I4(n8122), .O(n8129));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8130 (.I0(x3765), .I1(x3766), .I2(x3767), .I3(n8128), .I4(n8129), .O(n8130));
  LUT3 #(.INIT(8'hE8)) lut_n8131 (.I0(x3774), .I1(x3775), .I2(x3776), .O(n8131));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8132 (.I0(x3765), .I1(x3766), .I2(x3767), .I3(n8128), .I4(n8129), .O(n8132));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8133 (.I0(x3771), .I1(x3772), .I2(x3773), .I3(n8131), .I4(n8132), .O(n8133));
  LUT3 #(.INIT(8'h96)) lut_n8134 (.I0(n8120), .I1(n8123), .I2(n8124), .O(n8134));
  LUT3 #(.INIT(8'hE8)) lut_n8135 (.I0(n8130), .I1(n8133), .I2(n8134), .O(n8135));
  LUT3 #(.INIT(8'hE8)) lut_n8136 (.I0(x3780), .I1(x3781), .I2(x3782), .O(n8136));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8137 (.I0(x3771), .I1(x3772), .I2(x3773), .I3(n8131), .I4(n8132), .O(n8137));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8138 (.I0(x3777), .I1(x3778), .I2(x3779), .I3(n8136), .I4(n8137), .O(n8138));
  LUT3 #(.INIT(8'hE8)) lut_n8139 (.I0(x3786), .I1(x3787), .I2(x3788), .O(n8139));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8140 (.I0(x3777), .I1(x3778), .I2(x3779), .I3(n8136), .I4(n8137), .O(n8140));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8141 (.I0(x3783), .I1(x3784), .I2(x3785), .I3(n8139), .I4(n8140), .O(n8141));
  LUT3 #(.INIT(8'h96)) lut_n8142 (.I0(n8130), .I1(n8133), .I2(n8134), .O(n8142));
  LUT3 #(.INIT(8'hE8)) lut_n8143 (.I0(n8138), .I1(n8141), .I2(n8142), .O(n8143));
  LUT3 #(.INIT(8'h96)) lut_n8144 (.I0(n8117), .I1(n8125), .I2(n8126), .O(n8144));
  LUT3 #(.INIT(8'hE8)) lut_n8145 (.I0(n8135), .I1(n8143), .I2(n8144), .O(n8145));
  LUT3 #(.INIT(8'h96)) lut_n8146 (.I0(n8087), .I1(n8105), .I2(n8106), .O(n8146));
  LUT3 #(.INIT(8'hE8)) lut_n8147 (.I0(n8127), .I1(n8145), .I2(n8146), .O(n8147));
  LUT3 #(.INIT(8'hE8)) lut_n8148 (.I0(x3792), .I1(x3793), .I2(x3794), .O(n8148));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8149 (.I0(x3783), .I1(x3784), .I2(x3785), .I3(n8139), .I4(n8140), .O(n8149));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8150 (.I0(x3789), .I1(x3790), .I2(x3791), .I3(n8148), .I4(n8149), .O(n8150));
  LUT3 #(.INIT(8'hE8)) lut_n8151 (.I0(x3798), .I1(x3799), .I2(x3800), .O(n8151));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8152 (.I0(x3789), .I1(x3790), .I2(x3791), .I3(n8148), .I4(n8149), .O(n8152));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8153 (.I0(x3795), .I1(x3796), .I2(x3797), .I3(n8151), .I4(n8152), .O(n8153));
  LUT3 #(.INIT(8'h96)) lut_n8154 (.I0(n8138), .I1(n8141), .I2(n8142), .O(n8154));
  LUT3 #(.INIT(8'hE8)) lut_n8155 (.I0(n8150), .I1(n8153), .I2(n8154), .O(n8155));
  LUT3 #(.INIT(8'hE8)) lut_n8156 (.I0(x3804), .I1(x3805), .I2(x3806), .O(n8156));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8157 (.I0(x3795), .I1(x3796), .I2(x3797), .I3(n8151), .I4(n8152), .O(n8157));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8158 (.I0(x3801), .I1(x3802), .I2(x3803), .I3(n8156), .I4(n8157), .O(n8158));
  LUT3 #(.INIT(8'hE8)) lut_n8159 (.I0(x3810), .I1(x3811), .I2(x3812), .O(n8159));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8160 (.I0(x3801), .I1(x3802), .I2(x3803), .I3(n8156), .I4(n8157), .O(n8160));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8161 (.I0(x3807), .I1(x3808), .I2(x3809), .I3(n8159), .I4(n8160), .O(n8161));
  LUT3 #(.INIT(8'h96)) lut_n8162 (.I0(n8150), .I1(n8153), .I2(n8154), .O(n8162));
  LUT3 #(.INIT(8'hE8)) lut_n8163 (.I0(n8158), .I1(n8161), .I2(n8162), .O(n8163));
  LUT3 #(.INIT(8'h96)) lut_n8164 (.I0(n8135), .I1(n8143), .I2(n8144), .O(n8164));
  LUT3 #(.INIT(8'hE8)) lut_n8165 (.I0(n8155), .I1(n8163), .I2(n8164), .O(n8165));
  LUT3 #(.INIT(8'hE8)) lut_n8166 (.I0(x3816), .I1(x3817), .I2(x3818), .O(n8166));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8167 (.I0(x3807), .I1(x3808), .I2(x3809), .I3(n8159), .I4(n8160), .O(n8167));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8168 (.I0(x3813), .I1(x3814), .I2(x3815), .I3(n8166), .I4(n8167), .O(n8168));
  LUT3 #(.INIT(8'hE8)) lut_n8169 (.I0(x3822), .I1(x3823), .I2(x3824), .O(n8169));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8170 (.I0(x3813), .I1(x3814), .I2(x3815), .I3(n8166), .I4(n8167), .O(n8170));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8171 (.I0(x3819), .I1(x3820), .I2(x3821), .I3(n8169), .I4(n8170), .O(n8171));
  LUT3 #(.INIT(8'h96)) lut_n8172 (.I0(n8158), .I1(n8161), .I2(n8162), .O(n8172));
  LUT3 #(.INIT(8'hE8)) lut_n8173 (.I0(n8168), .I1(n8171), .I2(n8172), .O(n8173));
  LUT3 #(.INIT(8'hE8)) lut_n8174 (.I0(x3828), .I1(x3829), .I2(x3830), .O(n8174));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8175 (.I0(x3819), .I1(x3820), .I2(x3821), .I3(n8169), .I4(n8170), .O(n8175));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8176 (.I0(x3825), .I1(x3826), .I2(x3827), .I3(n8174), .I4(n8175), .O(n8176));
  LUT3 #(.INIT(8'hE8)) lut_n8177 (.I0(x3834), .I1(x3835), .I2(x3836), .O(n8177));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8178 (.I0(x3825), .I1(x3826), .I2(x3827), .I3(n8174), .I4(n8175), .O(n8178));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8179 (.I0(x3831), .I1(x3832), .I2(x3833), .I3(n8177), .I4(n8178), .O(n8179));
  LUT3 #(.INIT(8'h96)) lut_n8180 (.I0(n8168), .I1(n8171), .I2(n8172), .O(n8180));
  LUT3 #(.INIT(8'hE8)) lut_n8181 (.I0(n8176), .I1(n8179), .I2(n8180), .O(n8181));
  LUT3 #(.INIT(8'h96)) lut_n8182 (.I0(n8155), .I1(n8163), .I2(n8164), .O(n8182));
  LUT3 #(.INIT(8'hE8)) lut_n8183 (.I0(n8173), .I1(n8181), .I2(n8182), .O(n8183));
  LUT3 #(.INIT(8'h96)) lut_n8184 (.I0(n8127), .I1(n8145), .I2(n8146), .O(n8184));
  LUT3 #(.INIT(8'hE8)) lut_n8185 (.I0(n8165), .I1(n8183), .I2(n8184), .O(n8185));
  LUT3 #(.INIT(8'h96)) lut_n8186 (.I0(n8069), .I1(n8107), .I2(n8108), .O(n8186));
  LUT3 #(.INIT(8'hE8)) lut_n8187 (.I0(n8147), .I1(n8185), .I2(n8186), .O(n8187));
  LUT3 #(.INIT(8'h96)) lut_n8188 (.I0(n7951), .I1(n8029), .I2(n8030), .O(n8188));
  LUT3 #(.INIT(8'hE8)) lut_n8189 (.I0(n8109), .I1(n8187), .I2(n8188), .O(n8189));
  LUT3 #(.INIT(8'h96)) lut_n8190 (.I0(n7713), .I1(n7871), .I2(n7872), .O(n8190));
  LUT3 #(.INIT(8'hE8)) lut_n8191 (.I0(n8031), .I1(n8189), .I2(n8190), .O(n8191));
  LUT3 #(.INIT(8'h96)) lut_n8192 (.I0(n7234), .I1(n7552), .I2(n7553), .O(n8192));
  LUT3 #(.INIT(8'hE8)) lut_n8193 (.I0(n7873), .I1(n8191), .I2(n8192), .O(n8193));
  LUT3 #(.INIT(8'hE8)) lut_n8194 (.I0(x3840), .I1(x3841), .I2(x3842), .O(n8194));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8195 (.I0(x3831), .I1(x3832), .I2(x3833), .I3(n8177), .I4(n8178), .O(n8195));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8196 (.I0(x3837), .I1(x3838), .I2(x3839), .I3(n8194), .I4(n8195), .O(n8196));
  LUT3 #(.INIT(8'hE8)) lut_n8197 (.I0(x3846), .I1(x3847), .I2(x3848), .O(n8197));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8198 (.I0(x3837), .I1(x3838), .I2(x3839), .I3(n8194), .I4(n8195), .O(n8198));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8199 (.I0(x3843), .I1(x3844), .I2(x3845), .I3(n8197), .I4(n8198), .O(n8199));
  LUT3 #(.INIT(8'h96)) lut_n8200 (.I0(n8176), .I1(n8179), .I2(n8180), .O(n8200));
  LUT3 #(.INIT(8'hE8)) lut_n8201 (.I0(n8196), .I1(n8199), .I2(n8200), .O(n8201));
  LUT3 #(.INIT(8'hE8)) lut_n8202 (.I0(x3852), .I1(x3853), .I2(x3854), .O(n8202));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8203 (.I0(x3843), .I1(x3844), .I2(x3845), .I3(n8197), .I4(n8198), .O(n8203));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8204 (.I0(x3849), .I1(x3850), .I2(x3851), .I3(n8202), .I4(n8203), .O(n8204));
  LUT3 #(.INIT(8'hE8)) lut_n8205 (.I0(x3858), .I1(x3859), .I2(x3860), .O(n8205));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8206 (.I0(x3849), .I1(x3850), .I2(x3851), .I3(n8202), .I4(n8203), .O(n8206));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8207 (.I0(x3855), .I1(x3856), .I2(x3857), .I3(n8205), .I4(n8206), .O(n8207));
  LUT3 #(.INIT(8'h96)) lut_n8208 (.I0(n8196), .I1(n8199), .I2(n8200), .O(n8208));
  LUT3 #(.INIT(8'hE8)) lut_n8209 (.I0(n8204), .I1(n8207), .I2(n8208), .O(n8209));
  LUT3 #(.INIT(8'h96)) lut_n8210 (.I0(n8173), .I1(n8181), .I2(n8182), .O(n8210));
  LUT3 #(.INIT(8'hE8)) lut_n8211 (.I0(n8201), .I1(n8209), .I2(n8210), .O(n8211));
  LUT3 #(.INIT(8'hE8)) lut_n8212 (.I0(x3864), .I1(x3865), .I2(x3866), .O(n8212));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8213 (.I0(x3855), .I1(x3856), .I2(x3857), .I3(n8205), .I4(n8206), .O(n8213));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8214 (.I0(x3861), .I1(x3862), .I2(x3863), .I3(n8212), .I4(n8213), .O(n8214));
  LUT3 #(.INIT(8'hE8)) lut_n8215 (.I0(x3870), .I1(x3871), .I2(x3872), .O(n8215));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8216 (.I0(x3861), .I1(x3862), .I2(x3863), .I3(n8212), .I4(n8213), .O(n8216));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8217 (.I0(x3867), .I1(x3868), .I2(x3869), .I3(n8215), .I4(n8216), .O(n8217));
  LUT3 #(.INIT(8'h96)) lut_n8218 (.I0(n8204), .I1(n8207), .I2(n8208), .O(n8218));
  LUT3 #(.INIT(8'hE8)) lut_n8219 (.I0(n8214), .I1(n8217), .I2(n8218), .O(n8219));
  LUT3 #(.INIT(8'hE8)) lut_n8220 (.I0(x3876), .I1(x3877), .I2(x3878), .O(n8220));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8221 (.I0(x3867), .I1(x3868), .I2(x3869), .I3(n8215), .I4(n8216), .O(n8221));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8222 (.I0(x3873), .I1(x3874), .I2(x3875), .I3(n8220), .I4(n8221), .O(n8222));
  LUT3 #(.INIT(8'hE8)) lut_n8223 (.I0(x3882), .I1(x3883), .I2(x3884), .O(n8223));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8224 (.I0(x3873), .I1(x3874), .I2(x3875), .I3(n8220), .I4(n8221), .O(n8224));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8225 (.I0(x3879), .I1(x3880), .I2(x3881), .I3(n8223), .I4(n8224), .O(n8225));
  LUT3 #(.INIT(8'h96)) lut_n8226 (.I0(n8214), .I1(n8217), .I2(n8218), .O(n8226));
  LUT3 #(.INIT(8'hE8)) lut_n8227 (.I0(n8222), .I1(n8225), .I2(n8226), .O(n8227));
  LUT3 #(.INIT(8'h96)) lut_n8228 (.I0(n8201), .I1(n8209), .I2(n8210), .O(n8228));
  LUT3 #(.INIT(8'hE8)) lut_n8229 (.I0(n8219), .I1(n8227), .I2(n8228), .O(n8229));
  LUT3 #(.INIT(8'h96)) lut_n8230 (.I0(n8165), .I1(n8183), .I2(n8184), .O(n8230));
  LUT3 #(.INIT(8'hE8)) lut_n8231 (.I0(n8211), .I1(n8229), .I2(n8230), .O(n8231));
  LUT3 #(.INIT(8'hE8)) lut_n8232 (.I0(x3888), .I1(x3889), .I2(x3890), .O(n8232));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8233 (.I0(x3879), .I1(x3880), .I2(x3881), .I3(n8223), .I4(n8224), .O(n8233));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8234 (.I0(x3885), .I1(x3886), .I2(x3887), .I3(n8232), .I4(n8233), .O(n8234));
  LUT3 #(.INIT(8'hE8)) lut_n8235 (.I0(x3894), .I1(x3895), .I2(x3896), .O(n8235));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8236 (.I0(x3885), .I1(x3886), .I2(x3887), .I3(n8232), .I4(n8233), .O(n8236));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8237 (.I0(x3891), .I1(x3892), .I2(x3893), .I3(n8235), .I4(n8236), .O(n8237));
  LUT3 #(.INIT(8'h96)) lut_n8238 (.I0(n8222), .I1(n8225), .I2(n8226), .O(n8238));
  LUT3 #(.INIT(8'hE8)) lut_n8239 (.I0(n8234), .I1(n8237), .I2(n8238), .O(n8239));
  LUT3 #(.INIT(8'hE8)) lut_n8240 (.I0(x3900), .I1(x3901), .I2(x3902), .O(n8240));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8241 (.I0(x3891), .I1(x3892), .I2(x3893), .I3(n8235), .I4(n8236), .O(n8241));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8242 (.I0(x3897), .I1(x3898), .I2(x3899), .I3(n8240), .I4(n8241), .O(n8242));
  LUT3 #(.INIT(8'hE8)) lut_n8243 (.I0(x3906), .I1(x3907), .I2(x3908), .O(n8243));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8244 (.I0(x3897), .I1(x3898), .I2(x3899), .I3(n8240), .I4(n8241), .O(n8244));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8245 (.I0(x3903), .I1(x3904), .I2(x3905), .I3(n8243), .I4(n8244), .O(n8245));
  LUT3 #(.INIT(8'h96)) lut_n8246 (.I0(n8234), .I1(n8237), .I2(n8238), .O(n8246));
  LUT3 #(.INIT(8'hE8)) lut_n8247 (.I0(n8242), .I1(n8245), .I2(n8246), .O(n8247));
  LUT3 #(.INIT(8'h96)) lut_n8248 (.I0(n8219), .I1(n8227), .I2(n8228), .O(n8248));
  LUT3 #(.INIT(8'hE8)) lut_n8249 (.I0(n8239), .I1(n8247), .I2(n8248), .O(n8249));
  LUT3 #(.INIT(8'hE8)) lut_n8250 (.I0(x3912), .I1(x3913), .I2(x3914), .O(n8250));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8251 (.I0(x3903), .I1(x3904), .I2(x3905), .I3(n8243), .I4(n8244), .O(n8251));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8252 (.I0(x3909), .I1(x3910), .I2(x3911), .I3(n8250), .I4(n8251), .O(n8252));
  LUT3 #(.INIT(8'hE8)) lut_n8253 (.I0(x3918), .I1(x3919), .I2(x3920), .O(n8253));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8254 (.I0(x3909), .I1(x3910), .I2(x3911), .I3(n8250), .I4(n8251), .O(n8254));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8255 (.I0(x3915), .I1(x3916), .I2(x3917), .I3(n8253), .I4(n8254), .O(n8255));
  LUT3 #(.INIT(8'h96)) lut_n8256 (.I0(n8242), .I1(n8245), .I2(n8246), .O(n8256));
  LUT3 #(.INIT(8'hE8)) lut_n8257 (.I0(n8252), .I1(n8255), .I2(n8256), .O(n8257));
  LUT3 #(.INIT(8'hE8)) lut_n8258 (.I0(x3924), .I1(x3925), .I2(x3926), .O(n8258));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8259 (.I0(x3915), .I1(x3916), .I2(x3917), .I3(n8253), .I4(n8254), .O(n8259));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8260 (.I0(x3921), .I1(x3922), .I2(x3923), .I3(n8258), .I4(n8259), .O(n8260));
  LUT3 #(.INIT(8'hE8)) lut_n8261 (.I0(x3930), .I1(x3931), .I2(x3932), .O(n8261));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8262 (.I0(x3921), .I1(x3922), .I2(x3923), .I3(n8258), .I4(n8259), .O(n8262));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8263 (.I0(x3927), .I1(x3928), .I2(x3929), .I3(n8261), .I4(n8262), .O(n8263));
  LUT3 #(.INIT(8'h96)) lut_n8264 (.I0(n8252), .I1(n8255), .I2(n8256), .O(n8264));
  LUT3 #(.INIT(8'hE8)) lut_n8265 (.I0(n8260), .I1(n8263), .I2(n8264), .O(n8265));
  LUT3 #(.INIT(8'h96)) lut_n8266 (.I0(n8239), .I1(n8247), .I2(n8248), .O(n8266));
  LUT3 #(.INIT(8'hE8)) lut_n8267 (.I0(n8257), .I1(n8265), .I2(n8266), .O(n8267));
  LUT3 #(.INIT(8'h96)) lut_n8268 (.I0(n8211), .I1(n8229), .I2(n8230), .O(n8268));
  LUT3 #(.INIT(8'hE8)) lut_n8269 (.I0(n8249), .I1(n8267), .I2(n8268), .O(n8269));
  LUT3 #(.INIT(8'h96)) lut_n8270 (.I0(n8147), .I1(n8185), .I2(n8186), .O(n8270));
  LUT3 #(.INIT(8'hE8)) lut_n8271 (.I0(n8231), .I1(n8269), .I2(n8270), .O(n8271));
  LUT3 #(.INIT(8'hE8)) lut_n8272 (.I0(x3936), .I1(x3937), .I2(x3938), .O(n8272));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8273 (.I0(x3927), .I1(x3928), .I2(x3929), .I3(n8261), .I4(n8262), .O(n8273));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8274 (.I0(x3933), .I1(x3934), .I2(x3935), .I3(n8272), .I4(n8273), .O(n8274));
  LUT3 #(.INIT(8'hE8)) lut_n8275 (.I0(x3942), .I1(x3943), .I2(x3944), .O(n8275));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8276 (.I0(x3933), .I1(x3934), .I2(x3935), .I3(n8272), .I4(n8273), .O(n8276));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8277 (.I0(x3939), .I1(x3940), .I2(x3941), .I3(n8275), .I4(n8276), .O(n8277));
  LUT3 #(.INIT(8'h96)) lut_n8278 (.I0(n8260), .I1(n8263), .I2(n8264), .O(n8278));
  LUT3 #(.INIT(8'hE8)) lut_n8279 (.I0(n8274), .I1(n8277), .I2(n8278), .O(n8279));
  LUT3 #(.INIT(8'hE8)) lut_n8280 (.I0(x3948), .I1(x3949), .I2(x3950), .O(n8280));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8281 (.I0(x3939), .I1(x3940), .I2(x3941), .I3(n8275), .I4(n8276), .O(n8281));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8282 (.I0(x3945), .I1(x3946), .I2(x3947), .I3(n8280), .I4(n8281), .O(n8282));
  LUT3 #(.INIT(8'hE8)) lut_n8283 (.I0(x3954), .I1(x3955), .I2(x3956), .O(n8283));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8284 (.I0(x3945), .I1(x3946), .I2(x3947), .I3(n8280), .I4(n8281), .O(n8284));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8285 (.I0(x3951), .I1(x3952), .I2(x3953), .I3(n8283), .I4(n8284), .O(n8285));
  LUT3 #(.INIT(8'h96)) lut_n8286 (.I0(n8274), .I1(n8277), .I2(n8278), .O(n8286));
  LUT3 #(.INIT(8'hE8)) lut_n8287 (.I0(n8282), .I1(n8285), .I2(n8286), .O(n8287));
  LUT3 #(.INIT(8'h96)) lut_n8288 (.I0(n8257), .I1(n8265), .I2(n8266), .O(n8288));
  LUT3 #(.INIT(8'hE8)) lut_n8289 (.I0(n8279), .I1(n8287), .I2(n8288), .O(n8289));
  LUT3 #(.INIT(8'hE8)) lut_n8290 (.I0(x3960), .I1(x3961), .I2(x3962), .O(n8290));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8291 (.I0(x3951), .I1(x3952), .I2(x3953), .I3(n8283), .I4(n8284), .O(n8291));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8292 (.I0(x3957), .I1(x3958), .I2(x3959), .I3(n8290), .I4(n8291), .O(n8292));
  LUT3 #(.INIT(8'hE8)) lut_n8293 (.I0(x3966), .I1(x3967), .I2(x3968), .O(n8293));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8294 (.I0(x3957), .I1(x3958), .I2(x3959), .I3(n8290), .I4(n8291), .O(n8294));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8295 (.I0(x3963), .I1(x3964), .I2(x3965), .I3(n8293), .I4(n8294), .O(n8295));
  LUT3 #(.INIT(8'h96)) lut_n8296 (.I0(n8282), .I1(n8285), .I2(n8286), .O(n8296));
  LUT3 #(.INIT(8'hE8)) lut_n8297 (.I0(n8292), .I1(n8295), .I2(n8296), .O(n8297));
  LUT3 #(.INIT(8'hE8)) lut_n8298 (.I0(x3972), .I1(x3973), .I2(x3974), .O(n8298));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8299 (.I0(x3963), .I1(x3964), .I2(x3965), .I3(n8293), .I4(n8294), .O(n8299));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8300 (.I0(x3969), .I1(x3970), .I2(x3971), .I3(n8298), .I4(n8299), .O(n8300));
  LUT3 #(.INIT(8'hE8)) lut_n8301 (.I0(x3978), .I1(x3979), .I2(x3980), .O(n8301));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8302 (.I0(x3969), .I1(x3970), .I2(x3971), .I3(n8298), .I4(n8299), .O(n8302));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8303 (.I0(x3975), .I1(x3976), .I2(x3977), .I3(n8301), .I4(n8302), .O(n8303));
  LUT3 #(.INIT(8'h96)) lut_n8304 (.I0(n8292), .I1(n8295), .I2(n8296), .O(n8304));
  LUT3 #(.INIT(8'hE8)) lut_n8305 (.I0(n8300), .I1(n8303), .I2(n8304), .O(n8305));
  LUT3 #(.INIT(8'h96)) lut_n8306 (.I0(n8279), .I1(n8287), .I2(n8288), .O(n8306));
  LUT3 #(.INIT(8'hE8)) lut_n8307 (.I0(n8297), .I1(n8305), .I2(n8306), .O(n8307));
  LUT3 #(.INIT(8'h96)) lut_n8308 (.I0(n8249), .I1(n8267), .I2(n8268), .O(n8308));
  LUT3 #(.INIT(8'hE8)) lut_n8309 (.I0(n8289), .I1(n8307), .I2(n8308), .O(n8309));
  LUT3 #(.INIT(8'hE8)) lut_n8310 (.I0(x3984), .I1(x3985), .I2(x3986), .O(n8310));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8311 (.I0(x3975), .I1(x3976), .I2(x3977), .I3(n8301), .I4(n8302), .O(n8311));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8312 (.I0(x3981), .I1(x3982), .I2(x3983), .I3(n8310), .I4(n8311), .O(n8312));
  LUT3 #(.INIT(8'hE8)) lut_n8313 (.I0(x3990), .I1(x3991), .I2(x3992), .O(n8313));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8314 (.I0(x3981), .I1(x3982), .I2(x3983), .I3(n8310), .I4(n8311), .O(n8314));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8315 (.I0(x3987), .I1(x3988), .I2(x3989), .I3(n8313), .I4(n8314), .O(n8315));
  LUT3 #(.INIT(8'h96)) lut_n8316 (.I0(n8300), .I1(n8303), .I2(n8304), .O(n8316));
  LUT3 #(.INIT(8'hE8)) lut_n8317 (.I0(n8312), .I1(n8315), .I2(n8316), .O(n8317));
  LUT3 #(.INIT(8'hE8)) lut_n8318 (.I0(x3996), .I1(x3997), .I2(x3998), .O(n8318));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8319 (.I0(x3987), .I1(x3988), .I2(x3989), .I3(n8313), .I4(n8314), .O(n8319));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8320 (.I0(x3993), .I1(x3994), .I2(x3995), .I3(n8318), .I4(n8319), .O(n8320));
  LUT3 #(.INIT(8'hE8)) lut_n8321 (.I0(x4002), .I1(x4003), .I2(x4004), .O(n8321));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8322 (.I0(x3993), .I1(x3994), .I2(x3995), .I3(n8318), .I4(n8319), .O(n8322));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8323 (.I0(x3999), .I1(x4000), .I2(x4001), .I3(n8321), .I4(n8322), .O(n8323));
  LUT3 #(.INIT(8'h96)) lut_n8324 (.I0(n8312), .I1(n8315), .I2(n8316), .O(n8324));
  LUT3 #(.INIT(8'hE8)) lut_n8325 (.I0(n8320), .I1(n8323), .I2(n8324), .O(n8325));
  LUT3 #(.INIT(8'h96)) lut_n8326 (.I0(n8297), .I1(n8305), .I2(n8306), .O(n8326));
  LUT3 #(.INIT(8'hE8)) lut_n8327 (.I0(n8317), .I1(n8325), .I2(n8326), .O(n8327));
  LUT3 #(.INIT(8'hE8)) lut_n8328 (.I0(x4008), .I1(x4009), .I2(x4010), .O(n8328));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8329 (.I0(x3999), .I1(x4000), .I2(x4001), .I3(n8321), .I4(n8322), .O(n8329));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8330 (.I0(x4005), .I1(x4006), .I2(x4007), .I3(n8328), .I4(n8329), .O(n8330));
  LUT3 #(.INIT(8'hE8)) lut_n8331 (.I0(x4014), .I1(x4015), .I2(x4016), .O(n8331));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8332 (.I0(x4005), .I1(x4006), .I2(x4007), .I3(n8328), .I4(n8329), .O(n8332));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8333 (.I0(x4011), .I1(x4012), .I2(x4013), .I3(n8331), .I4(n8332), .O(n8333));
  LUT3 #(.INIT(8'h96)) lut_n8334 (.I0(n8320), .I1(n8323), .I2(n8324), .O(n8334));
  LUT3 #(.INIT(8'hE8)) lut_n8335 (.I0(n8330), .I1(n8333), .I2(n8334), .O(n8335));
  LUT3 #(.INIT(8'hE8)) lut_n8336 (.I0(x4020), .I1(x4021), .I2(x4022), .O(n8336));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8337 (.I0(x4011), .I1(x4012), .I2(x4013), .I3(n8331), .I4(n8332), .O(n8337));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8338 (.I0(x4017), .I1(x4018), .I2(x4019), .I3(n8336), .I4(n8337), .O(n8338));
  LUT3 #(.INIT(8'hE8)) lut_n8339 (.I0(x4026), .I1(x4027), .I2(x4028), .O(n8339));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8340 (.I0(x4017), .I1(x4018), .I2(x4019), .I3(n8336), .I4(n8337), .O(n8340));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8341 (.I0(x4023), .I1(x4024), .I2(x4025), .I3(n8339), .I4(n8340), .O(n8341));
  LUT3 #(.INIT(8'h96)) lut_n8342 (.I0(n8330), .I1(n8333), .I2(n8334), .O(n8342));
  LUT3 #(.INIT(8'hE8)) lut_n8343 (.I0(n8338), .I1(n8341), .I2(n8342), .O(n8343));
  LUT3 #(.INIT(8'h96)) lut_n8344 (.I0(n8317), .I1(n8325), .I2(n8326), .O(n8344));
  LUT3 #(.INIT(8'hE8)) lut_n8345 (.I0(n8335), .I1(n8343), .I2(n8344), .O(n8345));
  LUT3 #(.INIT(8'h96)) lut_n8346 (.I0(n8289), .I1(n8307), .I2(n8308), .O(n8346));
  LUT3 #(.INIT(8'hE8)) lut_n8347 (.I0(n8327), .I1(n8345), .I2(n8346), .O(n8347));
  LUT3 #(.INIT(8'h96)) lut_n8348 (.I0(n8231), .I1(n8269), .I2(n8270), .O(n8348));
  LUT3 #(.INIT(8'hE8)) lut_n8349 (.I0(n8309), .I1(n8347), .I2(n8348), .O(n8349));
  LUT3 #(.INIT(8'h96)) lut_n8350 (.I0(n8109), .I1(n8187), .I2(n8188), .O(n8350));
  LUT3 #(.INIT(8'hE8)) lut_n8351 (.I0(n8271), .I1(n8349), .I2(n8350), .O(n8351));
  LUT3 #(.INIT(8'hE8)) lut_n8352 (.I0(x4032), .I1(x4033), .I2(x4034), .O(n8352));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8353 (.I0(x4023), .I1(x4024), .I2(x4025), .I3(n8339), .I4(n8340), .O(n8353));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8354 (.I0(x4029), .I1(x4030), .I2(x4031), .I3(n8352), .I4(n8353), .O(n8354));
  LUT3 #(.INIT(8'hE8)) lut_n8355 (.I0(x4038), .I1(x4039), .I2(x4040), .O(n8355));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8356 (.I0(x4029), .I1(x4030), .I2(x4031), .I3(n8352), .I4(n8353), .O(n8356));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8357 (.I0(x4035), .I1(x4036), .I2(x4037), .I3(n8355), .I4(n8356), .O(n8357));
  LUT3 #(.INIT(8'h96)) lut_n8358 (.I0(n8338), .I1(n8341), .I2(n8342), .O(n8358));
  LUT3 #(.INIT(8'hE8)) lut_n8359 (.I0(n8354), .I1(n8357), .I2(n8358), .O(n8359));
  LUT3 #(.INIT(8'hE8)) lut_n8360 (.I0(x4044), .I1(x4045), .I2(x4046), .O(n8360));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8361 (.I0(x4035), .I1(x4036), .I2(x4037), .I3(n8355), .I4(n8356), .O(n8361));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8362 (.I0(x4041), .I1(x4042), .I2(x4043), .I3(n8360), .I4(n8361), .O(n8362));
  LUT3 #(.INIT(8'hE8)) lut_n8363 (.I0(x4050), .I1(x4051), .I2(x4052), .O(n8363));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8364 (.I0(x4041), .I1(x4042), .I2(x4043), .I3(n8360), .I4(n8361), .O(n8364));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8365 (.I0(x4047), .I1(x4048), .I2(x4049), .I3(n8363), .I4(n8364), .O(n8365));
  LUT3 #(.INIT(8'h96)) lut_n8366 (.I0(n8354), .I1(n8357), .I2(n8358), .O(n8366));
  LUT3 #(.INIT(8'hE8)) lut_n8367 (.I0(n8362), .I1(n8365), .I2(n8366), .O(n8367));
  LUT3 #(.INIT(8'h96)) lut_n8368 (.I0(n8335), .I1(n8343), .I2(n8344), .O(n8368));
  LUT3 #(.INIT(8'hE8)) lut_n8369 (.I0(n8359), .I1(n8367), .I2(n8368), .O(n8369));
  LUT3 #(.INIT(8'hE8)) lut_n8370 (.I0(x4056), .I1(x4057), .I2(x4058), .O(n8370));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8371 (.I0(x4047), .I1(x4048), .I2(x4049), .I3(n8363), .I4(n8364), .O(n8371));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8372 (.I0(x4053), .I1(x4054), .I2(x4055), .I3(n8370), .I4(n8371), .O(n8372));
  LUT3 #(.INIT(8'hE8)) lut_n8373 (.I0(x4062), .I1(x4063), .I2(x4064), .O(n8373));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8374 (.I0(x4053), .I1(x4054), .I2(x4055), .I3(n8370), .I4(n8371), .O(n8374));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8375 (.I0(x4059), .I1(x4060), .I2(x4061), .I3(n8373), .I4(n8374), .O(n8375));
  LUT3 #(.INIT(8'h96)) lut_n8376 (.I0(n8362), .I1(n8365), .I2(n8366), .O(n8376));
  LUT3 #(.INIT(8'hE8)) lut_n8377 (.I0(n8372), .I1(n8375), .I2(n8376), .O(n8377));
  LUT3 #(.INIT(8'hE8)) lut_n8378 (.I0(x4068), .I1(x4069), .I2(x4070), .O(n8378));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8379 (.I0(x4059), .I1(x4060), .I2(x4061), .I3(n8373), .I4(n8374), .O(n8379));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8380 (.I0(x4065), .I1(x4066), .I2(x4067), .I3(n8378), .I4(n8379), .O(n8380));
  LUT3 #(.INIT(8'hE8)) lut_n8381 (.I0(x4074), .I1(x4075), .I2(x4076), .O(n8381));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8382 (.I0(x4065), .I1(x4066), .I2(x4067), .I3(n8378), .I4(n8379), .O(n8382));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8383 (.I0(x4071), .I1(x4072), .I2(x4073), .I3(n8381), .I4(n8382), .O(n8383));
  LUT3 #(.INIT(8'h96)) lut_n8384 (.I0(n8372), .I1(n8375), .I2(n8376), .O(n8384));
  LUT3 #(.INIT(8'hE8)) lut_n8385 (.I0(n8380), .I1(n8383), .I2(n8384), .O(n8385));
  LUT3 #(.INIT(8'h96)) lut_n8386 (.I0(n8359), .I1(n8367), .I2(n8368), .O(n8386));
  LUT3 #(.INIT(8'hE8)) lut_n8387 (.I0(n8377), .I1(n8385), .I2(n8386), .O(n8387));
  LUT3 #(.INIT(8'h96)) lut_n8388 (.I0(n8327), .I1(n8345), .I2(n8346), .O(n8388));
  LUT3 #(.INIT(8'hE8)) lut_n8389 (.I0(n8369), .I1(n8387), .I2(n8388), .O(n8389));
  LUT3 #(.INIT(8'hE8)) lut_n8390 (.I0(x4080), .I1(x4081), .I2(x4082), .O(n8390));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8391 (.I0(x4071), .I1(x4072), .I2(x4073), .I3(n8381), .I4(n8382), .O(n8391));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8392 (.I0(x4077), .I1(x4078), .I2(x4079), .I3(n8390), .I4(n8391), .O(n8392));
  LUT3 #(.INIT(8'hE8)) lut_n8393 (.I0(x4086), .I1(x4087), .I2(x4088), .O(n8393));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8394 (.I0(x4077), .I1(x4078), .I2(x4079), .I3(n8390), .I4(n8391), .O(n8394));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8395 (.I0(x4083), .I1(x4084), .I2(x4085), .I3(n8393), .I4(n8394), .O(n8395));
  LUT3 #(.INIT(8'h96)) lut_n8396 (.I0(n8380), .I1(n8383), .I2(n8384), .O(n8396));
  LUT3 #(.INIT(8'hE8)) lut_n8397 (.I0(n8392), .I1(n8395), .I2(n8396), .O(n8397));
  LUT3 #(.INIT(8'hE8)) lut_n8398 (.I0(x4092), .I1(x4093), .I2(x4094), .O(n8398));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8399 (.I0(x4083), .I1(x4084), .I2(x4085), .I3(n8393), .I4(n8394), .O(n8399));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8400 (.I0(x4089), .I1(x4090), .I2(x4091), .I3(n8398), .I4(n8399), .O(n8400));
  LUT3 #(.INIT(8'hE8)) lut_n8401 (.I0(x4098), .I1(x4099), .I2(x4100), .O(n8401));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8402 (.I0(x4089), .I1(x4090), .I2(x4091), .I3(n8398), .I4(n8399), .O(n8402));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8403 (.I0(x4095), .I1(x4096), .I2(x4097), .I3(n8401), .I4(n8402), .O(n8403));
  LUT3 #(.INIT(8'h96)) lut_n8404 (.I0(n8392), .I1(n8395), .I2(n8396), .O(n8404));
  LUT3 #(.INIT(8'hE8)) lut_n8405 (.I0(n8400), .I1(n8403), .I2(n8404), .O(n8405));
  LUT3 #(.INIT(8'h96)) lut_n8406 (.I0(n8377), .I1(n8385), .I2(n8386), .O(n8406));
  LUT3 #(.INIT(8'hE8)) lut_n8407 (.I0(n8397), .I1(n8405), .I2(n8406), .O(n8407));
  LUT3 #(.INIT(8'hE8)) lut_n8408 (.I0(x4104), .I1(x4105), .I2(x4106), .O(n8408));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8409 (.I0(x4095), .I1(x4096), .I2(x4097), .I3(n8401), .I4(n8402), .O(n8409));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8410 (.I0(x4101), .I1(x4102), .I2(x4103), .I3(n8408), .I4(n8409), .O(n8410));
  LUT3 #(.INIT(8'hE8)) lut_n8411 (.I0(x4110), .I1(x4111), .I2(x4112), .O(n8411));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8412 (.I0(x4101), .I1(x4102), .I2(x4103), .I3(n8408), .I4(n8409), .O(n8412));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8413 (.I0(x4107), .I1(x4108), .I2(x4109), .I3(n8411), .I4(n8412), .O(n8413));
  LUT3 #(.INIT(8'h96)) lut_n8414 (.I0(n8400), .I1(n8403), .I2(n8404), .O(n8414));
  LUT3 #(.INIT(8'hE8)) lut_n8415 (.I0(n8410), .I1(n8413), .I2(n8414), .O(n8415));
  LUT3 #(.INIT(8'hE8)) lut_n8416 (.I0(x4116), .I1(x4117), .I2(x4118), .O(n8416));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8417 (.I0(x4107), .I1(x4108), .I2(x4109), .I3(n8411), .I4(n8412), .O(n8417));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8418 (.I0(x4113), .I1(x4114), .I2(x4115), .I3(n8416), .I4(n8417), .O(n8418));
  LUT3 #(.INIT(8'hE8)) lut_n8419 (.I0(x4122), .I1(x4123), .I2(x4124), .O(n8419));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8420 (.I0(x4113), .I1(x4114), .I2(x4115), .I3(n8416), .I4(n8417), .O(n8420));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8421 (.I0(x4119), .I1(x4120), .I2(x4121), .I3(n8419), .I4(n8420), .O(n8421));
  LUT3 #(.INIT(8'h96)) lut_n8422 (.I0(n8410), .I1(n8413), .I2(n8414), .O(n8422));
  LUT3 #(.INIT(8'hE8)) lut_n8423 (.I0(n8418), .I1(n8421), .I2(n8422), .O(n8423));
  LUT3 #(.INIT(8'h96)) lut_n8424 (.I0(n8397), .I1(n8405), .I2(n8406), .O(n8424));
  LUT3 #(.INIT(8'hE8)) lut_n8425 (.I0(n8415), .I1(n8423), .I2(n8424), .O(n8425));
  LUT3 #(.INIT(8'h96)) lut_n8426 (.I0(n8369), .I1(n8387), .I2(n8388), .O(n8426));
  LUT3 #(.INIT(8'hE8)) lut_n8427 (.I0(n8407), .I1(n8425), .I2(n8426), .O(n8427));
  LUT3 #(.INIT(8'h96)) lut_n8428 (.I0(n8309), .I1(n8347), .I2(n8348), .O(n8428));
  LUT3 #(.INIT(8'hE8)) lut_n8429 (.I0(n8389), .I1(n8427), .I2(n8428), .O(n8429));
  LUT3 #(.INIT(8'hE8)) lut_n8430 (.I0(x4128), .I1(x4129), .I2(x4130), .O(n8430));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8431 (.I0(x4119), .I1(x4120), .I2(x4121), .I3(n8419), .I4(n8420), .O(n8431));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8432 (.I0(x4125), .I1(x4126), .I2(x4127), .I3(n8430), .I4(n8431), .O(n8432));
  LUT3 #(.INIT(8'hE8)) lut_n8433 (.I0(x4134), .I1(x4135), .I2(x4136), .O(n8433));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8434 (.I0(x4125), .I1(x4126), .I2(x4127), .I3(n8430), .I4(n8431), .O(n8434));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8435 (.I0(x4131), .I1(x4132), .I2(x4133), .I3(n8433), .I4(n8434), .O(n8435));
  LUT3 #(.INIT(8'h96)) lut_n8436 (.I0(n8418), .I1(n8421), .I2(n8422), .O(n8436));
  LUT3 #(.INIT(8'hE8)) lut_n8437 (.I0(n8432), .I1(n8435), .I2(n8436), .O(n8437));
  LUT3 #(.INIT(8'hE8)) lut_n8438 (.I0(x4140), .I1(x4141), .I2(x4142), .O(n8438));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8439 (.I0(x4131), .I1(x4132), .I2(x4133), .I3(n8433), .I4(n8434), .O(n8439));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8440 (.I0(x4137), .I1(x4138), .I2(x4139), .I3(n8438), .I4(n8439), .O(n8440));
  LUT3 #(.INIT(8'hE8)) lut_n8441 (.I0(x4146), .I1(x4147), .I2(x4148), .O(n8441));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8442 (.I0(x4137), .I1(x4138), .I2(x4139), .I3(n8438), .I4(n8439), .O(n8442));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8443 (.I0(x4143), .I1(x4144), .I2(x4145), .I3(n8441), .I4(n8442), .O(n8443));
  LUT3 #(.INIT(8'h96)) lut_n8444 (.I0(n8432), .I1(n8435), .I2(n8436), .O(n8444));
  LUT3 #(.INIT(8'hE8)) lut_n8445 (.I0(n8440), .I1(n8443), .I2(n8444), .O(n8445));
  LUT3 #(.INIT(8'h96)) lut_n8446 (.I0(n8415), .I1(n8423), .I2(n8424), .O(n8446));
  LUT3 #(.INIT(8'hE8)) lut_n8447 (.I0(n8437), .I1(n8445), .I2(n8446), .O(n8447));
  LUT3 #(.INIT(8'hE8)) lut_n8448 (.I0(x4152), .I1(x4153), .I2(x4154), .O(n8448));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8449 (.I0(x4143), .I1(x4144), .I2(x4145), .I3(n8441), .I4(n8442), .O(n8449));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8450 (.I0(x4149), .I1(x4150), .I2(x4151), .I3(n8448), .I4(n8449), .O(n8450));
  LUT3 #(.INIT(8'hE8)) lut_n8451 (.I0(x4158), .I1(x4159), .I2(x4160), .O(n8451));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8452 (.I0(x4149), .I1(x4150), .I2(x4151), .I3(n8448), .I4(n8449), .O(n8452));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8453 (.I0(x4155), .I1(x4156), .I2(x4157), .I3(n8451), .I4(n8452), .O(n8453));
  LUT3 #(.INIT(8'h96)) lut_n8454 (.I0(n8440), .I1(n8443), .I2(n8444), .O(n8454));
  LUT3 #(.INIT(8'hE8)) lut_n8455 (.I0(n8450), .I1(n8453), .I2(n8454), .O(n8455));
  LUT3 #(.INIT(8'hE8)) lut_n8456 (.I0(x4164), .I1(x4165), .I2(x4166), .O(n8456));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8457 (.I0(x4155), .I1(x4156), .I2(x4157), .I3(n8451), .I4(n8452), .O(n8457));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8458 (.I0(x4161), .I1(x4162), .I2(x4163), .I3(n8456), .I4(n8457), .O(n8458));
  LUT3 #(.INIT(8'hE8)) lut_n8459 (.I0(x4170), .I1(x4171), .I2(x4172), .O(n8459));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8460 (.I0(x4161), .I1(x4162), .I2(x4163), .I3(n8456), .I4(n8457), .O(n8460));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8461 (.I0(x4167), .I1(x4168), .I2(x4169), .I3(n8459), .I4(n8460), .O(n8461));
  LUT3 #(.INIT(8'h96)) lut_n8462 (.I0(n8450), .I1(n8453), .I2(n8454), .O(n8462));
  LUT3 #(.INIT(8'hE8)) lut_n8463 (.I0(n8458), .I1(n8461), .I2(n8462), .O(n8463));
  LUT3 #(.INIT(8'h96)) lut_n8464 (.I0(n8437), .I1(n8445), .I2(n8446), .O(n8464));
  LUT3 #(.INIT(8'hE8)) lut_n8465 (.I0(n8455), .I1(n8463), .I2(n8464), .O(n8465));
  LUT3 #(.INIT(8'h96)) lut_n8466 (.I0(n8407), .I1(n8425), .I2(n8426), .O(n8466));
  LUT3 #(.INIT(8'hE8)) lut_n8467 (.I0(n8447), .I1(n8465), .I2(n8466), .O(n8467));
  LUT3 #(.INIT(8'hE8)) lut_n8468 (.I0(x4176), .I1(x4177), .I2(x4178), .O(n8468));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8469 (.I0(x4167), .I1(x4168), .I2(x4169), .I3(n8459), .I4(n8460), .O(n8469));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8470 (.I0(x4173), .I1(x4174), .I2(x4175), .I3(n8468), .I4(n8469), .O(n8470));
  LUT3 #(.INIT(8'hE8)) lut_n8471 (.I0(x4182), .I1(x4183), .I2(x4184), .O(n8471));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8472 (.I0(x4173), .I1(x4174), .I2(x4175), .I3(n8468), .I4(n8469), .O(n8472));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8473 (.I0(x4179), .I1(x4180), .I2(x4181), .I3(n8471), .I4(n8472), .O(n8473));
  LUT3 #(.INIT(8'h96)) lut_n8474 (.I0(n8458), .I1(n8461), .I2(n8462), .O(n8474));
  LUT3 #(.INIT(8'hE8)) lut_n8475 (.I0(n8470), .I1(n8473), .I2(n8474), .O(n8475));
  LUT3 #(.INIT(8'hE8)) lut_n8476 (.I0(x4188), .I1(x4189), .I2(x4190), .O(n8476));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8477 (.I0(x4179), .I1(x4180), .I2(x4181), .I3(n8471), .I4(n8472), .O(n8477));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8478 (.I0(x4185), .I1(x4186), .I2(x4187), .I3(n8476), .I4(n8477), .O(n8478));
  LUT3 #(.INIT(8'hE8)) lut_n8479 (.I0(x4194), .I1(x4195), .I2(x4196), .O(n8479));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8480 (.I0(x4185), .I1(x4186), .I2(x4187), .I3(n8476), .I4(n8477), .O(n8480));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8481 (.I0(x4191), .I1(x4192), .I2(x4193), .I3(n8479), .I4(n8480), .O(n8481));
  LUT3 #(.INIT(8'h96)) lut_n8482 (.I0(n8470), .I1(n8473), .I2(n8474), .O(n8482));
  LUT3 #(.INIT(8'hE8)) lut_n8483 (.I0(n8478), .I1(n8481), .I2(n8482), .O(n8483));
  LUT3 #(.INIT(8'h96)) lut_n8484 (.I0(n8455), .I1(n8463), .I2(n8464), .O(n8484));
  LUT3 #(.INIT(8'hE8)) lut_n8485 (.I0(n8475), .I1(n8483), .I2(n8484), .O(n8485));
  LUT3 #(.INIT(8'hE8)) lut_n8486 (.I0(x4200), .I1(x4201), .I2(x4202), .O(n8486));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8487 (.I0(x4191), .I1(x4192), .I2(x4193), .I3(n8479), .I4(n8480), .O(n8487));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8488 (.I0(x4197), .I1(x4198), .I2(x4199), .I3(n8486), .I4(n8487), .O(n8488));
  LUT3 #(.INIT(8'hE8)) lut_n8489 (.I0(x4206), .I1(x4207), .I2(x4208), .O(n8489));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8490 (.I0(x4197), .I1(x4198), .I2(x4199), .I3(n8486), .I4(n8487), .O(n8490));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8491 (.I0(x4203), .I1(x4204), .I2(x4205), .I3(n8489), .I4(n8490), .O(n8491));
  LUT3 #(.INIT(8'h96)) lut_n8492 (.I0(n8478), .I1(n8481), .I2(n8482), .O(n8492));
  LUT3 #(.INIT(8'hE8)) lut_n8493 (.I0(n8488), .I1(n8491), .I2(n8492), .O(n8493));
  LUT3 #(.INIT(8'hE8)) lut_n8494 (.I0(x4212), .I1(x4213), .I2(x4214), .O(n8494));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8495 (.I0(x4203), .I1(x4204), .I2(x4205), .I3(n8489), .I4(n8490), .O(n8495));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8496 (.I0(x4209), .I1(x4210), .I2(x4211), .I3(n8494), .I4(n8495), .O(n8496));
  LUT3 #(.INIT(8'hE8)) lut_n8497 (.I0(x4218), .I1(x4219), .I2(x4220), .O(n8497));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8498 (.I0(x4209), .I1(x4210), .I2(x4211), .I3(n8494), .I4(n8495), .O(n8498));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8499 (.I0(x4215), .I1(x4216), .I2(x4217), .I3(n8497), .I4(n8498), .O(n8499));
  LUT3 #(.INIT(8'h96)) lut_n8500 (.I0(n8488), .I1(n8491), .I2(n8492), .O(n8500));
  LUT3 #(.INIT(8'hE8)) lut_n8501 (.I0(n8496), .I1(n8499), .I2(n8500), .O(n8501));
  LUT3 #(.INIT(8'h96)) lut_n8502 (.I0(n8475), .I1(n8483), .I2(n8484), .O(n8502));
  LUT3 #(.INIT(8'hE8)) lut_n8503 (.I0(n8493), .I1(n8501), .I2(n8502), .O(n8503));
  LUT3 #(.INIT(8'h96)) lut_n8504 (.I0(n8447), .I1(n8465), .I2(n8466), .O(n8504));
  LUT3 #(.INIT(8'hE8)) lut_n8505 (.I0(n8485), .I1(n8503), .I2(n8504), .O(n8505));
  LUT3 #(.INIT(8'h96)) lut_n8506 (.I0(n8389), .I1(n8427), .I2(n8428), .O(n8506));
  LUT3 #(.INIT(8'hE8)) lut_n8507 (.I0(n8467), .I1(n8505), .I2(n8506), .O(n8507));
  LUT3 #(.INIT(8'h96)) lut_n8508 (.I0(n8271), .I1(n8349), .I2(n8350), .O(n8508));
  LUT3 #(.INIT(8'hE8)) lut_n8509 (.I0(n8429), .I1(n8507), .I2(n8508), .O(n8509));
  LUT3 #(.INIT(8'h96)) lut_n8510 (.I0(n8031), .I1(n8189), .I2(n8190), .O(n8510));
  LUT3 #(.INIT(8'hE8)) lut_n8511 (.I0(n8351), .I1(n8509), .I2(n8510), .O(n8511));
  LUT3 #(.INIT(8'hE8)) lut_n8512 (.I0(x4224), .I1(x4225), .I2(x4226), .O(n8512));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8513 (.I0(x4215), .I1(x4216), .I2(x4217), .I3(n8497), .I4(n8498), .O(n8513));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8514 (.I0(x4221), .I1(x4222), .I2(x4223), .I3(n8512), .I4(n8513), .O(n8514));
  LUT3 #(.INIT(8'hE8)) lut_n8515 (.I0(x4230), .I1(x4231), .I2(x4232), .O(n8515));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8516 (.I0(x4221), .I1(x4222), .I2(x4223), .I3(n8512), .I4(n8513), .O(n8516));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8517 (.I0(x4227), .I1(x4228), .I2(x4229), .I3(n8515), .I4(n8516), .O(n8517));
  LUT3 #(.INIT(8'h96)) lut_n8518 (.I0(n8496), .I1(n8499), .I2(n8500), .O(n8518));
  LUT3 #(.INIT(8'hE8)) lut_n8519 (.I0(n8514), .I1(n8517), .I2(n8518), .O(n8519));
  LUT3 #(.INIT(8'hE8)) lut_n8520 (.I0(x4236), .I1(x4237), .I2(x4238), .O(n8520));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8521 (.I0(x4227), .I1(x4228), .I2(x4229), .I3(n8515), .I4(n8516), .O(n8521));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8522 (.I0(x4233), .I1(x4234), .I2(x4235), .I3(n8520), .I4(n8521), .O(n8522));
  LUT3 #(.INIT(8'hE8)) lut_n8523 (.I0(x4242), .I1(x4243), .I2(x4244), .O(n8523));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8524 (.I0(x4233), .I1(x4234), .I2(x4235), .I3(n8520), .I4(n8521), .O(n8524));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8525 (.I0(x4239), .I1(x4240), .I2(x4241), .I3(n8523), .I4(n8524), .O(n8525));
  LUT3 #(.INIT(8'h96)) lut_n8526 (.I0(n8514), .I1(n8517), .I2(n8518), .O(n8526));
  LUT3 #(.INIT(8'hE8)) lut_n8527 (.I0(n8522), .I1(n8525), .I2(n8526), .O(n8527));
  LUT3 #(.INIT(8'h96)) lut_n8528 (.I0(n8493), .I1(n8501), .I2(n8502), .O(n8528));
  LUT3 #(.INIT(8'hE8)) lut_n8529 (.I0(n8519), .I1(n8527), .I2(n8528), .O(n8529));
  LUT3 #(.INIT(8'hE8)) lut_n8530 (.I0(x4248), .I1(x4249), .I2(x4250), .O(n8530));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8531 (.I0(x4239), .I1(x4240), .I2(x4241), .I3(n8523), .I4(n8524), .O(n8531));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8532 (.I0(x4245), .I1(x4246), .I2(x4247), .I3(n8530), .I4(n8531), .O(n8532));
  LUT3 #(.INIT(8'hE8)) lut_n8533 (.I0(x4254), .I1(x4255), .I2(x4256), .O(n8533));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8534 (.I0(x4245), .I1(x4246), .I2(x4247), .I3(n8530), .I4(n8531), .O(n8534));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8535 (.I0(x4251), .I1(x4252), .I2(x4253), .I3(n8533), .I4(n8534), .O(n8535));
  LUT3 #(.INIT(8'h96)) lut_n8536 (.I0(n8522), .I1(n8525), .I2(n8526), .O(n8536));
  LUT3 #(.INIT(8'hE8)) lut_n8537 (.I0(n8532), .I1(n8535), .I2(n8536), .O(n8537));
  LUT3 #(.INIT(8'hE8)) lut_n8538 (.I0(x4260), .I1(x4261), .I2(x4262), .O(n8538));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8539 (.I0(x4251), .I1(x4252), .I2(x4253), .I3(n8533), .I4(n8534), .O(n8539));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8540 (.I0(x4257), .I1(x4258), .I2(x4259), .I3(n8538), .I4(n8539), .O(n8540));
  LUT3 #(.INIT(8'hE8)) lut_n8541 (.I0(x4266), .I1(x4267), .I2(x4268), .O(n8541));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8542 (.I0(x4257), .I1(x4258), .I2(x4259), .I3(n8538), .I4(n8539), .O(n8542));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8543 (.I0(x4263), .I1(x4264), .I2(x4265), .I3(n8541), .I4(n8542), .O(n8543));
  LUT3 #(.INIT(8'h96)) lut_n8544 (.I0(n8532), .I1(n8535), .I2(n8536), .O(n8544));
  LUT3 #(.INIT(8'hE8)) lut_n8545 (.I0(n8540), .I1(n8543), .I2(n8544), .O(n8545));
  LUT3 #(.INIT(8'h96)) lut_n8546 (.I0(n8519), .I1(n8527), .I2(n8528), .O(n8546));
  LUT3 #(.INIT(8'hE8)) lut_n8547 (.I0(n8537), .I1(n8545), .I2(n8546), .O(n8547));
  LUT3 #(.INIT(8'h96)) lut_n8548 (.I0(n8485), .I1(n8503), .I2(n8504), .O(n8548));
  LUT3 #(.INIT(8'hE8)) lut_n8549 (.I0(n8529), .I1(n8547), .I2(n8548), .O(n8549));
  LUT3 #(.INIT(8'hE8)) lut_n8550 (.I0(x4272), .I1(x4273), .I2(x4274), .O(n8550));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8551 (.I0(x4263), .I1(x4264), .I2(x4265), .I3(n8541), .I4(n8542), .O(n8551));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8552 (.I0(x4269), .I1(x4270), .I2(x4271), .I3(n8550), .I4(n8551), .O(n8552));
  LUT3 #(.INIT(8'hE8)) lut_n8553 (.I0(x4278), .I1(x4279), .I2(x4280), .O(n8553));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8554 (.I0(x4269), .I1(x4270), .I2(x4271), .I3(n8550), .I4(n8551), .O(n8554));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8555 (.I0(x4275), .I1(x4276), .I2(x4277), .I3(n8553), .I4(n8554), .O(n8555));
  LUT3 #(.INIT(8'h96)) lut_n8556 (.I0(n8540), .I1(n8543), .I2(n8544), .O(n8556));
  LUT3 #(.INIT(8'hE8)) lut_n8557 (.I0(n8552), .I1(n8555), .I2(n8556), .O(n8557));
  LUT3 #(.INIT(8'hE8)) lut_n8558 (.I0(x4284), .I1(x4285), .I2(x4286), .O(n8558));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8559 (.I0(x4275), .I1(x4276), .I2(x4277), .I3(n8553), .I4(n8554), .O(n8559));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8560 (.I0(x4281), .I1(x4282), .I2(x4283), .I3(n8558), .I4(n8559), .O(n8560));
  LUT3 #(.INIT(8'hE8)) lut_n8561 (.I0(x4290), .I1(x4291), .I2(x4292), .O(n8561));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8562 (.I0(x4281), .I1(x4282), .I2(x4283), .I3(n8558), .I4(n8559), .O(n8562));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8563 (.I0(x4287), .I1(x4288), .I2(x4289), .I3(n8561), .I4(n8562), .O(n8563));
  LUT3 #(.INIT(8'h96)) lut_n8564 (.I0(n8552), .I1(n8555), .I2(n8556), .O(n8564));
  LUT3 #(.INIT(8'hE8)) lut_n8565 (.I0(n8560), .I1(n8563), .I2(n8564), .O(n8565));
  LUT3 #(.INIT(8'h96)) lut_n8566 (.I0(n8537), .I1(n8545), .I2(n8546), .O(n8566));
  LUT3 #(.INIT(8'hE8)) lut_n8567 (.I0(n8557), .I1(n8565), .I2(n8566), .O(n8567));
  LUT3 #(.INIT(8'hE8)) lut_n8568 (.I0(x4296), .I1(x4297), .I2(x4298), .O(n8568));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8569 (.I0(x4287), .I1(x4288), .I2(x4289), .I3(n8561), .I4(n8562), .O(n8569));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8570 (.I0(x4293), .I1(x4294), .I2(x4295), .I3(n8568), .I4(n8569), .O(n8570));
  LUT3 #(.INIT(8'hE8)) lut_n8571 (.I0(x4302), .I1(x4303), .I2(x4304), .O(n8571));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8572 (.I0(x4293), .I1(x4294), .I2(x4295), .I3(n8568), .I4(n8569), .O(n8572));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8573 (.I0(x4299), .I1(x4300), .I2(x4301), .I3(n8571), .I4(n8572), .O(n8573));
  LUT3 #(.INIT(8'h96)) lut_n8574 (.I0(n8560), .I1(n8563), .I2(n8564), .O(n8574));
  LUT3 #(.INIT(8'hE8)) lut_n8575 (.I0(n8570), .I1(n8573), .I2(n8574), .O(n8575));
  LUT3 #(.INIT(8'hE8)) lut_n8576 (.I0(x4308), .I1(x4309), .I2(x4310), .O(n8576));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8577 (.I0(x4299), .I1(x4300), .I2(x4301), .I3(n8571), .I4(n8572), .O(n8577));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8578 (.I0(x4305), .I1(x4306), .I2(x4307), .I3(n8576), .I4(n8577), .O(n8578));
  LUT3 #(.INIT(8'hE8)) lut_n8579 (.I0(x4314), .I1(x4315), .I2(x4316), .O(n8579));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8580 (.I0(x4305), .I1(x4306), .I2(x4307), .I3(n8576), .I4(n8577), .O(n8580));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8581 (.I0(x4311), .I1(x4312), .I2(x4313), .I3(n8579), .I4(n8580), .O(n8581));
  LUT3 #(.INIT(8'h96)) lut_n8582 (.I0(n8570), .I1(n8573), .I2(n8574), .O(n8582));
  LUT3 #(.INIT(8'hE8)) lut_n8583 (.I0(n8578), .I1(n8581), .I2(n8582), .O(n8583));
  LUT3 #(.INIT(8'h96)) lut_n8584 (.I0(n8557), .I1(n8565), .I2(n8566), .O(n8584));
  LUT3 #(.INIT(8'hE8)) lut_n8585 (.I0(n8575), .I1(n8583), .I2(n8584), .O(n8585));
  LUT3 #(.INIT(8'h96)) lut_n8586 (.I0(n8529), .I1(n8547), .I2(n8548), .O(n8586));
  LUT3 #(.INIT(8'hE8)) lut_n8587 (.I0(n8567), .I1(n8585), .I2(n8586), .O(n8587));
  LUT3 #(.INIT(8'h96)) lut_n8588 (.I0(n8467), .I1(n8505), .I2(n8506), .O(n8588));
  LUT3 #(.INIT(8'hE8)) lut_n8589 (.I0(n8549), .I1(n8587), .I2(n8588), .O(n8589));
  LUT3 #(.INIT(8'hE8)) lut_n8590 (.I0(x4320), .I1(x4321), .I2(x4322), .O(n8590));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8591 (.I0(x4311), .I1(x4312), .I2(x4313), .I3(n8579), .I4(n8580), .O(n8591));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8592 (.I0(x4317), .I1(x4318), .I2(x4319), .I3(n8590), .I4(n8591), .O(n8592));
  LUT3 #(.INIT(8'hE8)) lut_n8593 (.I0(x4326), .I1(x4327), .I2(x4328), .O(n8593));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8594 (.I0(x4317), .I1(x4318), .I2(x4319), .I3(n8590), .I4(n8591), .O(n8594));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8595 (.I0(x4323), .I1(x4324), .I2(x4325), .I3(n8593), .I4(n8594), .O(n8595));
  LUT3 #(.INIT(8'h96)) lut_n8596 (.I0(n8578), .I1(n8581), .I2(n8582), .O(n8596));
  LUT3 #(.INIT(8'hE8)) lut_n8597 (.I0(n8592), .I1(n8595), .I2(n8596), .O(n8597));
  LUT3 #(.INIT(8'hE8)) lut_n8598 (.I0(x4332), .I1(x4333), .I2(x4334), .O(n8598));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8599 (.I0(x4323), .I1(x4324), .I2(x4325), .I3(n8593), .I4(n8594), .O(n8599));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8600 (.I0(x4329), .I1(x4330), .I2(x4331), .I3(n8598), .I4(n8599), .O(n8600));
  LUT3 #(.INIT(8'hE8)) lut_n8601 (.I0(x4338), .I1(x4339), .I2(x4340), .O(n8601));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8602 (.I0(x4329), .I1(x4330), .I2(x4331), .I3(n8598), .I4(n8599), .O(n8602));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8603 (.I0(x4335), .I1(x4336), .I2(x4337), .I3(n8601), .I4(n8602), .O(n8603));
  LUT3 #(.INIT(8'h96)) lut_n8604 (.I0(n8592), .I1(n8595), .I2(n8596), .O(n8604));
  LUT3 #(.INIT(8'hE8)) lut_n8605 (.I0(n8600), .I1(n8603), .I2(n8604), .O(n8605));
  LUT3 #(.INIT(8'h96)) lut_n8606 (.I0(n8575), .I1(n8583), .I2(n8584), .O(n8606));
  LUT3 #(.INIT(8'hE8)) lut_n8607 (.I0(n8597), .I1(n8605), .I2(n8606), .O(n8607));
  LUT3 #(.INIT(8'hE8)) lut_n8608 (.I0(x4344), .I1(x4345), .I2(x4346), .O(n8608));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8609 (.I0(x4335), .I1(x4336), .I2(x4337), .I3(n8601), .I4(n8602), .O(n8609));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8610 (.I0(x4341), .I1(x4342), .I2(x4343), .I3(n8608), .I4(n8609), .O(n8610));
  LUT3 #(.INIT(8'hE8)) lut_n8611 (.I0(x4350), .I1(x4351), .I2(x4352), .O(n8611));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8612 (.I0(x4341), .I1(x4342), .I2(x4343), .I3(n8608), .I4(n8609), .O(n8612));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8613 (.I0(x4347), .I1(x4348), .I2(x4349), .I3(n8611), .I4(n8612), .O(n8613));
  LUT3 #(.INIT(8'h96)) lut_n8614 (.I0(n8600), .I1(n8603), .I2(n8604), .O(n8614));
  LUT3 #(.INIT(8'hE8)) lut_n8615 (.I0(n8610), .I1(n8613), .I2(n8614), .O(n8615));
  LUT3 #(.INIT(8'hE8)) lut_n8616 (.I0(x4356), .I1(x4357), .I2(x4358), .O(n8616));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8617 (.I0(x4347), .I1(x4348), .I2(x4349), .I3(n8611), .I4(n8612), .O(n8617));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8618 (.I0(x4353), .I1(x4354), .I2(x4355), .I3(n8616), .I4(n8617), .O(n8618));
  LUT3 #(.INIT(8'hE8)) lut_n8619 (.I0(x4362), .I1(x4363), .I2(x4364), .O(n8619));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8620 (.I0(x4353), .I1(x4354), .I2(x4355), .I3(n8616), .I4(n8617), .O(n8620));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8621 (.I0(x4359), .I1(x4360), .I2(x4361), .I3(n8619), .I4(n8620), .O(n8621));
  LUT3 #(.INIT(8'h96)) lut_n8622 (.I0(n8610), .I1(n8613), .I2(n8614), .O(n8622));
  LUT3 #(.INIT(8'hE8)) lut_n8623 (.I0(n8618), .I1(n8621), .I2(n8622), .O(n8623));
  LUT3 #(.INIT(8'h96)) lut_n8624 (.I0(n8597), .I1(n8605), .I2(n8606), .O(n8624));
  LUT3 #(.INIT(8'hE8)) lut_n8625 (.I0(n8615), .I1(n8623), .I2(n8624), .O(n8625));
  LUT3 #(.INIT(8'h96)) lut_n8626 (.I0(n8567), .I1(n8585), .I2(n8586), .O(n8626));
  LUT3 #(.INIT(8'hE8)) lut_n8627 (.I0(n8607), .I1(n8625), .I2(n8626), .O(n8627));
  LUT3 #(.INIT(8'hE8)) lut_n8628 (.I0(x4368), .I1(x4369), .I2(x4370), .O(n8628));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8629 (.I0(x4359), .I1(x4360), .I2(x4361), .I3(n8619), .I4(n8620), .O(n8629));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8630 (.I0(x4365), .I1(x4366), .I2(x4367), .I3(n8628), .I4(n8629), .O(n8630));
  LUT3 #(.INIT(8'hE8)) lut_n8631 (.I0(x4374), .I1(x4375), .I2(x4376), .O(n8631));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8632 (.I0(x4365), .I1(x4366), .I2(x4367), .I3(n8628), .I4(n8629), .O(n8632));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8633 (.I0(x4371), .I1(x4372), .I2(x4373), .I3(n8631), .I4(n8632), .O(n8633));
  LUT3 #(.INIT(8'h96)) lut_n8634 (.I0(n8618), .I1(n8621), .I2(n8622), .O(n8634));
  LUT3 #(.INIT(8'hE8)) lut_n8635 (.I0(n8630), .I1(n8633), .I2(n8634), .O(n8635));
  LUT3 #(.INIT(8'hE8)) lut_n8636 (.I0(x4380), .I1(x4381), .I2(x4382), .O(n8636));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8637 (.I0(x4371), .I1(x4372), .I2(x4373), .I3(n8631), .I4(n8632), .O(n8637));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8638 (.I0(x4377), .I1(x4378), .I2(x4379), .I3(n8636), .I4(n8637), .O(n8638));
  LUT3 #(.INIT(8'hE8)) lut_n8639 (.I0(x4386), .I1(x4387), .I2(x4388), .O(n8639));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8640 (.I0(x4377), .I1(x4378), .I2(x4379), .I3(n8636), .I4(n8637), .O(n8640));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8641 (.I0(x4383), .I1(x4384), .I2(x4385), .I3(n8639), .I4(n8640), .O(n8641));
  LUT3 #(.INIT(8'h96)) lut_n8642 (.I0(n8630), .I1(n8633), .I2(n8634), .O(n8642));
  LUT3 #(.INIT(8'hE8)) lut_n8643 (.I0(n8638), .I1(n8641), .I2(n8642), .O(n8643));
  LUT3 #(.INIT(8'h96)) lut_n8644 (.I0(n8615), .I1(n8623), .I2(n8624), .O(n8644));
  LUT3 #(.INIT(8'hE8)) lut_n8645 (.I0(n8635), .I1(n8643), .I2(n8644), .O(n8645));
  LUT3 #(.INIT(8'hE8)) lut_n8646 (.I0(x4392), .I1(x4393), .I2(x4394), .O(n8646));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8647 (.I0(x4383), .I1(x4384), .I2(x4385), .I3(n8639), .I4(n8640), .O(n8647));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8648 (.I0(x4389), .I1(x4390), .I2(x4391), .I3(n8646), .I4(n8647), .O(n8648));
  LUT3 #(.INIT(8'hE8)) lut_n8649 (.I0(x4398), .I1(x4399), .I2(x4400), .O(n8649));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8650 (.I0(x4389), .I1(x4390), .I2(x4391), .I3(n8646), .I4(n8647), .O(n8650));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8651 (.I0(x4395), .I1(x4396), .I2(x4397), .I3(n8649), .I4(n8650), .O(n8651));
  LUT3 #(.INIT(8'h96)) lut_n8652 (.I0(n8638), .I1(n8641), .I2(n8642), .O(n8652));
  LUT3 #(.INIT(8'hE8)) lut_n8653 (.I0(n8648), .I1(n8651), .I2(n8652), .O(n8653));
  LUT3 #(.INIT(8'hE8)) lut_n8654 (.I0(x4404), .I1(x4405), .I2(x4406), .O(n8654));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8655 (.I0(x4395), .I1(x4396), .I2(x4397), .I3(n8649), .I4(n8650), .O(n8655));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8656 (.I0(x4401), .I1(x4402), .I2(x4403), .I3(n8654), .I4(n8655), .O(n8656));
  LUT3 #(.INIT(8'hE8)) lut_n8657 (.I0(x4410), .I1(x4411), .I2(x4412), .O(n8657));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8658 (.I0(x4401), .I1(x4402), .I2(x4403), .I3(n8654), .I4(n8655), .O(n8658));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8659 (.I0(x4407), .I1(x4408), .I2(x4409), .I3(n8657), .I4(n8658), .O(n8659));
  LUT3 #(.INIT(8'h96)) lut_n8660 (.I0(n8648), .I1(n8651), .I2(n8652), .O(n8660));
  LUT3 #(.INIT(8'hE8)) lut_n8661 (.I0(n8656), .I1(n8659), .I2(n8660), .O(n8661));
  LUT3 #(.INIT(8'h96)) lut_n8662 (.I0(n8635), .I1(n8643), .I2(n8644), .O(n8662));
  LUT3 #(.INIT(8'hE8)) lut_n8663 (.I0(n8653), .I1(n8661), .I2(n8662), .O(n8663));
  LUT3 #(.INIT(8'h96)) lut_n8664 (.I0(n8607), .I1(n8625), .I2(n8626), .O(n8664));
  LUT3 #(.INIT(8'hE8)) lut_n8665 (.I0(n8645), .I1(n8663), .I2(n8664), .O(n8665));
  LUT3 #(.INIT(8'h96)) lut_n8666 (.I0(n8549), .I1(n8587), .I2(n8588), .O(n8666));
  LUT3 #(.INIT(8'hE8)) lut_n8667 (.I0(n8627), .I1(n8665), .I2(n8666), .O(n8667));
  LUT3 #(.INIT(8'h96)) lut_n8668 (.I0(n8429), .I1(n8507), .I2(n8508), .O(n8668));
  LUT3 #(.INIT(8'hE8)) lut_n8669 (.I0(n8589), .I1(n8667), .I2(n8668), .O(n8669));
  LUT3 #(.INIT(8'hE8)) lut_n8670 (.I0(x4416), .I1(x4417), .I2(x4418), .O(n8670));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8671 (.I0(x4407), .I1(x4408), .I2(x4409), .I3(n8657), .I4(n8658), .O(n8671));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8672 (.I0(x4413), .I1(x4414), .I2(x4415), .I3(n8670), .I4(n8671), .O(n8672));
  LUT3 #(.INIT(8'hE8)) lut_n8673 (.I0(x4422), .I1(x4423), .I2(x4424), .O(n8673));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8674 (.I0(x4413), .I1(x4414), .I2(x4415), .I3(n8670), .I4(n8671), .O(n8674));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8675 (.I0(x4419), .I1(x4420), .I2(x4421), .I3(n8673), .I4(n8674), .O(n8675));
  LUT3 #(.INIT(8'h96)) lut_n8676 (.I0(n8656), .I1(n8659), .I2(n8660), .O(n8676));
  LUT3 #(.INIT(8'hE8)) lut_n8677 (.I0(n8672), .I1(n8675), .I2(n8676), .O(n8677));
  LUT3 #(.INIT(8'hE8)) lut_n8678 (.I0(x4428), .I1(x4429), .I2(x4430), .O(n8678));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8679 (.I0(x4419), .I1(x4420), .I2(x4421), .I3(n8673), .I4(n8674), .O(n8679));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8680 (.I0(x4425), .I1(x4426), .I2(x4427), .I3(n8678), .I4(n8679), .O(n8680));
  LUT3 #(.INIT(8'hE8)) lut_n8681 (.I0(x4434), .I1(x4435), .I2(x4436), .O(n8681));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8682 (.I0(x4425), .I1(x4426), .I2(x4427), .I3(n8678), .I4(n8679), .O(n8682));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8683 (.I0(x4431), .I1(x4432), .I2(x4433), .I3(n8681), .I4(n8682), .O(n8683));
  LUT3 #(.INIT(8'h96)) lut_n8684 (.I0(n8672), .I1(n8675), .I2(n8676), .O(n8684));
  LUT3 #(.INIT(8'hE8)) lut_n8685 (.I0(n8680), .I1(n8683), .I2(n8684), .O(n8685));
  LUT3 #(.INIT(8'h96)) lut_n8686 (.I0(n8653), .I1(n8661), .I2(n8662), .O(n8686));
  LUT3 #(.INIT(8'hE8)) lut_n8687 (.I0(n8677), .I1(n8685), .I2(n8686), .O(n8687));
  LUT3 #(.INIT(8'hE8)) lut_n8688 (.I0(x4440), .I1(x4441), .I2(x4442), .O(n8688));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8689 (.I0(x4431), .I1(x4432), .I2(x4433), .I3(n8681), .I4(n8682), .O(n8689));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8690 (.I0(x4437), .I1(x4438), .I2(x4439), .I3(n8688), .I4(n8689), .O(n8690));
  LUT3 #(.INIT(8'hE8)) lut_n8691 (.I0(x4446), .I1(x4447), .I2(x4448), .O(n8691));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8692 (.I0(x4437), .I1(x4438), .I2(x4439), .I3(n8688), .I4(n8689), .O(n8692));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8693 (.I0(x4443), .I1(x4444), .I2(x4445), .I3(n8691), .I4(n8692), .O(n8693));
  LUT3 #(.INIT(8'h96)) lut_n8694 (.I0(n8680), .I1(n8683), .I2(n8684), .O(n8694));
  LUT3 #(.INIT(8'hE8)) lut_n8695 (.I0(n8690), .I1(n8693), .I2(n8694), .O(n8695));
  LUT3 #(.INIT(8'hE8)) lut_n8696 (.I0(x4452), .I1(x4453), .I2(x4454), .O(n8696));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8697 (.I0(x4443), .I1(x4444), .I2(x4445), .I3(n8691), .I4(n8692), .O(n8697));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8698 (.I0(x4449), .I1(x4450), .I2(x4451), .I3(n8696), .I4(n8697), .O(n8698));
  LUT3 #(.INIT(8'hE8)) lut_n8699 (.I0(x4458), .I1(x4459), .I2(x4460), .O(n8699));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8700 (.I0(x4449), .I1(x4450), .I2(x4451), .I3(n8696), .I4(n8697), .O(n8700));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8701 (.I0(x4455), .I1(x4456), .I2(x4457), .I3(n8699), .I4(n8700), .O(n8701));
  LUT3 #(.INIT(8'h96)) lut_n8702 (.I0(n8690), .I1(n8693), .I2(n8694), .O(n8702));
  LUT3 #(.INIT(8'hE8)) lut_n8703 (.I0(n8698), .I1(n8701), .I2(n8702), .O(n8703));
  LUT3 #(.INIT(8'h96)) lut_n8704 (.I0(n8677), .I1(n8685), .I2(n8686), .O(n8704));
  LUT3 #(.INIT(8'hE8)) lut_n8705 (.I0(n8695), .I1(n8703), .I2(n8704), .O(n8705));
  LUT3 #(.INIT(8'h96)) lut_n8706 (.I0(n8645), .I1(n8663), .I2(n8664), .O(n8706));
  LUT3 #(.INIT(8'hE8)) lut_n8707 (.I0(n8687), .I1(n8705), .I2(n8706), .O(n8707));
  LUT3 #(.INIT(8'hE8)) lut_n8708 (.I0(x4464), .I1(x4465), .I2(x4466), .O(n8708));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8709 (.I0(x4455), .I1(x4456), .I2(x4457), .I3(n8699), .I4(n8700), .O(n8709));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8710 (.I0(x4461), .I1(x4462), .I2(x4463), .I3(n8708), .I4(n8709), .O(n8710));
  LUT3 #(.INIT(8'hE8)) lut_n8711 (.I0(x4470), .I1(x4471), .I2(x4472), .O(n8711));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8712 (.I0(x4461), .I1(x4462), .I2(x4463), .I3(n8708), .I4(n8709), .O(n8712));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8713 (.I0(x4467), .I1(x4468), .I2(x4469), .I3(n8711), .I4(n8712), .O(n8713));
  LUT3 #(.INIT(8'h96)) lut_n8714 (.I0(n8698), .I1(n8701), .I2(n8702), .O(n8714));
  LUT3 #(.INIT(8'hE8)) lut_n8715 (.I0(n8710), .I1(n8713), .I2(n8714), .O(n8715));
  LUT3 #(.INIT(8'hE8)) lut_n8716 (.I0(x4476), .I1(x4477), .I2(x4478), .O(n8716));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8717 (.I0(x4467), .I1(x4468), .I2(x4469), .I3(n8711), .I4(n8712), .O(n8717));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8718 (.I0(x4473), .I1(x4474), .I2(x4475), .I3(n8716), .I4(n8717), .O(n8718));
  LUT3 #(.INIT(8'hE8)) lut_n8719 (.I0(x4482), .I1(x4483), .I2(x4484), .O(n8719));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8720 (.I0(x4473), .I1(x4474), .I2(x4475), .I3(n8716), .I4(n8717), .O(n8720));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8721 (.I0(x4479), .I1(x4480), .I2(x4481), .I3(n8719), .I4(n8720), .O(n8721));
  LUT3 #(.INIT(8'h96)) lut_n8722 (.I0(n8710), .I1(n8713), .I2(n8714), .O(n8722));
  LUT3 #(.INIT(8'hE8)) lut_n8723 (.I0(n8718), .I1(n8721), .I2(n8722), .O(n8723));
  LUT3 #(.INIT(8'h96)) lut_n8724 (.I0(n8695), .I1(n8703), .I2(n8704), .O(n8724));
  LUT3 #(.INIT(8'hE8)) lut_n8725 (.I0(n8715), .I1(n8723), .I2(n8724), .O(n8725));
  LUT3 #(.INIT(8'hE8)) lut_n8726 (.I0(x4488), .I1(x4489), .I2(x4490), .O(n8726));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8727 (.I0(x4479), .I1(x4480), .I2(x4481), .I3(n8719), .I4(n8720), .O(n8727));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8728 (.I0(x4485), .I1(x4486), .I2(x4487), .I3(n8726), .I4(n8727), .O(n8728));
  LUT3 #(.INIT(8'hE8)) lut_n8729 (.I0(x4494), .I1(x4495), .I2(x4496), .O(n8729));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8730 (.I0(x4485), .I1(x4486), .I2(x4487), .I3(n8726), .I4(n8727), .O(n8730));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8731 (.I0(x4491), .I1(x4492), .I2(x4493), .I3(n8729), .I4(n8730), .O(n8731));
  LUT3 #(.INIT(8'h96)) lut_n8732 (.I0(n8718), .I1(n8721), .I2(n8722), .O(n8732));
  LUT3 #(.INIT(8'hE8)) lut_n8733 (.I0(n8728), .I1(n8731), .I2(n8732), .O(n8733));
  LUT3 #(.INIT(8'hE8)) lut_n8734 (.I0(x4500), .I1(x4501), .I2(x4502), .O(n8734));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8735 (.I0(x4491), .I1(x4492), .I2(x4493), .I3(n8729), .I4(n8730), .O(n8735));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8736 (.I0(x4497), .I1(x4498), .I2(x4499), .I3(n8734), .I4(n8735), .O(n8736));
  LUT3 #(.INIT(8'hE8)) lut_n8737 (.I0(x4506), .I1(x4507), .I2(x4508), .O(n8737));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8738 (.I0(x4497), .I1(x4498), .I2(x4499), .I3(n8734), .I4(n8735), .O(n8738));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8739 (.I0(x4503), .I1(x4504), .I2(x4505), .I3(n8737), .I4(n8738), .O(n8739));
  LUT3 #(.INIT(8'h96)) lut_n8740 (.I0(n8728), .I1(n8731), .I2(n8732), .O(n8740));
  LUT3 #(.INIT(8'hE8)) lut_n8741 (.I0(n8736), .I1(n8739), .I2(n8740), .O(n8741));
  LUT3 #(.INIT(8'h96)) lut_n8742 (.I0(n8715), .I1(n8723), .I2(n8724), .O(n8742));
  LUT3 #(.INIT(8'hE8)) lut_n8743 (.I0(n8733), .I1(n8741), .I2(n8742), .O(n8743));
  LUT3 #(.INIT(8'h96)) lut_n8744 (.I0(n8687), .I1(n8705), .I2(n8706), .O(n8744));
  LUT3 #(.INIT(8'hE8)) lut_n8745 (.I0(n8725), .I1(n8743), .I2(n8744), .O(n8745));
  LUT3 #(.INIT(8'h96)) lut_n8746 (.I0(n8627), .I1(n8665), .I2(n8666), .O(n8746));
  LUT3 #(.INIT(8'hE8)) lut_n8747 (.I0(n8707), .I1(n8745), .I2(n8746), .O(n8747));
  LUT3 #(.INIT(8'hE8)) lut_n8748 (.I0(x4512), .I1(x4513), .I2(x4514), .O(n8748));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8749 (.I0(x4503), .I1(x4504), .I2(x4505), .I3(n8737), .I4(n8738), .O(n8749));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8750 (.I0(x4509), .I1(x4510), .I2(x4511), .I3(n8748), .I4(n8749), .O(n8750));
  LUT3 #(.INIT(8'hE8)) lut_n8751 (.I0(x4518), .I1(x4519), .I2(x4520), .O(n8751));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8752 (.I0(x4509), .I1(x4510), .I2(x4511), .I3(n8748), .I4(n8749), .O(n8752));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8753 (.I0(x4515), .I1(x4516), .I2(x4517), .I3(n8751), .I4(n8752), .O(n8753));
  LUT3 #(.INIT(8'h96)) lut_n8754 (.I0(n8736), .I1(n8739), .I2(n8740), .O(n8754));
  LUT3 #(.INIT(8'hE8)) lut_n8755 (.I0(n8750), .I1(n8753), .I2(n8754), .O(n8755));
  LUT3 #(.INIT(8'hE8)) lut_n8756 (.I0(x4524), .I1(x4525), .I2(x4526), .O(n8756));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8757 (.I0(x4515), .I1(x4516), .I2(x4517), .I3(n8751), .I4(n8752), .O(n8757));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8758 (.I0(x4521), .I1(x4522), .I2(x4523), .I3(n8756), .I4(n8757), .O(n8758));
  LUT3 #(.INIT(8'hE8)) lut_n8759 (.I0(x4530), .I1(x4531), .I2(x4532), .O(n8759));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8760 (.I0(x4521), .I1(x4522), .I2(x4523), .I3(n8756), .I4(n8757), .O(n8760));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8761 (.I0(x4527), .I1(x4528), .I2(x4529), .I3(n8759), .I4(n8760), .O(n8761));
  LUT3 #(.INIT(8'h96)) lut_n8762 (.I0(n8750), .I1(n8753), .I2(n8754), .O(n8762));
  LUT3 #(.INIT(8'hE8)) lut_n8763 (.I0(n8758), .I1(n8761), .I2(n8762), .O(n8763));
  LUT3 #(.INIT(8'h96)) lut_n8764 (.I0(n8733), .I1(n8741), .I2(n8742), .O(n8764));
  LUT3 #(.INIT(8'hE8)) lut_n8765 (.I0(n8755), .I1(n8763), .I2(n8764), .O(n8765));
  LUT3 #(.INIT(8'hE8)) lut_n8766 (.I0(x4536), .I1(x4537), .I2(x4538), .O(n8766));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8767 (.I0(x4527), .I1(x4528), .I2(x4529), .I3(n8759), .I4(n8760), .O(n8767));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8768 (.I0(x4533), .I1(x4534), .I2(x4535), .I3(n8766), .I4(n8767), .O(n8768));
  LUT3 #(.INIT(8'hE8)) lut_n8769 (.I0(x4542), .I1(x4543), .I2(x4544), .O(n8769));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8770 (.I0(x4533), .I1(x4534), .I2(x4535), .I3(n8766), .I4(n8767), .O(n8770));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8771 (.I0(x4539), .I1(x4540), .I2(x4541), .I3(n8769), .I4(n8770), .O(n8771));
  LUT3 #(.INIT(8'h96)) lut_n8772 (.I0(n8758), .I1(n8761), .I2(n8762), .O(n8772));
  LUT3 #(.INIT(8'hE8)) lut_n8773 (.I0(n8768), .I1(n8771), .I2(n8772), .O(n8773));
  LUT3 #(.INIT(8'hE8)) lut_n8774 (.I0(x4548), .I1(x4549), .I2(x4550), .O(n8774));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8775 (.I0(x4539), .I1(x4540), .I2(x4541), .I3(n8769), .I4(n8770), .O(n8775));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8776 (.I0(x4545), .I1(x4546), .I2(x4547), .I3(n8774), .I4(n8775), .O(n8776));
  LUT3 #(.INIT(8'hE8)) lut_n8777 (.I0(x4554), .I1(x4555), .I2(x4556), .O(n8777));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8778 (.I0(x4545), .I1(x4546), .I2(x4547), .I3(n8774), .I4(n8775), .O(n8778));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8779 (.I0(x4551), .I1(x4552), .I2(x4553), .I3(n8777), .I4(n8778), .O(n8779));
  LUT3 #(.INIT(8'h96)) lut_n8780 (.I0(n8768), .I1(n8771), .I2(n8772), .O(n8780));
  LUT3 #(.INIT(8'hE8)) lut_n8781 (.I0(n8776), .I1(n8779), .I2(n8780), .O(n8781));
  LUT3 #(.INIT(8'h96)) lut_n8782 (.I0(n8755), .I1(n8763), .I2(n8764), .O(n8782));
  LUT3 #(.INIT(8'hE8)) lut_n8783 (.I0(n8773), .I1(n8781), .I2(n8782), .O(n8783));
  LUT3 #(.INIT(8'h96)) lut_n8784 (.I0(n8725), .I1(n8743), .I2(n8744), .O(n8784));
  LUT3 #(.INIT(8'hE8)) lut_n8785 (.I0(n8765), .I1(n8783), .I2(n8784), .O(n8785));
  LUT3 #(.INIT(8'hE8)) lut_n8786 (.I0(x4560), .I1(x4561), .I2(x4562), .O(n8786));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8787 (.I0(x4551), .I1(x4552), .I2(x4553), .I3(n8777), .I4(n8778), .O(n8787));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8788 (.I0(x4557), .I1(x4558), .I2(x4559), .I3(n8786), .I4(n8787), .O(n8788));
  LUT3 #(.INIT(8'hE8)) lut_n8789 (.I0(x4566), .I1(x4567), .I2(x4568), .O(n8789));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8790 (.I0(x4557), .I1(x4558), .I2(x4559), .I3(n8786), .I4(n8787), .O(n8790));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8791 (.I0(x4563), .I1(x4564), .I2(x4565), .I3(n8789), .I4(n8790), .O(n8791));
  LUT3 #(.INIT(8'h96)) lut_n8792 (.I0(n8776), .I1(n8779), .I2(n8780), .O(n8792));
  LUT3 #(.INIT(8'hE8)) lut_n8793 (.I0(n8788), .I1(n8791), .I2(n8792), .O(n8793));
  LUT3 #(.INIT(8'hE8)) lut_n8794 (.I0(x4572), .I1(x4573), .I2(x4574), .O(n8794));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8795 (.I0(x4563), .I1(x4564), .I2(x4565), .I3(n8789), .I4(n8790), .O(n8795));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8796 (.I0(x4569), .I1(x4570), .I2(x4571), .I3(n8794), .I4(n8795), .O(n8796));
  LUT3 #(.INIT(8'hE8)) lut_n8797 (.I0(x4578), .I1(x4579), .I2(x4580), .O(n8797));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8798 (.I0(x4569), .I1(x4570), .I2(x4571), .I3(n8794), .I4(n8795), .O(n8798));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8799 (.I0(x4575), .I1(x4576), .I2(x4577), .I3(n8797), .I4(n8798), .O(n8799));
  LUT3 #(.INIT(8'h96)) lut_n8800 (.I0(n8788), .I1(n8791), .I2(n8792), .O(n8800));
  LUT3 #(.INIT(8'hE8)) lut_n8801 (.I0(n8796), .I1(n8799), .I2(n8800), .O(n8801));
  LUT3 #(.INIT(8'h96)) lut_n8802 (.I0(n8773), .I1(n8781), .I2(n8782), .O(n8802));
  LUT3 #(.INIT(8'hE8)) lut_n8803 (.I0(n8793), .I1(n8801), .I2(n8802), .O(n8803));
  LUT3 #(.INIT(8'hE8)) lut_n8804 (.I0(x4584), .I1(x4585), .I2(x4586), .O(n8804));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8805 (.I0(x4575), .I1(x4576), .I2(x4577), .I3(n8797), .I4(n8798), .O(n8805));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8806 (.I0(x4581), .I1(x4582), .I2(x4583), .I3(n8804), .I4(n8805), .O(n8806));
  LUT3 #(.INIT(8'hE8)) lut_n8807 (.I0(x4590), .I1(x4591), .I2(x4592), .O(n8807));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8808 (.I0(x4581), .I1(x4582), .I2(x4583), .I3(n8804), .I4(n8805), .O(n8808));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8809 (.I0(x4587), .I1(x4588), .I2(x4589), .I3(n8807), .I4(n8808), .O(n8809));
  LUT3 #(.INIT(8'h96)) lut_n8810 (.I0(n8796), .I1(n8799), .I2(n8800), .O(n8810));
  LUT3 #(.INIT(8'hE8)) lut_n8811 (.I0(n8806), .I1(n8809), .I2(n8810), .O(n8811));
  LUT3 #(.INIT(8'hE8)) lut_n8812 (.I0(x4596), .I1(x4597), .I2(x4598), .O(n8812));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8813 (.I0(x4587), .I1(x4588), .I2(x4589), .I3(n8807), .I4(n8808), .O(n8813));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8814 (.I0(x4593), .I1(x4594), .I2(x4595), .I3(n8812), .I4(n8813), .O(n8814));
  LUT3 #(.INIT(8'hE8)) lut_n8815 (.I0(x4602), .I1(x4603), .I2(x4604), .O(n8815));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8816 (.I0(x4593), .I1(x4594), .I2(x4595), .I3(n8812), .I4(n8813), .O(n8816));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8817 (.I0(x4599), .I1(x4600), .I2(x4601), .I3(n8815), .I4(n8816), .O(n8817));
  LUT3 #(.INIT(8'h96)) lut_n8818 (.I0(n8806), .I1(n8809), .I2(n8810), .O(n8818));
  LUT3 #(.INIT(8'hE8)) lut_n8819 (.I0(n8814), .I1(n8817), .I2(n8818), .O(n8819));
  LUT3 #(.INIT(8'h96)) lut_n8820 (.I0(n8793), .I1(n8801), .I2(n8802), .O(n8820));
  LUT3 #(.INIT(8'hE8)) lut_n8821 (.I0(n8811), .I1(n8819), .I2(n8820), .O(n8821));
  LUT3 #(.INIT(8'h96)) lut_n8822 (.I0(n8765), .I1(n8783), .I2(n8784), .O(n8822));
  LUT3 #(.INIT(8'hE8)) lut_n8823 (.I0(n8803), .I1(n8821), .I2(n8822), .O(n8823));
  LUT3 #(.INIT(8'h96)) lut_n8824 (.I0(n8707), .I1(n8745), .I2(n8746), .O(n8824));
  LUT3 #(.INIT(8'hE8)) lut_n8825 (.I0(n8785), .I1(n8823), .I2(n8824), .O(n8825));
  LUT3 #(.INIT(8'h96)) lut_n8826 (.I0(n8589), .I1(n8667), .I2(n8668), .O(n8826));
  LUT3 #(.INIT(8'hE8)) lut_n8827 (.I0(n8747), .I1(n8825), .I2(n8826), .O(n8827));
  LUT3 #(.INIT(8'h96)) lut_n8828 (.I0(n8351), .I1(n8509), .I2(n8510), .O(n8828));
  LUT3 #(.INIT(8'hE8)) lut_n8829 (.I0(n8669), .I1(n8827), .I2(n8828), .O(n8829));
  LUT3 #(.INIT(8'h96)) lut_n8830 (.I0(n7873), .I1(n8191), .I2(n8192), .O(n8830));
  LUT3 #(.INIT(8'hE8)) lut_n8831 (.I0(n8511), .I1(n8829), .I2(n8830), .O(n8831));
  LUT3 #(.INIT(8'h96)) lut_n8832 (.I0(n6278), .I1(n6916), .I2(n7554), .O(n8832));
  LUT3 #(.INIT(8'hE8)) lut_n8833 (.I0(n8193), .I1(n8831), .I2(n8832), .O(n8833));
  LUT3 #(.INIT(8'hE8)) lut_n8834 (.I0(x4608), .I1(x4609), .I2(x4610), .O(n8834));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8835 (.I0(x4599), .I1(x4600), .I2(x4601), .I3(n8815), .I4(n8816), .O(n8835));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8836 (.I0(x4605), .I1(x4606), .I2(x4607), .I3(n8834), .I4(n8835), .O(n8836));
  LUT3 #(.INIT(8'hE8)) lut_n8837 (.I0(x4614), .I1(x4615), .I2(x4616), .O(n8837));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8838 (.I0(x4605), .I1(x4606), .I2(x4607), .I3(n8834), .I4(n8835), .O(n8838));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8839 (.I0(x4611), .I1(x4612), .I2(x4613), .I3(n8837), .I4(n8838), .O(n8839));
  LUT3 #(.INIT(8'h96)) lut_n8840 (.I0(n8814), .I1(n8817), .I2(n8818), .O(n8840));
  LUT3 #(.INIT(8'hE8)) lut_n8841 (.I0(n8836), .I1(n8839), .I2(n8840), .O(n8841));
  LUT3 #(.INIT(8'hE8)) lut_n8842 (.I0(x4620), .I1(x4621), .I2(x4622), .O(n8842));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8843 (.I0(x4611), .I1(x4612), .I2(x4613), .I3(n8837), .I4(n8838), .O(n8843));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8844 (.I0(x4617), .I1(x4618), .I2(x4619), .I3(n8842), .I4(n8843), .O(n8844));
  LUT3 #(.INIT(8'hE8)) lut_n8845 (.I0(x4626), .I1(x4627), .I2(x4628), .O(n8845));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8846 (.I0(x4617), .I1(x4618), .I2(x4619), .I3(n8842), .I4(n8843), .O(n8846));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8847 (.I0(x4623), .I1(x4624), .I2(x4625), .I3(n8845), .I4(n8846), .O(n8847));
  LUT3 #(.INIT(8'h96)) lut_n8848 (.I0(n8836), .I1(n8839), .I2(n8840), .O(n8848));
  LUT3 #(.INIT(8'hE8)) lut_n8849 (.I0(n8844), .I1(n8847), .I2(n8848), .O(n8849));
  LUT3 #(.INIT(8'h96)) lut_n8850 (.I0(n8811), .I1(n8819), .I2(n8820), .O(n8850));
  LUT3 #(.INIT(8'hE8)) lut_n8851 (.I0(n8841), .I1(n8849), .I2(n8850), .O(n8851));
  LUT3 #(.INIT(8'hE8)) lut_n8852 (.I0(x4632), .I1(x4633), .I2(x4634), .O(n8852));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8853 (.I0(x4623), .I1(x4624), .I2(x4625), .I3(n8845), .I4(n8846), .O(n8853));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8854 (.I0(x4629), .I1(x4630), .I2(x4631), .I3(n8852), .I4(n8853), .O(n8854));
  LUT3 #(.INIT(8'hE8)) lut_n8855 (.I0(x4638), .I1(x4639), .I2(x4640), .O(n8855));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8856 (.I0(x4629), .I1(x4630), .I2(x4631), .I3(n8852), .I4(n8853), .O(n8856));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8857 (.I0(x4635), .I1(x4636), .I2(x4637), .I3(n8855), .I4(n8856), .O(n8857));
  LUT3 #(.INIT(8'h96)) lut_n8858 (.I0(n8844), .I1(n8847), .I2(n8848), .O(n8858));
  LUT3 #(.INIT(8'hE8)) lut_n8859 (.I0(n8854), .I1(n8857), .I2(n8858), .O(n8859));
  LUT3 #(.INIT(8'hE8)) lut_n8860 (.I0(x4644), .I1(x4645), .I2(x4646), .O(n8860));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8861 (.I0(x4635), .I1(x4636), .I2(x4637), .I3(n8855), .I4(n8856), .O(n8861));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8862 (.I0(x4641), .I1(x4642), .I2(x4643), .I3(n8860), .I4(n8861), .O(n8862));
  LUT3 #(.INIT(8'hE8)) lut_n8863 (.I0(x4650), .I1(x4651), .I2(x4652), .O(n8863));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8864 (.I0(x4641), .I1(x4642), .I2(x4643), .I3(n8860), .I4(n8861), .O(n8864));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8865 (.I0(x4647), .I1(x4648), .I2(x4649), .I3(n8863), .I4(n8864), .O(n8865));
  LUT3 #(.INIT(8'h96)) lut_n8866 (.I0(n8854), .I1(n8857), .I2(n8858), .O(n8866));
  LUT3 #(.INIT(8'hE8)) lut_n8867 (.I0(n8862), .I1(n8865), .I2(n8866), .O(n8867));
  LUT3 #(.INIT(8'h96)) lut_n8868 (.I0(n8841), .I1(n8849), .I2(n8850), .O(n8868));
  LUT3 #(.INIT(8'hE8)) lut_n8869 (.I0(n8859), .I1(n8867), .I2(n8868), .O(n8869));
  LUT3 #(.INIT(8'h96)) lut_n8870 (.I0(n8803), .I1(n8821), .I2(n8822), .O(n8870));
  LUT3 #(.INIT(8'hE8)) lut_n8871 (.I0(n8851), .I1(n8869), .I2(n8870), .O(n8871));
  LUT3 #(.INIT(8'hE8)) lut_n8872 (.I0(x4656), .I1(x4657), .I2(x4658), .O(n8872));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8873 (.I0(x4647), .I1(x4648), .I2(x4649), .I3(n8863), .I4(n8864), .O(n8873));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8874 (.I0(x4653), .I1(x4654), .I2(x4655), .I3(n8872), .I4(n8873), .O(n8874));
  LUT3 #(.INIT(8'hE8)) lut_n8875 (.I0(x4662), .I1(x4663), .I2(x4664), .O(n8875));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8876 (.I0(x4653), .I1(x4654), .I2(x4655), .I3(n8872), .I4(n8873), .O(n8876));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8877 (.I0(x4659), .I1(x4660), .I2(x4661), .I3(n8875), .I4(n8876), .O(n8877));
  LUT3 #(.INIT(8'h96)) lut_n8878 (.I0(n8862), .I1(n8865), .I2(n8866), .O(n8878));
  LUT3 #(.INIT(8'hE8)) lut_n8879 (.I0(n8874), .I1(n8877), .I2(n8878), .O(n8879));
  LUT3 #(.INIT(8'hE8)) lut_n8880 (.I0(x4668), .I1(x4669), .I2(x4670), .O(n8880));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8881 (.I0(x4659), .I1(x4660), .I2(x4661), .I3(n8875), .I4(n8876), .O(n8881));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8882 (.I0(x4665), .I1(x4666), .I2(x4667), .I3(n8880), .I4(n8881), .O(n8882));
  LUT3 #(.INIT(8'hE8)) lut_n8883 (.I0(x4674), .I1(x4675), .I2(x4676), .O(n8883));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8884 (.I0(x4665), .I1(x4666), .I2(x4667), .I3(n8880), .I4(n8881), .O(n8884));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8885 (.I0(x4671), .I1(x4672), .I2(x4673), .I3(n8883), .I4(n8884), .O(n8885));
  LUT3 #(.INIT(8'h96)) lut_n8886 (.I0(n8874), .I1(n8877), .I2(n8878), .O(n8886));
  LUT3 #(.INIT(8'hE8)) lut_n8887 (.I0(n8882), .I1(n8885), .I2(n8886), .O(n8887));
  LUT3 #(.INIT(8'h96)) lut_n8888 (.I0(n8859), .I1(n8867), .I2(n8868), .O(n8888));
  LUT3 #(.INIT(8'hE8)) lut_n8889 (.I0(n8879), .I1(n8887), .I2(n8888), .O(n8889));
  LUT3 #(.INIT(8'hE8)) lut_n8890 (.I0(x4680), .I1(x4681), .I2(x4682), .O(n8890));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8891 (.I0(x4671), .I1(x4672), .I2(x4673), .I3(n8883), .I4(n8884), .O(n8891));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8892 (.I0(x4677), .I1(x4678), .I2(x4679), .I3(n8890), .I4(n8891), .O(n8892));
  LUT3 #(.INIT(8'hE8)) lut_n8893 (.I0(x4686), .I1(x4687), .I2(x4688), .O(n8893));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8894 (.I0(x4677), .I1(x4678), .I2(x4679), .I3(n8890), .I4(n8891), .O(n8894));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8895 (.I0(x4683), .I1(x4684), .I2(x4685), .I3(n8893), .I4(n8894), .O(n8895));
  LUT3 #(.INIT(8'h96)) lut_n8896 (.I0(n8882), .I1(n8885), .I2(n8886), .O(n8896));
  LUT3 #(.INIT(8'hE8)) lut_n8897 (.I0(n8892), .I1(n8895), .I2(n8896), .O(n8897));
  LUT3 #(.INIT(8'hE8)) lut_n8898 (.I0(x4692), .I1(x4693), .I2(x4694), .O(n8898));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8899 (.I0(x4683), .I1(x4684), .I2(x4685), .I3(n8893), .I4(n8894), .O(n8899));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8900 (.I0(x4689), .I1(x4690), .I2(x4691), .I3(n8898), .I4(n8899), .O(n8900));
  LUT3 #(.INIT(8'hE8)) lut_n8901 (.I0(x4698), .I1(x4699), .I2(x4700), .O(n8901));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8902 (.I0(x4689), .I1(x4690), .I2(x4691), .I3(n8898), .I4(n8899), .O(n8902));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8903 (.I0(x4695), .I1(x4696), .I2(x4697), .I3(n8901), .I4(n8902), .O(n8903));
  LUT3 #(.INIT(8'h96)) lut_n8904 (.I0(n8892), .I1(n8895), .I2(n8896), .O(n8904));
  LUT3 #(.INIT(8'hE8)) lut_n8905 (.I0(n8900), .I1(n8903), .I2(n8904), .O(n8905));
  LUT3 #(.INIT(8'h96)) lut_n8906 (.I0(n8879), .I1(n8887), .I2(n8888), .O(n8906));
  LUT3 #(.INIT(8'hE8)) lut_n8907 (.I0(n8897), .I1(n8905), .I2(n8906), .O(n8907));
  LUT3 #(.INIT(8'h96)) lut_n8908 (.I0(n8851), .I1(n8869), .I2(n8870), .O(n8908));
  LUT3 #(.INIT(8'hE8)) lut_n8909 (.I0(n8889), .I1(n8907), .I2(n8908), .O(n8909));
  LUT3 #(.INIT(8'h96)) lut_n8910 (.I0(n8785), .I1(n8823), .I2(n8824), .O(n8910));
  LUT3 #(.INIT(8'hE8)) lut_n8911 (.I0(n8871), .I1(n8909), .I2(n8910), .O(n8911));
  LUT3 #(.INIT(8'hE8)) lut_n8912 (.I0(x4704), .I1(x4705), .I2(x4706), .O(n8912));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8913 (.I0(x4695), .I1(x4696), .I2(x4697), .I3(n8901), .I4(n8902), .O(n8913));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8914 (.I0(x4701), .I1(x4702), .I2(x4703), .I3(n8912), .I4(n8913), .O(n8914));
  LUT3 #(.INIT(8'hE8)) lut_n8915 (.I0(x4710), .I1(x4711), .I2(x4712), .O(n8915));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8916 (.I0(x4701), .I1(x4702), .I2(x4703), .I3(n8912), .I4(n8913), .O(n8916));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8917 (.I0(x4707), .I1(x4708), .I2(x4709), .I3(n8915), .I4(n8916), .O(n8917));
  LUT3 #(.INIT(8'h96)) lut_n8918 (.I0(n8900), .I1(n8903), .I2(n8904), .O(n8918));
  LUT3 #(.INIT(8'hE8)) lut_n8919 (.I0(n8914), .I1(n8917), .I2(n8918), .O(n8919));
  LUT3 #(.INIT(8'hE8)) lut_n8920 (.I0(x4716), .I1(x4717), .I2(x4718), .O(n8920));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8921 (.I0(x4707), .I1(x4708), .I2(x4709), .I3(n8915), .I4(n8916), .O(n8921));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8922 (.I0(x4713), .I1(x4714), .I2(x4715), .I3(n8920), .I4(n8921), .O(n8922));
  LUT3 #(.INIT(8'hE8)) lut_n8923 (.I0(x4722), .I1(x4723), .I2(x4724), .O(n8923));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8924 (.I0(x4713), .I1(x4714), .I2(x4715), .I3(n8920), .I4(n8921), .O(n8924));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8925 (.I0(x4719), .I1(x4720), .I2(x4721), .I3(n8923), .I4(n8924), .O(n8925));
  LUT3 #(.INIT(8'h96)) lut_n8926 (.I0(n8914), .I1(n8917), .I2(n8918), .O(n8926));
  LUT3 #(.INIT(8'hE8)) lut_n8927 (.I0(n8922), .I1(n8925), .I2(n8926), .O(n8927));
  LUT3 #(.INIT(8'h96)) lut_n8928 (.I0(n8897), .I1(n8905), .I2(n8906), .O(n8928));
  LUT3 #(.INIT(8'hE8)) lut_n8929 (.I0(n8919), .I1(n8927), .I2(n8928), .O(n8929));
  LUT3 #(.INIT(8'hE8)) lut_n8930 (.I0(x4728), .I1(x4729), .I2(x4730), .O(n8930));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8931 (.I0(x4719), .I1(x4720), .I2(x4721), .I3(n8923), .I4(n8924), .O(n8931));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8932 (.I0(x4725), .I1(x4726), .I2(x4727), .I3(n8930), .I4(n8931), .O(n8932));
  LUT3 #(.INIT(8'hE8)) lut_n8933 (.I0(x4734), .I1(x4735), .I2(x4736), .O(n8933));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8934 (.I0(x4725), .I1(x4726), .I2(x4727), .I3(n8930), .I4(n8931), .O(n8934));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8935 (.I0(x4731), .I1(x4732), .I2(x4733), .I3(n8933), .I4(n8934), .O(n8935));
  LUT3 #(.INIT(8'h96)) lut_n8936 (.I0(n8922), .I1(n8925), .I2(n8926), .O(n8936));
  LUT3 #(.INIT(8'hE8)) lut_n8937 (.I0(n8932), .I1(n8935), .I2(n8936), .O(n8937));
  LUT3 #(.INIT(8'hE8)) lut_n8938 (.I0(x4740), .I1(x4741), .I2(x4742), .O(n8938));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8939 (.I0(x4731), .I1(x4732), .I2(x4733), .I3(n8933), .I4(n8934), .O(n8939));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8940 (.I0(x4737), .I1(x4738), .I2(x4739), .I3(n8938), .I4(n8939), .O(n8940));
  LUT3 #(.INIT(8'hE8)) lut_n8941 (.I0(x4746), .I1(x4747), .I2(x4748), .O(n8941));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8942 (.I0(x4737), .I1(x4738), .I2(x4739), .I3(n8938), .I4(n8939), .O(n8942));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8943 (.I0(x4743), .I1(x4744), .I2(x4745), .I3(n8941), .I4(n8942), .O(n8943));
  LUT3 #(.INIT(8'h96)) lut_n8944 (.I0(n8932), .I1(n8935), .I2(n8936), .O(n8944));
  LUT3 #(.INIT(8'hE8)) lut_n8945 (.I0(n8940), .I1(n8943), .I2(n8944), .O(n8945));
  LUT3 #(.INIT(8'h96)) lut_n8946 (.I0(n8919), .I1(n8927), .I2(n8928), .O(n8946));
  LUT3 #(.INIT(8'hE8)) lut_n8947 (.I0(n8937), .I1(n8945), .I2(n8946), .O(n8947));
  LUT3 #(.INIT(8'h96)) lut_n8948 (.I0(n8889), .I1(n8907), .I2(n8908), .O(n8948));
  LUT3 #(.INIT(8'hE8)) lut_n8949 (.I0(n8929), .I1(n8947), .I2(n8948), .O(n8949));
  LUT3 #(.INIT(8'hE8)) lut_n8950 (.I0(x4752), .I1(x4753), .I2(x4754), .O(n8950));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8951 (.I0(x4743), .I1(x4744), .I2(x4745), .I3(n8941), .I4(n8942), .O(n8951));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8952 (.I0(x4749), .I1(x4750), .I2(x4751), .I3(n8950), .I4(n8951), .O(n8952));
  LUT3 #(.INIT(8'hE8)) lut_n8953 (.I0(x4758), .I1(x4759), .I2(x4760), .O(n8953));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8954 (.I0(x4749), .I1(x4750), .I2(x4751), .I3(n8950), .I4(n8951), .O(n8954));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8955 (.I0(x4755), .I1(x4756), .I2(x4757), .I3(n8953), .I4(n8954), .O(n8955));
  LUT3 #(.INIT(8'h96)) lut_n8956 (.I0(n8940), .I1(n8943), .I2(n8944), .O(n8956));
  LUT3 #(.INIT(8'hE8)) lut_n8957 (.I0(n8952), .I1(n8955), .I2(n8956), .O(n8957));
  LUT3 #(.INIT(8'hE8)) lut_n8958 (.I0(x4764), .I1(x4765), .I2(x4766), .O(n8958));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8959 (.I0(x4755), .I1(x4756), .I2(x4757), .I3(n8953), .I4(n8954), .O(n8959));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8960 (.I0(x4761), .I1(x4762), .I2(x4763), .I3(n8958), .I4(n8959), .O(n8960));
  LUT3 #(.INIT(8'hE8)) lut_n8961 (.I0(x4770), .I1(x4771), .I2(x4772), .O(n8961));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8962 (.I0(x4761), .I1(x4762), .I2(x4763), .I3(n8958), .I4(n8959), .O(n8962));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8963 (.I0(x4767), .I1(x4768), .I2(x4769), .I3(n8961), .I4(n8962), .O(n8963));
  LUT3 #(.INIT(8'h96)) lut_n8964 (.I0(n8952), .I1(n8955), .I2(n8956), .O(n8964));
  LUT3 #(.INIT(8'hE8)) lut_n8965 (.I0(n8960), .I1(n8963), .I2(n8964), .O(n8965));
  LUT3 #(.INIT(8'h96)) lut_n8966 (.I0(n8937), .I1(n8945), .I2(n8946), .O(n8966));
  LUT3 #(.INIT(8'hE8)) lut_n8967 (.I0(n8957), .I1(n8965), .I2(n8966), .O(n8967));
  LUT3 #(.INIT(8'hE8)) lut_n8968 (.I0(x4776), .I1(x4777), .I2(x4778), .O(n8968));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8969 (.I0(x4767), .I1(x4768), .I2(x4769), .I3(n8961), .I4(n8962), .O(n8969));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8970 (.I0(x4773), .I1(x4774), .I2(x4775), .I3(n8968), .I4(n8969), .O(n8970));
  LUT3 #(.INIT(8'hE8)) lut_n8971 (.I0(x4782), .I1(x4783), .I2(x4784), .O(n8971));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8972 (.I0(x4773), .I1(x4774), .I2(x4775), .I3(n8968), .I4(n8969), .O(n8972));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8973 (.I0(x4779), .I1(x4780), .I2(x4781), .I3(n8971), .I4(n8972), .O(n8973));
  LUT3 #(.INIT(8'h96)) lut_n8974 (.I0(n8960), .I1(n8963), .I2(n8964), .O(n8974));
  LUT3 #(.INIT(8'hE8)) lut_n8975 (.I0(n8970), .I1(n8973), .I2(n8974), .O(n8975));
  LUT3 #(.INIT(8'hE8)) lut_n8976 (.I0(x4788), .I1(x4789), .I2(x4790), .O(n8976));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8977 (.I0(x4779), .I1(x4780), .I2(x4781), .I3(n8971), .I4(n8972), .O(n8977));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8978 (.I0(x4785), .I1(x4786), .I2(x4787), .I3(n8976), .I4(n8977), .O(n8978));
  LUT3 #(.INIT(8'hE8)) lut_n8979 (.I0(x4794), .I1(x4795), .I2(x4796), .O(n8979));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8980 (.I0(x4785), .I1(x4786), .I2(x4787), .I3(n8976), .I4(n8977), .O(n8980));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8981 (.I0(x4791), .I1(x4792), .I2(x4793), .I3(n8979), .I4(n8980), .O(n8981));
  LUT3 #(.INIT(8'h96)) lut_n8982 (.I0(n8970), .I1(n8973), .I2(n8974), .O(n8982));
  LUT3 #(.INIT(8'hE8)) lut_n8983 (.I0(n8978), .I1(n8981), .I2(n8982), .O(n8983));
  LUT3 #(.INIT(8'h96)) lut_n8984 (.I0(n8957), .I1(n8965), .I2(n8966), .O(n8984));
  LUT3 #(.INIT(8'hE8)) lut_n8985 (.I0(n8975), .I1(n8983), .I2(n8984), .O(n8985));
  LUT3 #(.INIT(8'h96)) lut_n8986 (.I0(n8929), .I1(n8947), .I2(n8948), .O(n8986));
  LUT3 #(.INIT(8'hE8)) lut_n8987 (.I0(n8967), .I1(n8985), .I2(n8986), .O(n8987));
  LUT3 #(.INIT(8'h96)) lut_n8988 (.I0(n8871), .I1(n8909), .I2(n8910), .O(n8988));
  LUT3 #(.INIT(8'hE8)) lut_n8989 (.I0(n8949), .I1(n8987), .I2(n8988), .O(n8989));
  LUT3 #(.INIT(8'h96)) lut_n8990 (.I0(n8747), .I1(n8825), .I2(n8826), .O(n8990));
  LUT3 #(.INIT(8'hE8)) lut_n8991 (.I0(n8911), .I1(n8989), .I2(n8990), .O(n8991));
  LUT3 #(.INIT(8'hE8)) lut_n8992 (.I0(x4800), .I1(x4801), .I2(x4802), .O(n8992));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8993 (.I0(x4791), .I1(x4792), .I2(x4793), .I3(n8979), .I4(n8980), .O(n8993));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8994 (.I0(x4797), .I1(x4798), .I2(x4799), .I3(n8992), .I4(n8993), .O(n8994));
  LUT3 #(.INIT(8'hE8)) lut_n8995 (.I0(x4806), .I1(x4807), .I2(x4808), .O(n8995));
  LUT5 #(.INIT(32'hE81717E8)) lut_n8996 (.I0(x4797), .I1(x4798), .I2(x4799), .I3(n8992), .I4(n8993), .O(n8996));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n8997 (.I0(x4803), .I1(x4804), .I2(x4805), .I3(n8995), .I4(n8996), .O(n8997));
  LUT3 #(.INIT(8'h96)) lut_n8998 (.I0(n8978), .I1(n8981), .I2(n8982), .O(n8998));
  LUT3 #(.INIT(8'hE8)) lut_n8999 (.I0(n8994), .I1(n8997), .I2(n8998), .O(n8999));
  LUT3 #(.INIT(8'hE8)) lut_n9000 (.I0(x4812), .I1(x4813), .I2(x4814), .O(n9000));
  LUT5 #(.INIT(32'hE81717E8)) lut_n9001 (.I0(x4803), .I1(x4804), .I2(x4805), .I3(n8995), .I4(n8996), .O(n9001));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n9002 (.I0(x4809), .I1(x4810), .I2(x4811), .I3(n9000), .I4(n9001), .O(n9002));
  LUT3 #(.INIT(8'hE8)) lut_n9003 (.I0(x4818), .I1(x4819), .I2(x4820), .O(n9003));
  LUT5 #(.INIT(32'hE81717E8)) lut_n9004 (.I0(x4809), .I1(x4810), .I2(x4811), .I3(n9000), .I4(n9001), .O(n9004));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n9005 (.I0(x4815), .I1(x4816), .I2(x4817), .I3(n9003), .I4(n9004), .O(n9005));
  LUT3 #(.INIT(8'h96)) lut_n9006 (.I0(n8994), .I1(n8997), .I2(n8998), .O(n9006));
  LUT3 #(.INIT(8'hE8)) lut_n9007 (.I0(n9002), .I1(n9005), .I2(n9006), .O(n9007));
  LUT3 #(.INIT(8'h96)) lut_n9008 (.I0(n8975), .I1(n8983), .I2(n8984), .O(n9008));
  LUT3 #(.INIT(8'hE8)) lut_n9009 (.I0(n8999), .I1(n9007), .I2(n9008), .O(n9009));
  LUT3 #(.INIT(8'hE8)) lut_n9010 (.I0(x4824), .I1(x4825), .I2(x4826), .O(n9010));
  LUT5 #(.INIT(32'hE81717E8)) lut_n9011 (.I0(x4815), .I1(x4816), .I2(x4817), .I3(n9003), .I4(n9004), .O(n9011));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n9012 (.I0(x4821), .I1(x4822), .I2(x4823), .I3(n9010), .I4(n9011), .O(n9012));
  LUT3 #(.INIT(8'hE8)) lut_n9013 (.I0(x4830), .I1(x4831), .I2(x4832), .O(n9013));
  LUT5 #(.INIT(32'hE81717E8)) lut_n9014 (.I0(x4821), .I1(x4822), .I2(x4823), .I3(n9010), .I4(n9011), .O(n9014));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n9015 (.I0(x4827), .I1(x4828), .I2(x4829), .I3(n9013), .I4(n9014), .O(n9015));
  LUT3 #(.INIT(8'h96)) lut_n9016 (.I0(n9002), .I1(n9005), .I2(n9006), .O(n9016));
  LUT3 #(.INIT(8'hE8)) lut_n9017 (.I0(n9012), .I1(n9015), .I2(n9016), .O(n9017));
  LUT3 #(.INIT(8'hE8)) lut_n9018 (.I0(x4836), .I1(x4837), .I2(x4838), .O(n9018));
  LUT5 #(.INIT(32'hE81717E8)) lut_n9019 (.I0(x4827), .I1(x4828), .I2(x4829), .I3(n9013), .I4(n9014), .O(n9019));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n9020 (.I0(x4833), .I1(x4834), .I2(x4835), .I3(n9018), .I4(n9019), .O(n9020));
  LUT3 #(.INIT(8'hE8)) lut_n9021 (.I0(x4842), .I1(x4843), .I2(x4844), .O(n9021));
  LUT5 #(.INIT(32'hE81717E8)) lut_n9022 (.I0(x4833), .I1(x4834), .I2(x4835), .I3(n9018), .I4(n9019), .O(n9022));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n9023 (.I0(x4839), .I1(x4840), .I2(x4841), .I3(n9021), .I4(n9022), .O(n9023));
  LUT3 #(.INIT(8'h96)) lut_n9024 (.I0(n9012), .I1(n9015), .I2(n9016), .O(n9024));
  LUT3 #(.INIT(8'hE8)) lut_n9025 (.I0(n9020), .I1(n9023), .I2(n9024), .O(n9025));
  LUT3 #(.INIT(8'h96)) lut_n9026 (.I0(n8999), .I1(n9007), .I2(n9008), .O(n9026));
  LUT3 #(.INIT(8'hE8)) lut_n9027 (.I0(n9017), .I1(n9025), .I2(n9026), .O(n9027));
  LUT3 #(.INIT(8'h96)) lut_n9028 (.I0(n8967), .I1(n8985), .I2(n8986), .O(n9028));
  LUT3 #(.INIT(8'hE8)) lut_n9029 (.I0(n9009), .I1(n9027), .I2(n9028), .O(n9029));
  LUT3 #(.INIT(8'hE8)) lut_n9030 (.I0(x4848), .I1(x4849), .I2(x4850), .O(n9030));
  LUT5 #(.INIT(32'hE81717E8)) lut_n9031 (.I0(x4839), .I1(x4840), .I2(x4841), .I3(n9021), .I4(n9022), .O(n9031));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n9032 (.I0(x4845), .I1(x4846), .I2(x4847), .I3(n9030), .I4(n9031), .O(n9032));
  LUT3 #(.INIT(8'hE8)) lut_n9033 (.I0(x4854), .I1(x4855), .I2(x4856), .O(n9033));
  LUT5 #(.INIT(32'hE81717E8)) lut_n9034 (.I0(x4845), .I1(x4846), .I2(x4847), .I3(n9030), .I4(n9031), .O(n9034));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n9035 (.I0(x4851), .I1(x4852), .I2(x4853), .I3(n9033), .I4(n9034), .O(n9035));
  LUT3 #(.INIT(8'h96)) lut_n9036 (.I0(n9020), .I1(n9023), .I2(n9024), .O(n9036));
  LUT3 #(.INIT(8'hE8)) lut_n9037 (.I0(n9032), .I1(n9035), .I2(n9036), .O(n9037));
  LUT3 #(.INIT(8'hE8)) lut_n9038 (.I0(x4860), .I1(x4861), .I2(x4862), .O(n9038));
  LUT5 #(.INIT(32'hE81717E8)) lut_n9039 (.I0(x4851), .I1(x4852), .I2(x4853), .I3(n9033), .I4(n9034), .O(n9039));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n9040 (.I0(x4857), .I1(x4858), .I2(x4859), .I3(n9038), .I4(n9039), .O(n9040));
  LUT3 #(.INIT(8'hE8)) lut_n9041 (.I0(x4866), .I1(x4867), .I2(x4868), .O(n9041));
  LUT5 #(.INIT(32'hE81717E8)) lut_n9042 (.I0(x4857), .I1(x4858), .I2(x4859), .I3(n9038), .I4(n9039), .O(n9042));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n9043 (.I0(x4863), .I1(x4864), .I2(x4865), .I3(n9041), .I4(n9042), .O(n9043));
  LUT3 #(.INIT(8'h96)) lut_n9044 (.I0(n9032), .I1(n9035), .I2(n9036), .O(n9044));
  LUT3 #(.INIT(8'hE8)) lut_n9045 (.I0(n9040), .I1(n9043), .I2(n9044), .O(n9045));
  LUT3 #(.INIT(8'h96)) lut_n9046 (.I0(n9017), .I1(n9025), .I2(n9026), .O(n9046));
  LUT3 #(.INIT(8'hE8)) lut_n9047 (.I0(n9037), .I1(n9045), .I2(n9046), .O(n9047));
  LUT3 #(.INIT(8'hE8)) lut_n9048 (.I0(x4872), .I1(x4873), .I2(x4874), .O(n9048));
  LUT5 #(.INIT(32'hE81717E8)) lut_n9049 (.I0(x4863), .I1(x4864), .I2(x4865), .I3(n9041), .I4(n9042), .O(n9049));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n9050 (.I0(x4869), .I1(x4870), .I2(x4871), .I3(n9048), .I4(n9049), .O(n9050));
  LUT3 #(.INIT(8'hE8)) lut_n9051 (.I0(x4878), .I1(x4879), .I2(x4880), .O(n9051));
  LUT5 #(.INIT(32'hE81717E8)) lut_n9052 (.I0(x4869), .I1(x4870), .I2(x4871), .I3(n9048), .I4(n9049), .O(n9052));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n9053 (.I0(x4875), .I1(x4876), .I2(x4877), .I3(n9051), .I4(n9052), .O(n9053));
  LUT3 #(.INIT(8'h96)) lut_n9054 (.I0(n9040), .I1(n9043), .I2(n9044), .O(n9054));
  LUT3 #(.INIT(8'hE8)) lut_n9055 (.I0(n9050), .I1(n9053), .I2(n9054), .O(n9055));
  LUT3 #(.INIT(8'hE8)) lut_n9056 (.I0(x4884), .I1(x4885), .I2(x4886), .O(n9056));
  LUT5 #(.INIT(32'hE81717E8)) lut_n9057 (.I0(x4875), .I1(x4876), .I2(x4877), .I3(n9051), .I4(n9052), .O(n9057));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n9058 (.I0(x4881), .I1(x4882), .I2(x4883), .I3(n9056), .I4(n9057), .O(n9058));
  LUT3 #(.INIT(8'hE8)) lut_n9059 (.I0(x4890), .I1(x4891), .I2(x4892), .O(n9059));
  LUT5 #(.INIT(32'hE81717E8)) lut_n9060 (.I0(x4881), .I1(x4882), .I2(x4883), .I3(n9056), .I4(n9057), .O(n9060));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n9061 (.I0(x4887), .I1(x4888), .I2(x4889), .I3(n9059), .I4(n9060), .O(n9061));
  LUT3 #(.INIT(8'h96)) lut_n9062 (.I0(n9050), .I1(n9053), .I2(n9054), .O(n9062));
  LUT3 #(.INIT(8'hE8)) lut_n9063 (.I0(n9058), .I1(n9061), .I2(n9062), .O(n9063));
  LUT3 #(.INIT(8'h96)) lut_n9064 (.I0(n9037), .I1(n9045), .I2(n9046), .O(n9064));
  LUT3 #(.INIT(8'hE8)) lut_n9065 (.I0(n9055), .I1(n9063), .I2(n9064), .O(n9065));
  LUT3 #(.INIT(8'h96)) lut_n9066 (.I0(n9009), .I1(n9027), .I2(n9028), .O(n9066));
  LUT3 #(.INIT(8'hE8)) lut_n9067 (.I0(n9047), .I1(n9065), .I2(n9066), .O(n9067));
  LUT3 #(.INIT(8'h96)) lut_n9068 (.I0(n8949), .I1(n8987), .I2(n8988), .O(n9068));
  LUT3 #(.INIT(8'hE8)) lut_n9069 (.I0(n9029), .I1(n9067), .I2(n9068), .O(n9069));
  LUT3 #(.INIT(8'hE8)) lut_n9070 (.I0(x4896), .I1(x4897), .I2(x4898), .O(n9070));
  LUT5 #(.INIT(32'hE81717E8)) lut_n9071 (.I0(x4887), .I1(x4888), .I2(x4889), .I3(n9059), .I4(n9060), .O(n9071));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n9072 (.I0(x4893), .I1(x4894), .I2(x4895), .I3(n9070), .I4(n9071), .O(n9072));
  LUT3 #(.INIT(8'hE8)) lut_n9073 (.I0(x4902), .I1(x4903), .I2(x4904), .O(n9073));
  LUT5 #(.INIT(32'hE81717E8)) lut_n9074 (.I0(x4893), .I1(x4894), .I2(x4895), .I3(n9070), .I4(n9071), .O(n9074));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n9075 (.I0(x4899), .I1(x4900), .I2(x4901), .I3(n9073), .I4(n9074), .O(n9075));
  LUT3 #(.INIT(8'h96)) lut_n9076 (.I0(n9058), .I1(n9061), .I2(n9062), .O(n9076));
  LUT3 #(.INIT(8'hE8)) lut_n9077 (.I0(n9072), .I1(n9075), .I2(n9076), .O(n9077));
  LUT3 #(.INIT(8'hE8)) lut_n9078 (.I0(x4908), .I1(x4909), .I2(x4910), .O(n9078));
  LUT5 #(.INIT(32'hE81717E8)) lut_n9079 (.I0(x4899), .I1(x4900), .I2(x4901), .I3(n9073), .I4(n9074), .O(n9079));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n9080 (.I0(x4905), .I1(x4906), .I2(x4907), .I3(n9078), .I4(n9079), .O(n9080));
  LUT3 #(.INIT(8'hE8)) lut_n9081 (.I0(x4914), .I1(x4915), .I2(x4916), .O(n9081));
  LUT5 #(.INIT(32'hE81717E8)) lut_n9082 (.I0(x4905), .I1(x4906), .I2(x4907), .I3(n9078), .I4(n9079), .O(n9082));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n9083 (.I0(x4911), .I1(x4912), .I2(x4913), .I3(n9081), .I4(n9082), .O(n9083));
  LUT3 #(.INIT(8'h96)) lut_n9084 (.I0(n9072), .I1(n9075), .I2(n9076), .O(n9084));
  LUT3 #(.INIT(8'hE8)) lut_n9085 (.I0(n9080), .I1(n9083), .I2(n9084), .O(n9085));
  LUT3 #(.INIT(8'h96)) lut_n9086 (.I0(n9055), .I1(n9063), .I2(n9064), .O(n9086));
  LUT3 #(.INIT(8'hE8)) lut_n9087 (.I0(n9077), .I1(n9085), .I2(n9086), .O(n9087));
  LUT3 #(.INIT(8'hE8)) lut_n9088 (.I0(x4920), .I1(x4921), .I2(x4922), .O(n9088));
  LUT5 #(.INIT(32'hE81717E8)) lut_n9089 (.I0(x4911), .I1(x4912), .I2(x4913), .I3(n9081), .I4(n9082), .O(n9089));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n9090 (.I0(x4917), .I1(x4918), .I2(x4919), .I3(n9088), .I4(n9089), .O(n9090));
  LUT3 #(.INIT(8'hE8)) lut_n9091 (.I0(x4926), .I1(x4927), .I2(x4928), .O(n9091));
  LUT5 #(.INIT(32'hE81717E8)) lut_n9092 (.I0(x4917), .I1(x4918), .I2(x4919), .I3(n9088), .I4(n9089), .O(n9092));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n9093 (.I0(x4923), .I1(x4924), .I2(x4925), .I3(n9091), .I4(n9092), .O(n9093));
  LUT3 #(.INIT(8'h96)) lut_n9094 (.I0(n9080), .I1(n9083), .I2(n9084), .O(n9094));
  LUT3 #(.INIT(8'hE8)) lut_n9095 (.I0(n9090), .I1(n9093), .I2(n9094), .O(n9095));
  LUT3 #(.INIT(8'hE8)) lut_n9096 (.I0(x4932), .I1(x4933), .I2(x4934), .O(n9096));
  LUT5 #(.INIT(32'hE81717E8)) lut_n9097 (.I0(x4923), .I1(x4924), .I2(x4925), .I3(n9091), .I4(n9092), .O(n9097));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n9098 (.I0(x4929), .I1(x4930), .I2(x4931), .I3(n9096), .I4(n9097), .O(n9098));
  LUT3 #(.INIT(8'hE8)) lut_n9099 (.I0(x4938), .I1(x4939), .I2(x4940), .O(n9099));
  LUT5 #(.INIT(32'hE81717E8)) lut_n9100 (.I0(x4929), .I1(x4930), .I2(x4931), .I3(n9096), .I4(n9097), .O(n9100));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n9101 (.I0(x4935), .I1(x4936), .I2(x4937), .I3(n9099), .I4(n9100), .O(n9101));
  LUT3 #(.INIT(8'h96)) lut_n9102 (.I0(n9090), .I1(n9093), .I2(n9094), .O(n9102));
  LUT3 #(.INIT(8'hE8)) lut_n9103 (.I0(n9098), .I1(n9101), .I2(n9102), .O(n9103));
  LUT3 #(.INIT(8'h96)) lut_n9104 (.I0(n9077), .I1(n9085), .I2(n9086), .O(n9104));
  LUT3 #(.INIT(8'hE8)) lut_n9105 (.I0(n9095), .I1(n9103), .I2(n9104), .O(n9105));
  LUT3 #(.INIT(8'h96)) lut_n9106 (.I0(n9047), .I1(n9065), .I2(n9066), .O(n9106));
  LUT3 #(.INIT(8'hE8)) lut_n9107 (.I0(n9087), .I1(n9105), .I2(n9106), .O(n9107));
  LUT3 #(.INIT(8'hE8)) lut_n9108 (.I0(x4944), .I1(x4945), .I2(x4946), .O(n9108));
  LUT5 #(.INIT(32'hE81717E8)) lut_n9109 (.I0(x4935), .I1(x4936), .I2(x4937), .I3(n9099), .I4(n9100), .O(n9109));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n9110 (.I0(x4941), .I1(x4942), .I2(x4943), .I3(n9108), .I4(n9109), .O(n9110));
  LUT3 #(.INIT(8'hE8)) lut_n9111 (.I0(x4950), .I1(x4951), .I2(x4952), .O(n9111));
  LUT5 #(.INIT(32'hE81717E8)) lut_n9112 (.I0(x4941), .I1(x4942), .I2(x4943), .I3(n9108), .I4(n9109), .O(n9112));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n9113 (.I0(x4947), .I1(x4948), .I2(x4949), .I3(n9111), .I4(n9112), .O(n9113));
  LUT3 #(.INIT(8'h96)) lut_n9114 (.I0(n9098), .I1(n9101), .I2(n9102), .O(n9114));
  LUT3 #(.INIT(8'hE8)) lut_n9115 (.I0(n9110), .I1(n9113), .I2(n9114), .O(n9115));
  LUT3 #(.INIT(8'hE8)) lut_n9116 (.I0(x4956), .I1(x4957), .I2(x4958), .O(n9116));
  LUT5 #(.INIT(32'hE81717E8)) lut_n9117 (.I0(x4947), .I1(x4948), .I2(x4949), .I3(n9111), .I4(n9112), .O(n9117));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n9118 (.I0(x4953), .I1(x4954), .I2(x4955), .I3(n9116), .I4(n9117), .O(n9118));
  LUT3 #(.INIT(8'hE8)) lut_n9119 (.I0(x4962), .I1(x4963), .I2(x4964), .O(n9119));
  LUT5 #(.INIT(32'hE81717E8)) lut_n9120 (.I0(x4953), .I1(x4954), .I2(x4955), .I3(n9116), .I4(n9117), .O(n9120));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n9121 (.I0(x4959), .I1(x4960), .I2(x4961), .I3(n9119), .I4(n9120), .O(n9121));
  LUT3 #(.INIT(8'h96)) lut_n9122 (.I0(n9110), .I1(n9113), .I2(n9114), .O(n9122));
  LUT3 #(.INIT(8'hE8)) lut_n9123 (.I0(n9118), .I1(n9121), .I2(n9122), .O(n9123));
  LUT3 #(.INIT(8'h96)) lut_n9124 (.I0(n9095), .I1(n9103), .I2(n9104), .O(n9124));
  LUT3 #(.INIT(8'hE8)) lut_n9125 (.I0(n9115), .I1(n9123), .I2(n9124), .O(n9125));
  LUT3 #(.INIT(8'hE8)) lut_n9126 (.I0(x4968), .I1(x4969), .I2(x4970), .O(n9126));
  LUT5 #(.INIT(32'hE81717E8)) lut_n9127 (.I0(x4959), .I1(x4960), .I2(x4961), .I3(n9119), .I4(n9120), .O(n9127));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n9128 (.I0(x4965), .I1(x4966), .I2(x4967), .I3(n9126), .I4(n9127), .O(n9128));
  LUT3 #(.INIT(8'hE8)) lut_n9129 (.I0(x4974), .I1(x4975), .I2(x4976), .O(n9129));
  LUT5 #(.INIT(32'hE81717E8)) lut_n9130 (.I0(x4965), .I1(x4966), .I2(x4967), .I3(n9126), .I4(n9127), .O(n9130));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n9131 (.I0(x4971), .I1(x4972), .I2(x4973), .I3(n9129), .I4(n9130), .O(n9131));
  LUT3 #(.INIT(8'h96)) lut_n9132 (.I0(n9118), .I1(n9121), .I2(n9122), .O(n9132));
  LUT3 #(.INIT(8'hE8)) lut_n9133 (.I0(n9128), .I1(n9131), .I2(n9132), .O(n9133));
  LUT3 #(.INIT(8'hE8)) lut_n9134 (.I0(x4980), .I1(x4981), .I2(x4982), .O(n9134));
  LUT5 #(.INIT(32'hE81717E8)) lut_n9135 (.I0(x4971), .I1(x4972), .I2(x4973), .I3(n9129), .I4(n9130), .O(n9135));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n9136 (.I0(x4977), .I1(x4978), .I2(x4979), .I3(n9134), .I4(n9135), .O(n9136));
  LUT3 #(.INIT(8'hE8)) lut_n9137 (.I0(x4986), .I1(x4987), .I2(x4988), .O(n9137));
  LUT5 #(.INIT(32'hE81717E8)) lut_n9138 (.I0(x4977), .I1(x4978), .I2(x4979), .I3(n9134), .I4(n9135), .O(n9138));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n9139 (.I0(x4983), .I1(x4984), .I2(x4985), .I3(n9137), .I4(n9138), .O(n9139));
  LUT3 #(.INIT(8'h96)) lut_n9140 (.I0(n9128), .I1(n9131), .I2(n9132), .O(n9140));
  LUT3 #(.INIT(8'hE8)) lut_n9141 (.I0(n9136), .I1(n9139), .I2(n9140), .O(n9141));
  LUT3 #(.INIT(8'h96)) lut_n9142 (.I0(n9115), .I1(n9123), .I2(n9124), .O(n9142));
  LUT3 #(.INIT(8'hE8)) lut_n9143 (.I0(n9133), .I1(n9141), .I2(n9142), .O(n9143));
  LUT3 #(.INIT(8'h96)) lut_n9144 (.I0(n9087), .I1(n9105), .I2(n9106), .O(n9144));
  LUT3 #(.INIT(8'hE8)) lut_n9145 (.I0(n9125), .I1(n9143), .I2(n9144), .O(n9145));
  LUT3 #(.INIT(8'h96)) lut_n9146 (.I0(n9029), .I1(n9067), .I2(n9068), .O(n9146));
  LUT3 #(.INIT(8'hE8)) lut_n9147 (.I0(n9107), .I1(n9145), .I2(n9146), .O(n9147));
  LUT3 #(.INIT(8'h96)) lut_n9148 (.I0(n8911), .I1(n8989), .I2(n8990), .O(n9148));
  LUT3 #(.INIT(8'hE8)) lut_n9149 (.I0(n9069), .I1(n9147), .I2(n9148), .O(n9149));
  LUT3 #(.INIT(8'h96)) lut_n9150 (.I0(n8669), .I1(n8827), .I2(n8828), .O(n9150));
  LUT3 #(.INIT(8'hE8)) lut_n9151 (.I0(n8991), .I1(n9149), .I2(n9150), .O(n9151));
  LUT3 #(.INIT(8'hE8)) lut_n9152 (.I0(x4992), .I1(x4993), .I2(x4994), .O(n9152));
  LUT5 #(.INIT(32'hE81717E8)) lut_n9153 (.I0(x4983), .I1(x4984), .I2(x4985), .I3(n9137), .I4(n9138), .O(n9153));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n9154 (.I0(x4989), .I1(x4990), .I2(x4991), .I3(n9152), .I4(n9153), .O(n9154));
  LUT3 #(.INIT(8'hE8)) lut_n9155 (.I0(x4998), .I1(x4999), .I2(x5000), .O(n9155));
  LUT5 #(.INIT(32'hE81717E8)) lut_n9156 (.I0(x4989), .I1(x4990), .I2(x4991), .I3(n9152), .I4(n9153), .O(n9156));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n9157 (.I0(x4995), .I1(x4996), .I2(x4997), .I3(n9155), .I4(n9156), .O(n9157));
  LUT3 #(.INIT(8'h96)) lut_n9158 (.I0(n9136), .I1(n9139), .I2(n9140), .O(n9158));
  LUT3 #(.INIT(8'hE8)) lut_n9159 (.I0(n9154), .I1(n9157), .I2(n9158), .O(n9159));
  LUT3 #(.INIT(8'hE8)) lut_n9160 (.I0(x5004), .I1(x5005), .I2(x5006), .O(n9160));
  LUT5 #(.INIT(32'hE81717E8)) lut_n9161 (.I0(x4995), .I1(x4996), .I2(x4997), .I3(n9155), .I4(n9156), .O(n9161));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n9162 (.I0(x5001), .I1(x5002), .I2(x5003), .I3(n9160), .I4(n9161), .O(n9162));
  LUT3 #(.INIT(8'hE8)) lut_n9163 (.I0(x5010), .I1(x5011), .I2(x5012), .O(n9163));
  LUT5 #(.INIT(32'hE81717E8)) lut_n9164 (.I0(x5001), .I1(x5002), .I2(x5003), .I3(n9160), .I4(n9161), .O(n9164));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n9165 (.I0(x5007), .I1(x5008), .I2(x5009), .I3(n9163), .I4(n9164), .O(n9165));
  LUT3 #(.INIT(8'h96)) lut_n9166 (.I0(n9154), .I1(n9157), .I2(n9158), .O(n9166));
  LUT3 #(.INIT(8'hE8)) lut_n9167 (.I0(n9162), .I1(n9165), .I2(n9166), .O(n9167));
  LUT3 #(.INIT(8'h96)) lut_n9168 (.I0(n9133), .I1(n9141), .I2(n9142), .O(n9168));
  LUT3 #(.INIT(8'hE8)) lut_n9169 (.I0(n9159), .I1(n9167), .I2(n9168), .O(n9169));
  LUT3 #(.INIT(8'hE8)) lut_n9170 (.I0(x5016), .I1(x5017), .I2(x5018), .O(n9170));
  LUT5 #(.INIT(32'hE81717E8)) lut_n9171 (.I0(x5007), .I1(x5008), .I2(x5009), .I3(n9163), .I4(n9164), .O(n9171));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n9172 (.I0(x5013), .I1(x5014), .I2(x5015), .I3(n9170), .I4(n9171), .O(n9172));
  LUT3 #(.INIT(8'hE8)) lut_n9173 (.I0(x5022), .I1(x5023), .I2(x5024), .O(n9173));
  LUT5 #(.INIT(32'hE81717E8)) lut_n9174 (.I0(x5013), .I1(x5014), .I2(x5015), .I3(n9170), .I4(n9171), .O(n9174));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n9175 (.I0(x5019), .I1(x5020), .I2(x5021), .I3(n9173), .I4(n9174), .O(n9175));
  LUT3 #(.INIT(8'h96)) lut_n9176 (.I0(n9162), .I1(n9165), .I2(n9166), .O(n9176));
  LUT3 #(.INIT(8'hE8)) lut_n9177 (.I0(n9172), .I1(n9175), .I2(n9176), .O(n9177));
  LUT3 #(.INIT(8'h96)) lut_n9178 (.I0(x0), .I1(x1), .I2(x2), .O(n9178));
  LUT3 #(.INIT(8'h96)) lut_n9179 (.I0(x6), .I1(x7), .I2(x8), .O(n9179));
  LUT5 #(.INIT(32'hFF969600)) lut_n9180 (.I0(x3), .I1(x4), .I2(x5), .I3(n9178), .I4(n9179), .O(n9180));
  LUT3 #(.INIT(8'h96)) lut_n9181 (.I0(x12), .I1(x13), .I2(x14), .O(n9181));
  LUT5 #(.INIT(32'h96696996)) lut_n9182 (.I0(x3), .I1(x4), .I2(x5), .I3(n9178), .I4(n9179), .O(n9182));
  LUT5 #(.INIT(32'hFF969600)) lut_n9183 (.I0(x9), .I1(x10), .I2(x11), .I3(n9181), .I4(n9182), .O(n9183));
  LUT5 #(.INIT(32'hE81717E8)) lut_n9184 (.I0(x5019), .I1(x5020), .I2(x5021), .I3(n9173), .I4(n9174), .O(n9184));
  LUT3 #(.INIT(8'hE8)) lut_n9185 (.I0(n9180), .I1(n9183), .I2(n9184), .O(n9185));
  LUT3 #(.INIT(8'h96)) lut_n9186 (.I0(x18), .I1(x19), .I2(x20), .O(n9186));
  LUT5 #(.INIT(32'h96696996)) lut_n9187 (.I0(x9), .I1(x10), .I2(x11), .I3(n9181), .I4(n9182), .O(n9187));
  LUT5 #(.INIT(32'hFF969600)) lut_n9188 (.I0(x15), .I1(x16), .I2(x17), .I3(n9186), .I4(n9187), .O(n9188));
  LUT3 #(.INIT(8'h96)) lut_n9189 (.I0(x24), .I1(x25), .I2(x26), .O(n9189));
  LUT5 #(.INIT(32'h96696996)) lut_n9190 (.I0(x15), .I1(x16), .I2(x17), .I3(n9186), .I4(n9187), .O(n9190));
  LUT5 #(.INIT(32'hFF969600)) lut_n9191 (.I0(x21), .I1(x22), .I2(x23), .I3(n9189), .I4(n9190), .O(n9191));
  LUT3 #(.INIT(8'h96)) lut_n9192 (.I0(n9180), .I1(n9183), .I2(n9184), .O(n9192));
  LUT3 #(.INIT(8'hE8)) lut_n9193 (.I0(n9188), .I1(n9191), .I2(n9192), .O(n9193));
  LUT3 #(.INIT(8'h96)) lut_n9194 (.I0(n9172), .I1(n9175), .I2(n9176), .O(n9194));
  LUT3 #(.INIT(8'hE8)) lut_n9195 (.I0(n9185), .I1(n9193), .I2(n9194), .O(n9195));
  LUT3 #(.INIT(8'h96)) lut_n9196 (.I0(n9159), .I1(n9167), .I2(n9168), .O(n9196));
  LUT3 #(.INIT(8'hE8)) lut_n9197 (.I0(n9177), .I1(n9195), .I2(n9196), .O(n9197));
  LUT3 #(.INIT(8'h96)) lut_n9198 (.I0(n9125), .I1(n9143), .I2(n9144), .O(n9198));
  LUT3 #(.INIT(8'hE8)) lut_n9199 (.I0(n9169), .I1(n9197), .I2(n9198), .O(n9199));
  LUT3 #(.INIT(8'h96)) lut_n9200 (.I0(x27), .I1(x28), .I2(x29), .O(n9200));
  LUT5 #(.INIT(32'h96696996)) lut_n9201 (.I0(x21), .I1(x22), .I2(x23), .I3(n9189), .I4(n9190), .O(n9201));
  LUT5 #(.INIT(32'hFF969600)) lut_n9202 (.I0(x30), .I1(x31), .I2(x32), .I3(n9200), .I4(n9201), .O(n9202));
  LUT3 #(.INIT(8'h96)) lut_n9203 (.I0(x36), .I1(x37), .I2(x38), .O(n9203));
  LUT5 #(.INIT(32'h96696996)) lut_n9204 (.I0(x30), .I1(x31), .I2(x32), .I3(n9200), .I4(n9201), .O(n9204));
  LUT5 #(.INIT(32'hFF969600)) lut_n9205 (.I0(x33), .I1(x34), .I2(x35), .I3(n9203), .I4(n9204), .O(n9205));
  LUT3 #(.INIT(8'h96)) lut_n9206 (.I0(n9188), .I1(n9191), .I2(n9192), .O(n9206));
  LUT3 #(.INIT(8'hE8)) lut_n9207 (.I0(n9202), .I1(n9205), .I2(n9206), .O(n9207));
  LUT3 #(.INIT(8'h96)) lut_n9208 (.I0(x42), .I1(x43), .I2(x44), .O(n9208));
  LUT5 #(.INIT(32'h96696996)) lut_n9209 (.I0(x33), .I1(x34), .I2(x35), .I3(n9203), .I4(n9204), .O(n9209));
  LUT5 #(.INIT(32'hFF969600)) lut_n9210 (.I0(x39), .I1(x40), .I2(x41), .I3(n9208), .I4(n9209), .O(n9210));
  LUT3 #(.INIT(8'h96)) lut_n9211 (.I0(x48), .I1(x49), .I2(x50), .O(n9211));
  LUT5 #(.INIT(32'h96696996)) lut_n9212 (.I0(x39), .I1(x40), .I2(x41), .I3(n9208), .I4(n9209), .O(n9212));
  LUT5 #(.INIT(32'hFF969600)) lut_n9213 (.I0(x45), .I1(x46), .I2(x47), .I3(n9211), .I4(n9212), .O(n9213));
  LUT3 #(.INIT(8'h96)) lut_n9214 (.I0(n9202), .I1(n9205), .I2(n9206), .O(n9214));
  LUT3 #(.INIT(8'hE8)) lut_n9215 (.I0(n9210), .I1(n9213), .I2(n9214), .O(n9215));
  LUT3 #(.INIT(8'h96)) lut_n9216 (.I0(n9185), .I1(n9193), .I2(n9194), .O(n9216));
  LUT3 #(.INIT(8'hE8)) lut_n9217 (.I0(n9207), .I1(n9215), .I2(n9216), .O(n9217));
  LUT3 #(.INIT(8'h96)) lut_n9218 (.I0(x54), .I1(x55), .I2(x56), .O(n9218));
  LUT5 #(.INIT(32'h96696996)) lut_n9219 (.I0(x45), .I1(x46), .I2(x47), .I3(n9211), .I4(n9212), .O(n9219));
  LUT5 #(.INIT(32'hFF969600)) lut_n9220 (.I0(x51), .I1(x52), .I2(x53), .I3(n9218), .I4(n9219), .O(n9220));
  LUT3 #(.INIT(8'h96)) lut_n9221 (.I0(x60), .I1(x61), .I2(x62), .O(n9221));
  LUT5 #(.INIT(32'h96696996)) lut_n9222 (.I0(x51), .I1(x52), .I2(x53), .I3(n9218), .I4(n9219), .O(n9222));
  LUT5 #(.INIT(32'hFF969600)) lut_n9223 (.I0(x57), .I1(x58), .I2(x59), .I3(n9221), .I4(n9222), .O(n9223));
  LUT3 #(.INIT(8'h96)) lut_n9224 (.I0(n9210), .I1(n9213), .I2(n9214), .O(n9224));
  LUT3 #(.INIT(8'hE8)) lut_n9225 (.I0(n9220), .I1(n9223), .I2(n9224), .O(n9225));
  LUT3 #(.INIT(8'h96)) lut_n9226 (.I0(x66), .I1(x67), .I2(x68), .O(n9226));
  LUT5 #(.INIT(32'h96696996)) lut_n9227 (.I0(x57), .I1(x58), .I2(x59), .I3(n9221), .I4(n9222), .O(n9227));
  LUT5 #(.INIT(32'hFF969600)) lut_n9228 (.I0(x63), .I1(x64), .I2(x65), .I3(n9226), .I4(n9227), .O(n9228));
  LUT3 #(.INIT(8'h96)) lut_n9229 (.I0(x72), .I1(x73), .I2(x74), .O(n9229));
  LUT5 #(.INIT(32'h96696996)) lut_n9230 (.I0(x63), .I1(x64), .I2(x65), .I3(n9226), .I4(n9227), .O(n9230));
  LUT5 #(.INIT(32'hFF969600)) lut_n9231 (.I0(x69), .I1(x70), .I2(x71), .I3(n9229), .I4(n9230), .O(n9231));
  LUT3 #(.INIT(8'h96)) lut_n9232 (.I0(n9220), .I1(n9223), .I2(n9224), .O(n9232));
  LUT3 #(.INIT(8'hE8)) lut_n9233 (.I0(n9228), .I1(n9231), .I2(n9232), .O(n9233));
  LUT3 #(.INIT(8'h96)) lut_n9234 (.I0(n9207), .I1(n9215), .I2(n9216), .O(n9234));
  LUT3 #(.INIT(8'hE8)) lut_n9235 (.I0(n9225), .I1(n9233), .I2(n9234), .O(n9235));
  LUT3 #(.INIT(8'h96)) lut_n9236 (.I0(n9177), .I1(n9195), .I2(n9196), .O(n9236));
  LUT3 #(.INIT(8'hE8)) lut_n9237 (.I0(n9217), .I1(n9235), .I2(n9236), .O(n9237));
  LUT3 #(.INIT(8'h96)) lut_n9238 (.I0(x78), .I1(x79), .I2(x80), .O(n9238));
  LUT5 #(.INIT(32'h96696996)) lut_n9239 (.I0(x69), .I1(x70), .I2(x71), .I3(n9229), .I4(n9230), .O(n9239));
  LUT5 #(.INIT(32'hFF969600)) lut_n9240 (.I0(x75), .I1(x76), .I2(x77), .I3(n9238), .I4(n9239), .O(n9240));
  LUT3 #(.INIT(8'h96)) lut_n9241 (.I0(x84), .I1(x85), .I2(x86), .O(n9241));
  LUT5 #(.INIT(32'h96696996)) lut_n9242 (.I0(x75), .I1(x76), .I2(x77), .I3(n9238), .I4(n9239), .O(n9242));
  LUT5 #(.INIT(32'hFF969600)) lut_n9243 (.I0(x81), .I1(x82), .I2(x83), .I3(n9241), .I4(n9242), .O(n9243));
  LUT3 #(.INIT(8'h96)) lut_n9244 (.I0(n9228), .I1(n9231), .I2(n9232), .O(n9244));
  LUT3 #(.INIT(8'hE8)) lut_n9245 (.I0(n9240), .I1(n9243), .I2(n9244), .O(n9245));
  LUT3 #(.INIT(8'h96)) lut_n9246 (.I0(x90), .I1(x91), .I2(x92), .O(n9246));
  LUT5 #(.INIT(32'h96696996)) lut_n9247 (.I0(x81), .I1(x82), .I2(x83), .I3(n9241), .I4(n9242), .O(n9247));
  LUT5 #(.INIT(32'hFF969600)) lut_n9248 (.I0(x87), .I1(x88), .I2(x89), .I3(n9246), .I4(n9247), .O(n9248));
  LUT3 #(.INIT(8'h96)) lut_n9249 (.I0(x96), .I1(x97), .I2(x98), .O(n9249));
  LUT5 #(.INIT(32'h96696996)) lut_n9250 (.I0(x87), .I1(x88), .I2(x89), .I3(n9246), .I4(n9247), .O(n9250));
  LUT5 #(.INIT(32'hFF969600)) lut_n9251 (.I0(x93), .I1(x94), .I2(x95), .I3(n9249), .I4(n9250), .O(n9251));
  LUT3 #(.INIT(8'h96)) lut_n9252 (.I0(n9240), .I1(n9243), .I2(n9244), .O(n9252));
  LUT3 #(.INIT(8'hE8)) lut_n9253 (.I0(n9248), .I1(n9251), .I2(n9252), .O(n9253));
  LUT3 #(.INIT(8'h96)) lut_n9254 (.I0(n9225), .I1(n9233), .I2(n9234), .O(n9254));
  LUT3 #(.INIT(8'hE8)) lut_n9255 (.I0(n9245), .I1(n9253), .I2(n9254), .O(n9255));
  LUT3 #(.INIT(8'h96)) lut_n9256 (.I0(x102), .I1(x103), .I2(x104), .O(n9256));
  LUT5 #(.INIT(32'h96696996)) lut_n9257 (.I0(x93), .I1(x94), .I2(x95), .I3(n9249), .I4(n9250), .O(n9257));
  LUT5 #(.INIT(32'hFF969600)) lut_n9258 (.I0(x99), .I1(x100), .I2(x101), .I3(n9256), .I4(n9257), .O(n9258));
  LUT3 #(.INIT(8'h96)) lut_n9259 (.I0(x108), .I1(x109), .I2(x110), .O(n9259));
  LUT5 #(.INIT(32'h96696996)) lut_n9260 (.I0(x99), .I1(x100), .I2(x101), .I3(n9256), .I4(n9257), .O(n9260));
  LUT5 #(.INIT(32'hFF969600)) lut_n9261 (.I0(x105), .I1(x106), .I2(x107), .I3(n9259), .I4(n9260), .O(n9261));
  LUT3 #(.INIT(8'h96)) lut_n9262 (.I0(n9248), .I1(n9251), .I2(n9252), .O(n9262));
  LUT3 #(.INIT(8'hE8)) lut_n9263 (.I0(n9258), .I1(n9261), .I2(n9262), .O(n9263));
  LUT3 #(.INIT(8'h96)) lut_n9264 (.I0(x114), .I1(x115), .I2(x116), .O(n9264));
  LUT5 #(.INIT(32'h96696996)) lut_n9265 (.I0(x105), .I1(x106), .I2(x107), .I3(n9259), .I4(n9260), .O(n9265));
  LUT5 #(.INIT(32'hFF969600)) lut_n9266 (.I0(x111), .I1(x112), .I2(x113), .I3(n9264), .I4(n9265), .O(n9266));
  LUT3 #(.INIT(8'h96)) lut_n9267 (.I0(x120), .I1(x121), .I2(x122), .O(n9267));
  LUT5 #(.INIT(32'h96696996)) lut_n9268 (.I0(x111), .I1(x112), .I2(x113), .I3(n9264), .I4(n9265), .O(n9268));
  LUT5 #(.INIT(32'hFF969600)) lut_n9269 (.I0(x117), .I1(x118), .I2(x119), .I3(n9267), .I4(n9268), .O(n9269));
  LUT3 #(.INIT(8'h96)) lut_n9270 (.I0(n9258), .I1(n9261), .I2(n9262), .O(n9270));
  LUT3 #(.INIT(8'hE8)) lut_n9271 (.I0(n9266), .I1(n9269), .I2(n9270), .O(n9271));
  LUT3 #(.INIT(8'h96)) lut_n9272 (.I0(n9245), .I1(n9253), .I2(n9254), .O(n9272));
  LUT3 #(.INIT(8'hE8)) lut_n9273 (.I0(n9263), .I1(n9271), .I2(n9272), .O(n9273));
  LUT3 #(.INIT(8'h96)) lut_n9274 (.I0(n9217), .I1(n9235), .I2(n9236), .O(n9274));
  LUT3 #(.INIT(8'hE8)) lut_n9275 (.I0(n9255), .I1(n9273), .I2(n9274), .O(n9275));
  LUT3 #(.INIT(8'h96)) lut_n9276 (.I0(n9169), .I1(n9197), .I2(n9198), .O(n9276));
  LUT3 #(.INIT(8'hE8)) lut_n9277 (.I0(n9237), .I1(n9275), .I2(n9276), .O(n9277));
  LUT3 #(.INIT(8'h96)) lut_n9278 (.I0(n9107), .I1(n9145), .I2(n9146), .O(n9278));
  LUT3 #(.INIT(8'hE8)) lut_n9279 (.I0(n9199), .I1(n9277), .I2(n9278), .O(n9279));
  LUT3 #(.INIT(8'h96)) lut_n9280 (.I0(x126), .I1(x127), .I2(x128), .O(n9280));
  LUT5 #(.INIT(32'h96696996)) lut_n9281 (.I0(x117), .I1(x118), .I2(x119), .I3(n9267), .I4(n9268), .O(n9281));
  LUT5 #(.INIT(32'hFF969600)) lut_n9282 (.I0(x123), .I1(x124), .I2(x125), .I3(n9280), .I4(n9281), .O(n9282));
  LUT3 #(.INIT(8'h96)) lut_n9283 (.I0(x132), .I1(x133), .I2(x134), .O(n9283));
  LUT5 #(.INIT(32'h96696996)) lut_n9284 (.I0(x123), .I1(x124), .I2(x125), .I3(n9280), .I4(n9281), .O(n9284));
  LUT5 #(.INIT(32'hFF969600)) lut_n9285 (.I0(x129), .I1(x130), .I2(x131), .I3(n9283), .I4(n9284), .O(n9285));
  LUT3 #(.INIT(8'h96)) lut_n9286 (.I0(n9266), .I1(n9269), .I2(n9270), .O(n9286));
  LUT3 #(.INIT(8'hE8)) lut_n9287 (.I0(n9282), .I1(n9285), .I2(n9286), .O(n9287));
  LUT3 #(.INIT(8'h96)) lut_n9288 (.I0(x138), .I1(x139), .I2(x140), .O(n9288));
  LUT5 #(.INIT(32'h96696996)) lut_n9289 (.I0(x129), .I1(x130), .I2(x131), .I3(n9283), .I4(n9284), .O(n9289));
  LUT5 #(.INIT(32'hFF969600)) lut_n9290 (.I0(x135), .I1(x136), .I2(x137), .I3(n9288), .I4(n9289), .O(n9290));
  LUT3 #(.INIT(8'h96)) lut_n9291 (.I0(x144), .I1(x145), .I2(x146), .O(n9291));
  LUT5 #(.INIT(32'h96696996)) lut_n9292 (.I0(x135), .I1(x136), .I2(x137), .I3(n9288), .I4(n9289), .O(n9292));
  LUT5 #(.INIT(32'hFF969600)) lut_n9293 (.I0(x141), .I1(x142), .I2(x143), .I3(n9291), .I4(n9292), .O(n9293));
  LUT3 #(.INIT(8'h96)) lut_n9294 (.I0(n9282), .I1(n9285), .I2(n9286), .O(n9294));
  LUT3 #(.INIT(8'hE8)) lut_n9295 (.I0(n9290), .I1(n9293), .I2(n9294), .O(n9295));
  LUT3 #(.INIT(8'h96)) lut_n9296 (.I0(n9263), .I1(n9271), .I2(n9272), .O(n9296));
  LUT3 #(.INIT(8'hE8)) lut_n9297 (.I0(n9287), .I1(n9295), .I2(n9296), .O(n9297));
  LUT3 #(.INIT(8'h96)) lut_n9298 (.I0(x150), .I1(x151), .I2(x152), .O(n9298));
  LUT5 #(.INIT(32'h96696996)) lut_n9299 (.I0(x141), .I1(x142), .I2(x143), .I3(n9291), .I4(n9292), .O(n9299));
  LUT5 #(.INIT(32'hFF969600)) lut_n9300 (.I0(x147), .I1(x148), .I2(x149), .I3(n9298), .I4(n9299), .O(n9300));
  LUT3 #(.INIT(8'h96)) lut_n9301 (.I0(x156), .I1(x157), .I2(x158), .O(n9301));
  LUT5 #(.INIT(32'h96696996)) lut_n9302 (.I0(x147), .I1(x148), .I2(x149), .I3(n9298), .I4(n9299), .O(n9302));
  LUT5 #(.INIT(32'hFF969600)) lut_n9303 (.I0(x153), .I1(x154), .I2(x155), .I3(n9301), .I4(n9302), .O(n9303));
  LUT3 #(.INIT(8'h96)) lut_n9304 (.I0(n9290), .I1(n9293), .I2(n9294), .O(n9304));
  LUT3 #(.INIT(8'hE8)) lut_n9305 (.I0(n9300), .I1(n9303), .I2(n9304), .O(n9305));
  LUT3 #(.INIT(8'h96)) lut_n9306 (.I0(x162), .I1(x163), .I2(x164), .O(n9306));
  LUT5 #(.INIT(32'h96696996)) lut_n9307 (.I0(x153), .I1(x154), .I2(x155), .I3(n9301), .I4(n9302), .O(n9307));
  LUT5 #(.INIT(32'hFF969600)) lut_n9308 (.I0(x159), .I1(x160), .I2(x161), .I3(n9306), .I4(n9307), .O(n9308));
  LUT3 #(.INIT(8'h96)) lut_n9309 (.I0(x168), .I1(x169), .I2(x170), .O(n9309));
  LUT5 #(.INIT(32'h96696996)) lut_n9310 (.I0(x159), .I1(x160), .I2(x161), .I3(n9306), .I4(n9307), .O(n9310));
  LUT5 #(.INIT(32'hFF969600)) lut_n9311 (.I0(x165), .I1(x166), .I2(x167), .I3(n9309), .I4(n9310), .O(n9311));
  LUT3 #(.INIT(8'h96)) lut_n9312 (.I0(n9300), .I1(n9303), .I2(n9304), .O(n9312));
  LUT3 #(.INIT(8'hE8)) lut_n9313 (.I0(n9308), .I1(n9311), .I2(n9312), .O(n9313));
  LUT3 #(.INIT(8'h96)) lut_n9314 (.I0(n9287), .I1(n9295), .I2(n9296), .O(n9314));
  LUT3 #(.INIT(8'hE8)) lut_n9315 (.I0(n9305), .I1(n9313), .I2(n9314), .O(n9315));
  LUT3 #(.INIT(8'h96)) lut_n9316 (.I0(n9255), .I1(n9273), .I2(n9274), .O(n9316));
  LUT3 #(.INIT(8'hE8)) lut_n9317 (.I0(n9297), .I1(n9315), .I2(n9316), .O(n9317));
  LUT3 #(.INIT(8'h96)) lut_n9318 (.I0(x174), .I1(x175), .I2(x176), .O(n9318));
  LUT5 #(.INIT(32'h96696996)) lut_n9319 (.I0(x165), .I1(x166), .I2(x167), .I3(n9309), .I4(n9310), .O(n9319));
  LUT5 #(.INIT(32'hFF969600)) lut_n9320 (.I0(x171), .I1(x172), .I2(x173), .I3(n9318), .I4(n9319), .O(n9320));
  LUT3 #(.INIT(8'h96)) lut_n9321 (.I0(x180), .I1(x181), .I2(x182), .O(n9321));
  LUT5 #(.INIT(32'h96696996)) lut_n9322 (.I0(x171), .I1(x172), .I2(x173), .I3(n9318), .I4(n9319), .O(n9322));
  LUT5 #(.INIT(32'hFF969600)) lut_n9323 (.I0(x177), .I1(x178), .I2(x179), .I3(n9321), .I4(n9322), .O(n9323));
  LUT3 #(.INIT(8'h96)) lut_n9324 (.I0(n9308), .I1(n9311), .I2(n9312), .O(n9324));
  LUT3 #(.INIT(8'hE8)) lut_n9325 (.I0(n9320), .I1(n9323), .I2(n9324), .O(n9325));
  LUT3 #(.INIT(8'h96)) lut_n9326 (.I0(x186), .I1(x187), .I2(x188), .O(n9326));
  LUT5 #(.INIT(32'h96696996)) lut_n9327 (.I0(x177), .I1(x178), .I2(x179), .I3(n9321), .I4(n9322), .O(n9327));
  LUT5 #(.INIT(32'hFF969600)) lut_n9328 (.I0(x183), .I1(x184), .I2(x185), .I3(n9326), .I4(n9327), .O(n9328));
  LUT3 #(.INIT(8'h96)) lut_n9329 (.I0(x192), .I1(x193), .I2(x194), .O(n9329));
  LUT5 #(.INIT(32'h96696996)) lut_n9330 (.I0(x183), .I1(x184), .I2(x185), .I3(n9326), .I4(n9327), .O(n9330));
  LUT5 #(.INIT(32'hFF969600)) lut_n9331 (.I0(x189), .I1(x190), .I2(x191), .I3(n9329), .I4(n9330), .O(n9331));
  LUT3 #(.INIT(8'h96)) lut_n9332 (.I0(n9320), .I1(n9323), .I2(n9324), .O(n9332));
  LUT3 #(.INIT(8'hE8)) lut_n9333 (.I0(n9328), .I1(n9331), .I2(n9332), .O(n9333));
  LUT3 #(.INIT(8'h96)) lut_n9334 (.I0(n9305), .I1(n9313), .I2(n9314), .O(n9334));
  LUT3 #(.INIT(8'hE8)) lut_n9335 (.I0(n9325), .I1(n9333), .I2(n9334), .O(n9335));
  LUT3 #(.INIT(8'h96)) lut_n9336 (.I0(x198), .I1(x199), .I2(x200), .O(n9336));
  LUT5 #(.INIT(32'h96696996)) lut_n9337 (.I0(x189), .I1(x190), .I2(x191), .I3(n9329), .I4(n9330), .O(n9337));
  LUT5 #(.INIT(32'hFF969600)) lut_n9338 (.I0(x195), .I1(x196), .I2(x197), .I3(n9336), .I4(n9337), .O(n9338));
  LUT3 #(.INIT(8'h96)) lut_n9339 (.I0(x204), .I1(x205), .I2(x206), .O(n9339));
  LUT5 #(.INIT(32'h96696996)) lut_n9340 (.I0(x195), .I1(x196), .I2(x197), .I3(n9336), .I4(n9337), .O(n9340));
  LUT5 #(.INIT(32'hFF969600)) lut_n9341 (.I0(x201), .I1(x202), .I2(x203), .I3(n9339), .I4(n9340), .O(n9341));
  LUT3 #(.INIT(8'h96)) lut_n9342 (.I0(n9328), .I1(n9331), .I2(n9332), .O(n9342));
  LUT3 #(.INIT(8'hE8)) lut_n9343 (.I0(n9338), .I1(n9341), .I2(n9342), .O(n9343));
  LUT3 #(.INIT(8'h96)) lut_n9344 (.I0(x210), .I1(x211), .I2(x212), .O(n9344));
  LUT5 #(.INIT(32'h96696996)) lut_n9345 (.I0(x201), .I1(x202), .I2(x203), .I3(n9339), .I4(n9340), .O(n9345));
  LUT5 #(.INIT(32'hFF969600)) lut_n9346 (.I0(x207), .I1(x208), .I2(x209), .I3(n9344), .I4(n9345), .O(n9346));
  LUT3 #(.INIT(8'h96)) lut_n9347 (.I0(x216), .I1(x217), .I2(x218), .O(n9347));
  LUT5 #(.INIT(32'h96696996)) lut_n9348 (.I0(x207), .I1(x208), .I2(x209), .I3(n9344), .I4(n9345), .O(n9348));
  LUT5 #(.INIT(32'hFF969600)) lut_n9349 (.I0(x213), .I1(x214), .I2(x215), .I3(n9347), .I4(n9348), .O(n9349));
  LUT3 #(.INIT(8'h96)) lut_n9350 (.I0(n9338), .I1(n9341), .I2(n9342), .O(n9350));
  LUT3 #(.INIT(8'hE8)) lut_n9351 (.I0(n9346), .I1(n9349), .I2(n9350), .O(n9351));
  LUT3 #(.INIT(8'h96)) lut_n9352 (.I0(n9325), .I1(n9333), .I2(n9334), .O(n9352));
  LUT3 #(.INIT(8'hE8)) lut_n9353 (.I0(n9343), .I1(n9351), .I2(n9352), .O(n9353));
  LUT3 #(.INIT(8'h96)) lut_n9354 (.I0(n9297), .I1(n9315), .I2(n9316), .O(n9354));
  LUT3 #(.INIT(8'hE8)) lut_n9355 (.I0(n9335), .I1(n9353), .I2(n9354), .O(n9355));
  LUT3 #(.INIT(8'h96)) lut_n9356 (.I0(n9237), .I1(n9275), .I2(n9276), .O(n9356));
  LUT3 #(.INIT(8'hE8)) lut_n9357 (.I0(n9317), .I1(n9355), .I2(n9356), .O(n9357));
  LUT3 #(.INIT(8'h96)) lut_n9358 (.I0(x222), .I1(x223), .I2(x224), .O(n9358));
  LUT5 #(.INIT(32'h96696996)) lut_n9359 (.I0(x213), .I1(x214), .I2(x215), .I3(n9347), .I4(n9348), .O(n9359));
  LUT5 #(.INIT(32'hFF969600)) lut_n9360 (.I0(x219), .I1(x220), .I2(x221), .I3(n9358), .I4(n9359), .O(n9360));
  LUT3 #(.INIT(8'h96)) lut_n9361 (.I0(x228), .I1(x229), .I2(x230), .O(n9361));
  LUT5 #(.INIT(32'h96696996)) lut_n9362 (.I0(x219), .I1(x220), .I2(x221), .I3(n9358), .I4(n9359), .O(n9362));
  LUT5 #(.INIT(32'hFF969600)) lut_n9363 (.I0(x225), .I1(x226), .I2(x227), .I3(n9361), .I4(n9362), .O(n9363));
  LUT3 #(.INIT(8'h96)) lut_n9364 (.I0(n9346), .I1(n9349), .I2(n9350), .O(n9364));
  LUT3 #(.INIT(8'hE8)) lut_n9365 (.I0(n9360), .I1(n9363), .I2(n9364), .O(n9365));
  LUT3 #(.INIT(8'h96)) lut_n9366 (.I0(x234), .I1(x235), .I2(x236), .O(n9366));
  LUT5 #(.INIT(32'h96696996)) lut_n9367 (.I0(x225), .I1(x226), .I2(x227), .I3(n9361), .I4(n9362), .O(n9367));
  LUT5 #(.INIT(32'hFF969600)) lut_n9368 (.I0(x231), .I1(x232), .I2(x233), .I3(n9366), .I4(n9367), .O(n9368));
  LUT3 #(.INIT(8'h96)) lut_n9369 (.I0(x240), .I1(x241), .I2(x242), .O(n9369));
  LUT5 #(.INIT(32'h96696996)) lut_n9370 (.I0(x231), .I1(x232), .I2(x233), .I3(n9366), .I4(n9367), .O(n9370));
  LUT5 #(.INIT(32'hFF969600)) lut_n9371 (.I0(x237), .I1(x238), .I2(x239), .I3(n9369), .I4(n9370), .O(n9371));
  LUT3 #(.INIT(8'h96)) lut_n9372 (.I0(n9360), .I1(n9363), .I2(n9364), .O(n9372));
  LUT3 #(.INIT(8'hE8)) lut_n9373 (.I0(n9368), .I1(n9371), .I2(n9372), .O(n9373));
  LUT3 #(.INIT(8'h96)) lut_n9374 (.I0(n9343), .I1(n9351), .I2(n9352), .O(n9374));
  LUT3 #(.INIT(8'hE8)) lut_n9375 (.I0(n9365), .I1(n9373), .I2(n9374), .O(n9375));
  LUT3 #(.INIT(8'h96)) lut_n9376 (.I0(x246), .I1(x247), .I2(x248), .O(n9376));
  LUT5 #(.INIT(32'h96696996)) lut_n9377 (.I0(x237), .I1(x238), .I2(x239), .I3(n9369), .I4(n9370), .O(n9377));
  LUT5 #(.INIT(32'hFF969600)) lut_n9378 (.I0(x243), .I1(x244), .I2(x245), .I3(n9376), .I4(n9377), .O(n9378));
  LUT3 #(.INIT(8'h96)) lut_n9379 (.I0(x252), .I1(x253), .I2(x254), .O(n9379));
  LUT5 #(.INIT(32'h96696996)) lut_n9380 (.I0(x243), .I1(x244), .I2(x245), .I3(n9376), .I4(n9377), .O(n9380));
  LUT5 #(.INIT(32'hFF969600)) lut_n9381 (.I0(x249), .I1(x250), .I2(x251), .I3(n9379), .I4(n9380), .O(n9381));
  LUT3 #(.INIT(8'h96)) lut_n9382 (.I0(n9368), .I1(n9371), .I2(n9372), .O(n9382));
  LUT3 #(.INIT(8'hE8)) lut_n9383 (.I0(n9378), .I1(n9381), .I2(n9382), .O(n9383));
  LUT3 #(.INIT(8'h96)) lut_n9384 (.I0(x258), .I1(x259), .I2(x260), .O(n9384));
  LUT5 #(.INIT(32'h96696996)) lut_n9385 (.I0(x249), .I1(x250), .I2(x251), .I3(n9379), .I4(n9380), .O(n9385));
  LUT5 #(.INIT(32'hFF969600)) lut_n9386 (.I0(x255), .I1(x256), .I2(x257), .I3(n9384), .I4(n9385), .O(n9386));
  LUT3 #(.INIT(8'h96)) lut_n9387 (.I0(x264), .I1(x265), .I2(x266), .O(n9387));
  LUT5 #(.INIT(32'h96696996)) lut_n9388 (.I0(x255), .I1(x256), .I2(x257), .I3(n9384), .I4(n9385), .O(n9388));
  LUT5 #(.INIT(32'hFF969600)) lut_n9389 (.I0(x261), .I1(x262), .I2(x263), .I3(n9387), .I4(n9388), .O(n9389));
  LUT3 #(.INIT(8'h96)) lut_n9390 (.I0(n9378), .I1(n9381), .I2(n9382), .O(n9390));
  LUT3 #(.INIT(8'hE8)) lut_n9391 (.I0(n9386), .I1(n9389), .I2(n9390), .O(n9391));
  LUT3 #(.INIT(8'h96)) lut_n9392 (.I0(n9365), .I1(n9373), .I2(n9374), .O(n9392));
  LUT3 #(.INIT(8'hE8)) lut_n9393 (.I0(n9383), .I1(n9391), .I2(n9392), .O(n9393));
  LUT3 #(.INIT(8'h96)) lut_n9394 (.I0(n9335), .I1(n9353), .I2(n9354), .O(n9394));
  LUT3 #(.INIT(8'hE8)) lut_n9395 (.I0(n9375), .I1(n9393), .I2(n9394), .O(n9395));
  LUT3 #(.INIT(8'h96)) lut_n9396 (.I0(x270), .I1(x271), .I2(x272), .O(n9396));
  LUT5 #(.INIT(32'h96696996)) lut_n9397 (.I0(x261), .I1(x262), .I2(x263), .I3(n9387), .I4(n9388), .O(n9397));
  LUT5 #(.INIT(32'hFF969600)) lut_n9398 (.I0(x267), .I1(x268), .I2(x269), .I3(n9396), .I4(n9397), .O(n9398));
  LUT3 #(.INIT(8'h96)) lut_n9399 (.I0(x276), .I1(x277), .I2(x278), .O(n9399));
  LUT5 #(.INIT(32'h96696996)) lut_n9400 (.I0(x267), .I1(x268), .I2(x269), .I3(n9396), .I4(n9397), .O(n9400));
  LUT5 #(.INIT(32'hFF969600)) lut_n9401 (.I0(x273), .I1(x274), .I2(x275), .I3(n9399), .I4(n9400), .O(n9401));
  LUT3 #(.INIT(8'h96)) lut_n9402 (.I0(n9386), .I1(n9389), .I2(n9390), .O(n9402));
  LUT3 #(.INIT(8'hE8)) lut_n9403 (.I0(n9398), .I1(n9401), .I2(n9402), .O(n9403));
  LUT3 #(.INIT(8'h96)) lut_n9404 (.I0(x282), .I1(x283), .I2(x284), .O(n9404));
  LUT5 #(.INIT(32'h96696996)) lut_n9405 (.I0(x273), .I1(x274), .I2(x275), .I3(n9399), .I4(n9400), .O(n9405));
  LUT5 #(.INIT(32'hFF969600)) lut_n9406 (.I0(x279), .I1(x280), .I2(x281), .I3(n9404), .I4(n9405), .O(n9406));
  LUT3 #(.INIT(8'h96)) lut_n9407 (.I0(x288), .I1(x289), .I2(x290), .O(n9407));
  LUT5 #(.INIT(32'h96696996)) lut_n9408 (.I0(x279), .I1(x280), .I2(x281), .I3(n9404), .I4(n9405), .O(n9408));
  LUT5 #(.INIT(32'hFF969600)) lut_n9409 (.I0(x285), .I1(x286), .I2(x287), .I3(n9407), .I4(n9408), .O(n9409));
  LUT3 #(.INIT(8'h96)) lut_n9410 (.I0(n9398), .I1(n9401), .I2(n9402), .O(n9410));
  LUT3 #(.INIT(8'hE8)) lut_n9411 (.I0(n9406), .I1(n9409), .I2(n9410), .O(n9411));
  LUT3 #(.INIT(8'h96)) lut_n9412 (.I0(n9383), .I1(n9391), .I2(n9392), .O(n9412));
  LUT3 #(.INIT(8'hE8)) lut_n9413 (.I0(n9403), .I1(n9411), .I2(n9412), .O(n9413));
  LUT3 #(.INIT(8'h96)) lut_n9414 (.I0(x294), .I1(x295), .I2(x296), .O(n9414));
  LUT5 #(.INIT(32'h96696996)) lut_n9415 (.I0(x285), .I1(x286), .I2(x287), .I3(n9407), .I4(n9408), .O(n9415));
  LUT5 #(.INIT(32'hFF969600)) lut_n9416 (.I0(x291), .I1(x292), .I2(x293), .I3(n9414), .I4(n9415), .O(n9416));
  LUT3 #(.INIT(8'h96)) lut_n9417 (.I0(x297), .I1(x298), .I2(x299), .O(n9417));
  LUT5 #(.INIT(32'h96696996)) lut_n9418 (.I0(x291), .I1(x292), .I2(x293), .I3(n9414), .I4(n9415), .O(n9418));
  LUT5 #(.INIT(32'hFF969600)) lut_n9419 (.I0(x300), .I1(x301), .I2(x302), .I3(n9417), .I4(n9418), .O(n9419));
  LUT3 #(.INIT(8'h96)) lut_n9420 (.I0(n9406), .I1(n9409), .I2(n9410), .O(n9420));
  LUT3 #(.INIT(8'hE8)) lut_n9421 (.I0(n9416), .I1(n9419), .I2(n9420), .O(n9421));
  LUT3 #(.INIT(8'h96)) lut_n9422 (.I0(x306), .I1(x307), .I2(x308), .O(n9422));
  LUT5 #(.INIT(32'h96696996)) lut_n9423 (.I0(x300), .I1(x301), .I2(x302), .I3(n9417), .I4(n9418), .O(n9423));
  LUT5 #(.INIT(32'hFF969600)) lut_n9424 (.I0(x303), .I1(x304), .I2(x305), .I3(n9422), .I4(n9423), .O(n9424));
  LUT3 #(.INIT(8'h96)) lut_n9425 (.I0(x312), .I1(x313), .I2(x314), .O(n9425));
  LUT5 #(.INIT(32'h96696996)) lut_n9426 (.I0(x303), .I1(x304), .I2(x305), .I3(n9422), .I4(n9423), .O(n9426));
  LUT5 #(.INIT(32'hFF969600)) lut_n9427 (.I0(x309), .I1(x310), .I2(x311), .I3(n9425), .I4(n9426), .O(n9427));
  LUT3 #(.INIT(8'h96)) lut_n9428 (.I0(n9416), .I1(n9419), .I2(n9420), .O(n9428));
  LUT3 #(.INIT(8'hE8)) lut_n9429 (.I0(n9424), .I1(n9427), .I2(n9428), .O(n9429));
  LUT3 #(.INIT(8'h96)) lut_n9430 (.I0(n9403), .I1(n9411), .I2(n9412), .O(n9430));
  LUT3 #(.INIT(8'hE8)) lut_n9431 (.I0(n9421), .I1(n9429), .I2(n9430), .O(n9431));
  LUT3 #(.INIT(8'h96)) lut_n9432 (.I0(n9375), .I1(n9393), .I2(n9394), .O(n9432));
  LUT3 #(.INIT(8'hE8)) lut_n9433 (.I0(n9413), .I1(n9431), .I2(n9432), .O(n9433));
  LUT3 #(.INIT(8'h96)) lut_n9434 (.I0(n9317), .I1(n9355), .I2(n9356), .O(n9434));
  LUT3 #(.INIT(8'hE8)) lut_n9435 (.I0(n9395), .I1(n9433), .I2(n9434), .O(n9435));
  LUT3 #(.INIT(8'h96)) lut_n9436 (.I0(n9199), .I1(n9277), .I2(n9278), .O(n9436));
  LUT3 #(.INIT(8'hE8)) lut_n9437 (.I0(n9357), .I1(n9435), .I2(n9436), .O(n9437));
  LUT3 #(.INIT(8'h96)) lut_n9438 (.I0(n9069), .I1(n9147), .I2(n9148), .O(n9438));
  LUT3 #(.INIT(8'hE8)) lut_n9439 (.I0(n9279), .I1(n9437), .I2(n9438), .O(n9439));
  LUT3 #(.INIT(8'h96)) lut_n9440 (.I0(x318), .I1(x319), .I2(x320), .O(n9440));
  LUT5 #(.INIT(32'h96696996)) lut_n9441 (.I0(x309), .I1(x310), .I2(x311), .I3(n9425), .I4(n9426), .O(n9441));
  LUT5 #(.INIT(32'hFF969600)) lut_n9442 (.I0(x315), .I1(x316), .I2(x317), .I3(n9440), .I4(n9441), .O(n9442));
  LUT3 #(.INIT(8'h96)) lut_n9443 (.I0(x324), .I1(x325), .I2(x326), .O(n9443));
  LUT5 #(.INIT(32'h96696996)) lut_n9444 (.I0(x315), .I1(x316), .I2(x317), .I3(n9440), .I4(n9441), .O(n9444));
  LUT5 #(.INIT(32'hFF969600)) lut_n9445 (.I0(x321), .I1(x322), .I2(x323), .I3(n9443), .I4(n9444), .O(n9445));
  LUT3 #(.INIT(8'h96)) lut_n9446 (.I0(n9424), .I1(n9427), .I2(n9428), .O(n9446));
  LUT3 #(.INIT(8'hE8)) lut_n9447 (.I0(n9442), .I1(n9445), .I2(n9446), .O(n9447));
  LUT3 #(.INIT(8'h96)) lut_n9448 (.I0(x330), .I1(x331), .I2(x332), .O(n9448));
  LUT5 #(.INIT(32'h96696996)) lut_n9449 (.I0(x321), .I1(x322), .I2(x323), .I3(n9443), .I4(n9444), .O(n9449));
  LUT5 #(.INIT(32'hFF969600)) lut_n9450 (.I0(x327), .I1(x328), .I2(x329), .I3(n9448), .I4(n9449), .O(n9450));
  LUT3 #(.INIT(8'h96)) lut_n9451 (.I0(x336), .I1(x337), .I2(x338), .O(n9451));
  LUT5 #(.INIT(32'h96696996)) lut_n9452 (.I0(x327), .I1(x328), .I2(x329), .I3(n9448), .I4(n9449), .O(n9452));
  LUT5 #(.INIT(32'hFF969600)) lut_n9453 (.I0(x333), .I1(x334), .I2(x335), .I3(n9451), .I4(n9452), .O(n9453));
  LUT3 #(.INIT(8'h96)) lut_n9454 (.I0(n9442), .I1(n9445), .I2(n9446), .O(n9454));
  LUT3 #(.INIT(8'hE8)) lut_n9455 (.I0(n9450), .I1(n9453), .I2(n9454), .O(n9455));
  LUT3 #(.INIT(8'h96)) lut_n9456 (.I0(n9421), .I1(n9429), .I2(n9430), .O(n9456));
  LUT3 #(.INIT(8'hE8)) lut_n9457 (.I0(n9447), .I1(n9455), .I2(n9456), .O(n9457));
  LUT3 #(.INIT(8'h96)) lut_n9458 (.I0(x342), .I1(x343), .I2(x344), .O(n9458));
  LUT5 #(.INIT(32'h96696996)) lut_n9459 (.I0(x333), .I1(x334), .I2(x335), .I3(n9451), .I4(n9452), .O(n9459));
  LUT5 #(.INIT(32'hFF969600)) lut_n9460 (.I0(x339), .I1(x340), .I2(x341), .I3(n9458), .I4(n9459), .O(n9460));
  LUT3 #(.INIT(8'h96)) lut_n9461 (.I0(x348), .I1(x349), .I2(x350), .O(n9461));
  LUT5 #(.INIT(32'h96696996)) lut_n9462 (.I0(x339), .I1(x340), .I2(x341), .I3(n9458), .I4(n9459), .O(n9462));
  LUT5 #(.INIT(32'hFF969600)) lut_n9463 (.I0(x345), .I1(x346), .I2(x347), .I3(n9461), .I4(n9462), .O(n9463));
  LUT3 #(.INIT(8'h96)) lut_n9464 (.I0(n9450), .I1(n9453), .I2(n9454), .O(n9464));
  LUT3 #(.INIT(8'hE8)) lut_n9465 (.I0(n9460), .I1(n9463), .I2(n9464), .O(n9465));
  LUT3 #(.INIT(8'h96)) lut_n9466 (.I0(x354), .I1(x355), .I2(x356), .O(n9466));
  LUT5 #(.INIT(32'h96696996)) lut_n9467 (.I0(x345), .I1(x346), .I2(x347), .I3(n9461), .I4(n9462), .O(n9467));
  LUT5 #(.INIT(32'hFF969600)) lut_n9468 (.I0(x351), .I1(x352), .I2(x353), .I3(n9466), .I4(n9467), .O(n9468));
  LUT3 #(.INIT(8'h96)) lut_n9469 (.I0(x360), .I1(x361), .I2(x362), .O(n9469));
  LUT5 #(.INIT(32'h96696996)) lut_n9470 (.I0(x351), .I1(x352), .I2(x353), .I3(n9466), .I4(n9467), .O(n9470));
  LUT5 #(.INIT(32'hFF969600)) lut_n9471 (.I0(x357), .I1(x358), .I2(x359), .I3(n9469), .I4(n9470), .O(n9471));
  LUT3 #(.INIT(8'h96)) lut_n9472 (.I0(n9460), .I1(n9463), .I2(n9464), .O(n9472));
  LUT3 #(.INIT(8'hE8)) lut_n9473 (.I0(n9468), .I1(n9471), .I2(n9472), .O(n9473));
  LUT3 #(.INIT(8'h96)) lut_n9474 (.I0(n9447), .I1(n9455), .I2(n9456), .O(n9474));
  LUT3 #(.INIT(8'hE8)) lut_n9475 (.I0(n9465), .I1(n9473), .I2(n9474), .O(n9475));
  LUT3 #(.INIT(8'h96)) lut_n9476 (.I0(n9413), .I1(n9431), .I2(n9432), .O(n9476));
  LUT3 #(.INIT(8'hE8)) lut_n9477 (.I0(n9457), .I1(n9475), .I2(n9476), .O(n9477));
  LUT3 #(.INIT(8'h96)) lut_n9478 (.I0(x366), .I1(x367), .I2(x368), .O(n9478));
  LUT5 #(.INIT(32'h96696996)) lut_n9479 (.I0(x357), .I1(x358), .I2(x359), .I3(n9469), .I4(n9470), .O(n9479));
  LUT5 #(.INIT(32'hFF969600)) lut_n9480 (.I0(x363), .I1(x364), .I2(x365), .I3(n9478), .I4(n9479), .O(n9480));
  LUT3 #(.INIT(8'h96)) lut_n9481 (.I0(x372), .I1(x373), .I2(x374), .O(n9481));
  LUT5 #(.INIT(32'h96696996)) lut_n9482 (.I0(x363), .I1(x364), .I2(x365), .I3(n9478), .I4(n9479), .O(n9482));
  LUT5 #(.INIT(32'hFF969600)) lut_n9483 (.I0(x369), .I1(x370), .I2(x371), .I3(n9481), .I4(n9482), .O(n9483));
  LUT3 #(.INIT(8'h96)) lut_n9484 (.I0(n9468), .I1(n9471), .I2(n9472), .O(n9484));
  LUT3 #(.INIT(8'hE8)) lut_n9485 (.I0(n9480), .I1(n9483), .I2(n9484), .O(n9485));
  LUT3 #(.INIT(8'h96)) lut_n9486 (.I0(x378), .I1(x379), .I2(x380), .O(n9486));
  LUT5 #(.INIT(32'h96696996)) lut_n9487 (.I0(x369), .I1(x370), .I2(x371), .I3(n9481), .I4(n9482), .O(n9487));
  LUT5 #(.INIT(32'hFF969600)) lut_n9488 (.I0(x375), .I1(x376), .I2(x377), .I3(n9486), .I4(n9487), .O(n9488));
  LUT3 #(.INIT(8'h96)) lut_n9489 (.I0(x384), .I1(x385), .I2(x386), .O(n9489));
  LUT5 #(.INIT(32'h96696996)) lut_n9490 (.I0(x375), .I1(x376), .I2(x377), .I3(n9486), .I4(n9487), .O(n9490));
  LUT5 #(.INIT(32'hFF969600)) lut_n9491 (.I0(x381), .I1(x382), .I2(x383), .I3(n9489), .I4(n9490), .O(n9491));
  LUT3 #(.INIT(8'h96)) lut_n9492 (.I0(n9480), .I1(n9483), .I2(n9484), .O(n9492));
  LUT3 #(.INIT(8'hE8)) lut_n9493 (.I0(n9488), .I1(n9491), .I2(n9492), .O(n9493));
  LUT3 #(.INIT(8'h96)) lut_n9494 (.I0(n9465), .I1(n9473), .I2(n9474), .O(n9494));
  LUT3 #(.INIT(8'hE8)) lut_n9495 (.I0(n9485), .I1(n9493), .I2(n9494), .O(n9495));
  LUT3 #(.INIT(8'h96)) lut_n9496 (.I0(x390), .I1(x391), .I2(x392), .O(n9496));
  LUT5 #(.INIT(32'h96696996)) lut_n9497 (.I0(x381), .I1(x382), .I2(x383), .I3(n9489), .I4(n9490), .O(n9497));
  LUT5 #(.INIT(32'hFF969600)) lut_n9498 (.I0(x387), .I1(x388), .I2(x389), .I3(n9496), .I4(n9497), .O(n9498));
  LUT3 #(.INIT(8'h96)) lut_n9499 (.I0(x396), .I1(x397), .I2(x398), .O(n9499));
  LUT5 #(.INIT(32'h96696996)) lut_n9500 (.I0(x387), .I1(x388), .I2(x389), .I3(n9496), .I4(n9497), .O(n9500));
  LUT5 #(.INIT(32'hFF969600)) lut_n9501 (.I0(x393), .I1(x394), .I2(x395), .I3(n9499), .I4(n9500), .O(n9501));
  LUT3 #(.INIT(8'h96)) lut_n9502 (.I0(n9488), .I1(n9491), .I2(n9492), .O(n9502));
  LUT3 #(.INIT(8'hE8)) lut_n9503 (.I0(n9498), .I1(n9501), .I2(n9502), .O(n9503));
  LUT3 #(.INIT(8'h96)) lut_n9504 (.I0(x402), .I1(x403), .I2(x404), .O(n9504));
  LUT5 #(.INIT(32'h96696996)) lut_n9505 (.I0(x393), .I1(x394), .I2(x395), .I3(n9499), .I4(n9500), .O(n9505));
  LUT5 #(.INIT(32'hFF969600)) lut_n9506 (.I0(x399), .I1(x400), .I2(x401), .I3(n9504), .I4(n9505), .O(n9506));
  LUT3 #(.INIT(8'h96)) lut_n9507 (.I0(x408), .I1(x409), .I2(x410), .O(n9507));
  LUT5 #(.INIT(32'h96696996)) lut_n9508 (.I0(x399), .I1(x400), .I2(x401), .I3(n9504), .I4(n9505), .O(n9508));
  LUT5 #(.INIT(32'hFF969600)) lut_n9509 (.I0(x405), .I1(x406), .I2(x407), .I3(n9507), .I4(n9508), .O(n9509));
  LUT3 #(.INIT(8'h96)) lut_n9510 (.I0(n9498), .I1(n9501), .I2(n9502), .O(n9510));
  LUT3 #(.INIT(8'hE8)) lut_n9511 (.I0(n9506), .I1(n9509), .I2(n9510), .O(n9511));
  LUT3 #(.INIT(8'h96)) lut_n9512 (.I0(n9485), .I1(n9493), .I2(n9494), .O(n9512));
  LUT3 #(.INIT(8'hE8)) lut_n9513 (.I0(n9503), .I1(n9511), .I2(n9512), .O(n9513));
  LUT3 #(.INIT(8'h96)) lut_n9514 (.I0(n9457), .I1(n9475), .I2(n9476), .O(n9514));
  LUT3 #(.INIT(8'hE8)) lut_n9515 (.I0(n9495), .I1(n9513), .I2(n9514), .O(n9515));
  LUT3 #(.INIT(8'h96)) lut_n9516 (.I0(n9395), .I1(n9433), .I2(n9434), .O(n9516));
  LUT3 #(.INIT(8'hE8)) lut_n9517 (.I0(n9477), .I1(n9515), .I2(n9516), .O(n9517));
  LUT3 #(.INIT(8'h96)) lut_n9518 (.I0(x414), .I1(x415), .I2(x416), .O(n9518));
  LUT5 #(.INIT(32'h96696996)) lut_n9519 (.I0(x405), .I1(x406), .I2(x407), .I3(n9507), .I4(n9508), .O(n9519));
  LUT5 #(.INIT(32'hFF969600)) lut_n9520 (.I0(x411), .I1(x412), .I2(x413), .I3(n9518), .I4(n9519), .O(n9520));
  LUT3 #(.INIT(8'h96)) lut_n9521 (.I0(x420), .I1(x421), .I2(x422), .O(n9521));
  LUT5 #(.INIT(32'h96696996)) lut_n9522 (.I0(x411), .I1(x412), .I2(x413), .I3(n9518), .I4(n9519), .O(n9522));
  LUT5 #(.INIT(32'hFF969600)) lut_n9523 (.I0(x417), .I1(x418), .I2(x419), .I3(n9521), .I4(n9522), .O(n9523));
  LUT3 #(.INIT(8'h96)) lut_n9524 (.I0(n9506), .I1(n9509), .I2(n9510), .O(n9524));
  LUT3 #(.INIT(8'hE8)) lut_n9525 (.I0(n9520), .I1(n9523), .I2(n9524), .O(n9525));
  LUT3 #(.INIT(8'h96)) lut_n9526 (.I0(x426), .I1(x427), .I2(x428), .O(n9526));
  LUT5 #(.INIT(32'h96696996)) lut_n9527 (.I0(x417), .I1(x418), .I2(x419), .I3(n9521), .I4(n9522), .O(n9527));
  LUT5 #(.INIT(32'hFF969600)) lut_n9528 (.I0(x423), .I1(x424), .I2(x425), .I3(n9526), .I4(n9527), .O(n9528));
  LUT3 #(.INIT(8'h96)) lut_n9529 (.I0(x432), .I1(x433), .I2(x434), .O(n9529));
  LUT5 #(.INIT(32'h96696996)) lut_n9530 (.I0(x423), .I1(x424), .I2(x425), .I3(n9526), .I4(n9527), .O(n9530));
  LUT5 #(.INIT(32'hFF969600)) lut_n9531 (.I0(x429), .I1(x430), .I2(x431), .I3(n9529), .I4(n9530), .O(n9531));
  LUT3 #(.INIT(8'h96)) lut_n9532 (.I0(n9520), .I1(n9523), .I2(n9524), .O(n9532));
  LUT3 #(.INIT(8'hE8)) lut_n9533 (.I0(n9528), .I1(n9531), .I2(n9532), .O(n9533));
  LUT3 #(.INIT(8'h96)) lut_n9534 (.I0(n9503), .I1(n9511), .I2(n9512), .O(n9534));
  LUT3 #(.INIT(8'hE8)) lut_n9535 (.I0(n9525), .I1(n9533), .I2(n9534), .O(n9535));
  LUT3 #(.INIT(8'h96)) lut_n9536 (.I0(x438), .I1(x439), .I2(x440), .O(n9536));
  LUT5 #(.INIT(32'h96696996)) lut_n9537 (.I0(x429), .I1(x430), .I2(x431), .I3(n9529), .I4(n9530), .O(n9537));
  LUT5 #(.INIT(32'hFF969600)) lut_n9538 (.I0(x435), .I1(x436), .I2(x437), .I3(n9536), .I4(n9537), .O(n9538));
  LUT3 #(.INIT(8'h96)) lut_n9539 (.I0(x444), .I1(x445), .I2(x446), .O(n9539));
  LUT5 #(.INIT(32'h96696996)) lut_n9540 (.I0(x435), .I1(x436), .I2(x437), .I3(n9536), .I4(n9537), .O(n9540));
  LUT5 #(.INIT(32'hFF969600)) lut_n9541 (.I0(x441), .I1(x442), .I2(x443), .I3(n9539), .I4(n9540), .O(n9541));
  LUT3 #(.INIT(8'h96)) lut_n9542 (.I0(n9528), .I1(n9531), .I2(n9532), .O(n9542));
  LUT3 #(.INIT(8'hE8)) lut_n9543 (.I0(n9538), .I1(n9541), .I2(n9542), .O(n9543));
  LUT3 #(.INIT(8'h96)) lut_n9544 (.I0(x450), .I1(x451), .I2(x452), .O(n9544));
  LUT5 #(.INIT(32'h96696996)) lut_n9545 (.I0(x441), .I1(x442), .I2(x443), .I3(n9539), .I4(n9540), .O(n9545));
  LUT5 #(.INIT(32'hFF969600)) lut_n9546 (.I0(x447), .I1(x448), .I2(x449), .I3(n9544), .I4(n9545), .O(n9546));
  LUT3 #(.INIT(8'h96)) lut_n9547 (.I0(x456), .I1(x457), .I2(x458), .O(n9547));
  LUT5 #(.INIT(32'h96696996)) lut_n9548 (.I0(x447), .I1(x448), .I2(x449), .I3(n9544), .I4(n9545), .O(n9548));
  LUT5 #(.INIT(32'hFF969600)) lut_n9549 (.I0(x453), .I1(x454), .I2(x455), .I3(n9547), .I4(n9548), .O(n9549));
  LUT3 #(.INIT(8'h96)) lut_n9550 (.I0(n9538), .I1(n9541), .I2(n9542), .O(n9550));
  LUT3 #(.INIT(8'hE8)) lut_n9551 (.I0(n9546), .I1(n9549), .I2(n9550), .O(n9551));
  LUT3 #(.INIT(8'h96)) lut_n9552 (.I0(n9525), .I1(n9533), .I2(n9534), .O(n9552));
  LUT3 #(.INIT(8'hE8)) lut_n9553 (.I0(n9543), .I1(n9551), .I2(n9552), .O(n9553));
  LUT3 #(.INIT(8'h96)) lut_n9554 (.I0(n9495), .I1(n9513), .I2(n9514), .O(n9554));
  LUT3 #(.INIT(8'hE8)) lut_n9555 (.I0(n9535), .I1(n9553), .I2(n9554), .O(n9555));
  LUT3 #(.INIT(8'h96)) lut_n9556 (.I0(x462), .I1(x463), .I2(x464), .O(n9556));
  LUT5 #(.INIT(32'h96696996)) lut_n9557 (.I0(x453), .I1(x454), .I2(x455), .I3(n9547), .I4(n9548), .O(n9557));
  LUT5 #(.INIT(32'hFF969600)) lut_n9558 (.I0(x459), .I1(x460), .I2(x461), .I3(n9556), .I4(n9557), .O(n9558));
  LUT3 #(.INIT(8'h96)) lut_n9559 (.I0(x468), .I1(x469), .I2(x470), .O(n9559));
  LUT5 #(.INIT(32'h96696996)) lut_n9560 (.I0(x459), .I1(x460), .I2(x461), .I3(n9556), .I4(n9557), .O(n9560));
  LUT5 #(.INIT(32'hFF969600)) lut_n9561 (.I0(x465), .I1(x466), .I2(x467), .I3(n9559), .I4(n9560), .O(n9561));
  LUT3 #(.INIT(8'h96)) lut_n9562 (.I0(n9546), .I1(n9549), .I2(n9550), .O(n9562));
  LUT3 #(.INIT(8'hE8)) lut_n9563 (.I0(n9558), .I1(n9561), .I2(n9562), .O(n9563));
  LUT3 #(.INIT(8'h96)) lut_n9564 (.I0(x474), .I1(x475), .I2(x476), .O(n9564));
  LUT5 #(.INIT(32'h96696996)) lut_n9565 (.I0(x465), .I1(x466), .I2(x467), .I3(n9559), .I4(n9560), .O(n9565));
  LUT5 #(.INIT(32'hFF969600)) lut_n9566 (.I0(x471), .I1(x472), .I2(x473), .I3(n9564), .I4(n9565), .O(n9566));
  LUT3 #(.INIT(8'h96)) lut_n9567 (.I0(x480), .I1(x481), .I2(x482), .O(n9567));
  LUT5 #(.INIT(32'h96696996)) lut_n9568 (.I0(x471), .I1(x472), .I2(x473), .I3(n9564), .I4(n9565), .O(n9568));
  LUT5 #(.INIT(32'hFF969600)) lut_n9569 (.I0(x477), .I1(x478), .I2(x479), .I3(n9567), .I4(n9568), .O(n9569));
  LUT3 #(.INIT(8'h96)) lut_n9570 (.I0(n9558), .I1(n9561), .I2(n9562), .O(n9570));
  LUT3 #(.INIT(8'hE8)) lut_n9571 (.I0(n9566), .I1(n9569), .I2(n9570), .O(n9571));
  LUT3 #(.INIT(8'h96)) lut_n9572 (.I0(n9543), .I1(n9551), .I2(n9552), .O(n9572));
  LUT3 #(.INIT(8'hE8)) lut_n9573 (.I0(n9563), .I1(n9571), .I2(n9572), .O(n9573));
  LUT3 #(.INIT(8'h96)) lut_n9574 (.I0(x486), .I1(x487), .I2(x488), .O(n9574));
  LUT5 #(.INIT(32'h96696996)) lut_n9575 (.I0(x477), .I1(x478), .I2(x479), .I3(n9567), .I4(n9568), .O(n9575));
  LUT5 #(.INIT(32'hFF969600)) lut_n9576 (.I0(x483), .I1(x484), .I2(x485), .I3(n9574), .I4(n9575), .O(n9576));
  LUT3 #(.INIT(8'h96)) lut_n9577 (.I0(x492), .I1(x493), .I2(x494), .O(n9577));
  LUT5 #(.INIT(32'h96696996)) lut_n9578 (.I0(x483), .I1(x484), .I2(x485), .I3(n9574), .I4(n9575), .O(n9578));
  LUT5 #(.INIT(32'hFF969600)) lut_n9579 (.I0(x489), .I1(x490), .I2(x491), .I3(n9577), .I4(n9578), .O(n9579));
  LUT3 #(.INIT(8'h96)) lut_n9580 (.I0(n9566), .I1(n9569), .I2(n9570), .O(n9580));
  LUT3 #(.INIT(8'hE8)) lut_n9581 (.I0(n9576), .I1(n9579), .I2(n9580), .O(n9581));
  LUT3 #(.INIT(8'h96)) lut_n9582 (.I0(x498), .I1(x499), .I2(x500), .O(n9582));
  LUT5 #(.INIT(32'h96696996)) lut_n9583 (.I0(x489), .I1(x490), .I2(x491), .I3(n9577), .I4(n9578), .O(n9583));
  LUT5 #(.INIT(32'hFF969600)) lut_n9584 (.I0(x495), .I1(x496), .I2(x497), .I3(n9582), .I4(n9583), .O(n9584));
  LUT3 #(.INIT(8'h96)) lut_n9585 (.I0(x504), .I1(x505), .I2(x506), .O(n9585));
  LUT5 #(.INIT(32'h96696996)) lut_n9586 (.I0(x495), .I1(x496), .I2(x497), .I3(n9582), .I4(n9583), .O(n9586));
  LUT5 #(.INIT(32'hFF969600)) lut_n9587 (.I0(x501), .I1(x502), .I2(x503), .I3(n9585), .I4(n9586), .O(n9587));
  LUT3 #(.INIT(8'h96)) lut_n9588 (.I0(n9576), .I1(n9579), .I2(n9580), .O(n9588));
  LUT3 #(.INIT(8'hE8)) lut_n9589 (.I0(n9584), .I1(n9587), .I2(n9588), .O(n9589));
  LUT3 #(.INIT(8'h96)) lut_n9590 (.I0(n9563), .I1(n9571), .I2(n9572), .O(n9590));
  LUT3 #(.INIT(8'hE8)) lut_n9591 (.I0(n9581), .I1(n9589), .I2(n9590), .O(n9591));
  LUT3 #(.INIT(8'h96)) lut_n9592 (.I0(n9535), .I1(n9553), .I2(n9554), .O(n9592));
  LUT3 #(.INIT(8'hE8)) lut_n9593 (.I0(n9573), .I1(n9591), .I2(n9592), .O(n9593));
  LUT3 #(.INIT(8'h96)) lut_n9594 (.I0(n9477), .I1(n9515), .I2(n9516), .O(n9594));
  LUT3 #(.INIT(8'hE8)) lut_n9595 (.I0(n9555), .I1(n9593), .I2(n9594), .O(n9595));
  LUT3 #(.INIT(8'h96)) lut_n9596 (.I0(n9357), .I1(n9435), .I2(n9436), .O(n9596));
  LUT3 #(.INIT(8'hE8)) lut_n9597 (.I0(n9517), .I1(n9595), .I2(n9596), .O(n9597));
  LUT3 #(.INIT(8'h96)) lut_n9598 (.I0(x510), .I1(x511), .I2(x512), .O(n9598));
  LUT5 #(.INIT(32'h96696996)) lut_n9599 (.I0(x501), .I1(x502), .I2(x503), .I3(n9585), .I4(n9586), .O(n9599));
  LUT5 #(.INIT(32'hFF969600)) lut_n9600 (.I0(x507), .I1(x508), .I2(x509), .I3(n9598), .I4(n9599), .O(n9600));
  LUT3 #(.INIT(8'h96)) lut_n9601 (.I0(x516), .I1(x517), .I2(x518), .O(n9601));
  LUT5 #(.INIT(32'h96696996)) lut_n9602 (.I0(x507), .I1(x508), .I2(x509), .I3(n9598), .I4(n9599), .O(n9602));
  LUT5 #(.INIT(32'hFF969600)) lut_n9603 (.I0(x513), .I1(x514), .I2(x515), .I3(n9601), .I4(n9602), .O(n9603));
  LUT3 #(.INIT(8'h96)) lut_n9604 (.I0(n9584), .I1(n9587), .I2(n9588), .O(n9604));
  LUT3 #(.INIT(8'hE8)) lut_n9605 (.I0(n9600), .I1(n9603), .I2(n9604), .O(n9605));
  LUT3 #(.INIT(8'h96)) lut_n9606 (.I0(x522), .I1(x523), .I2(x524), .O(n9606));
  LUT5 #(.INIT(32'h96696996)) lut_n9607 (.I0(x513), .I1(x514), .I2(x515), .I3(n9601), .I4(n9602), .O(n9607));
  LUT5 #(.INIT(32'hFF969600)) lut_n9608 (.I0(x519), .I1(x520), .I2(x521), .I3(n9606), .I4(n9607), .O(n9608));
  LUT3 #(.INIT(8'h96)) lut_n9609 (.I0(x528), .I1(x529), .I2(x530), .O(n9609));
  LUT5 #(.INIT(32'h96696996)) lut_n9610 (.I0(x519), .I1(x520), .I2(x521), .I3(n9606), .I4(n9607), .O(n9610));
  LUT5 #(.INIT(32'hFF969600)) lut_n9611 (.I0(x525), .I1(x526), .I2(x527), .I3(n9609), .I4(n9610), .O(n9611));
  LUT3 #(.INIT(8'h96)) lut_n9612 (.I0(n9600), .I1(n9603), .I2(n9604), .O(n9612));
  LUT3 #(.INIT(8'hE8)) lut_n9613 (.I0(n9608), .I1(n9611), .I2(n9612), .O(n9613));
  LUT3 #(.INIT(8'h96)) lut_n9614 (.I0(n9581), .I1(n9589), .I2(n9590), .O(n9614));
  LUT3 #(.INIT(8'hE8)) lut_n9615 (.I0(n9605), .I1(n9613), .I2(n9614), .O(n9615));
  LUT3 #(.INIT(8'h96)) lut_n9616 (.I0(x534), .I1(x535), .I2(x536), .O(n9616));
  LUT5 #(.INIT(32'h96696996)) lut_n9617 (.I0(x525), .I1(x526), .I2(x527), .I3(n9609), .I4(n9610), .O(n9617));
  LUT5 #(.INIT(32'hFF969600)) lut_n9618 (.I0(x531), .I1(x532), .I2(x533), .I3(n9616), .I4(n9617), .O(n9618));
  LUT3 #(.INIT(8'h96)) lut_n9619 (.I0(x540), .I1(x541), .I2(x542), .O(n9619));
  LUT5 #(.INIT(32'h96696996)) lut_n9620 (.I0(x531), .I1(x532), .I2(x533), .I3(n9616), .I4(n9617), .O(n9620));
  LUT5 #(.INIT(32'hFF969600)) lut_n9621 (.I0(x537), .I1(x538), .I2(x539), .I3(n9619), .I4(n9620), .O(n9621));
  LUT3 #(.INIT(8'h96)) lut_n9622 (.I0(n9608), .I1(n9611), .I2(n9612), .O(n9622));
  LUT3 #(.INIT(8'hE8)) lut_n9623 (.I0(n9618), .I1(n9621), .I2(n9622), .O(n9623));
  LUT3 #(.INIT(8'h96)) lut_n9624 (.I0(x546), .I1(x547), .I2(x548), .O(n9624));
  LUT5 #(.INIT(32'h96696996)) lut_n9625 (.I0(x537), .I1(x538), .I2(x539), .I3(n9619), .I4(n9620), .O(n9625));
  LUT5 #(.INIT(32'hFF969600)) lut_n9626 (.I0(x543), .I1(x544), .I2(x545), .I3(n9624), .I4(n9625), .O(n9626));
  LUT3 #(.INIT(8'h96)) lut_n9627 (.I0(x552), .I1(x553), .I2(x554), .O(n9627));
  LUT5 #(.INIT(32'h96696996)) lut_n9628 (.I0(x543), .I1(x544), .I2(x545), .I3(n9624), .I4(n9625), .O(n9628));
  LUT5 #(.INIT(32'hFF969600)) lut_n9629 (.I0(x549), .I1(x550), .I2(x551), .I3(n9627), .I4(n9628), .O(n9629));
  LUT3 #(.INIT(8'h96)) lut_n9630 (.I0(n9618), .I1(n9621), .I2(n9622), .O(n9630));
  LUT3 #(.INIT(8'hE8)) lut_n9631 (.I0(n9626), .I1(n9629), .I2(n9630), .O(n9631));
  LUT3 #(.INIT(8'h96)) lut_n9632 (.I0(n9605), .I1(n9613), .I2(n9614), .O(n9632));
  LUT3 #(.INIT(8'hE8)) lut_n9633 (.I0(n9623), .I1(n9631), .I2(n9632), .O(n9633));
  LUT3 #(.INIT(8'h96)) lut_n9634 (.I0(n9573), .I1(n9591), .I2(n9592), .O(n9634));
  LUT3 #(.INIT(8'hE8)) lut_n9635 (.I0(n9615), .I1(n9633), .I2(n9634), .O(n9635));
  LUT3 #(.INIT(8'h96)) lut_n9636 (.I0(x558), .I1(x559), .I2(x560), .O(n9636));
  LUT5 #(.INIT(32'h96696996)) lut_n9637 (.I0(x549), .I1(x550), .I2(x551), .I3(n9627), .I4(n9628), .O(n9637));
  LUT5 #(.INIT(32'hFF969600)) lut_n9638 (.I0(x555), .I1(x556), .I2(x557), .I3(n9636), .I4(n9637), .O(n9638));
  LUT3 #(.INIT(8'h96)) lut_n9639 (.I0(x564), .I1(x565), .I2(x566), .O(n9639));
  LUT5 #(.INIT(32'h96696996)) lut_n9640 (.I0(x555), .I1(x556), .I2(x557), .I3(n9636), .I4(n9637), .O(n9640));
  LUT5 #(.INIT(32'hFF969600)) lut_n9641 (.I0(x561), .I1(x562), .I2(x563), .I3(n9639), .I4(n9640), .O(n9641));
  LUT3 #(.INIT(8'h96)) lut_n9642 (.I0(n9626), .I1(n9629), .I2(n9630), .O(n9642));
  LUT3 #(.INIT(8'hE8)) lut_n9643 (.I0(n9638), .I1(n9641), .I2(n9642), .O(n9643));
  LUT3 #(.INIT(8'h96)) lut_n9644 (.I0(x570), .I1(x571), .I2(x572), .O(n9644));
  LUT5 #(.INIT(32'h96696996)) lut_n9645 (.I0(x561), .I1(x562), .I2(x563), .I3(n9639), .I4(n9640), .O(n9645));
  LUT5 #(.INIT(32'hFF969600)) lut_n9646 (.I0(x567), .I1(x568), .I2(x569), .I3(n9644), .I4(n9645), .O(n9646));
  LUT3 #(.INIT(8'h96)) lut_n9647 (.I0(x576), .I1(x577), .I2(x578), .O(n9647));
  LUT5 #(.INIT(32'h96696996)) lut_n9648 (.I0(x567), .I1(x568), .I2(x569), .I3(n9644), .I4(n9645), .O(n9648));
  LUT5 #(.INIT(32'hFF969600)) lut_n9649 (.I0(x573), .I1(x574), .I2(x575), .I3(n9647), .I4(n9648), .O(n9649));
  LUT3 #(.INIT(8'h96)) lut_n9650 (.I0(n9638), .I1(n9641), .I2(n9642), .O(n9650));
  LUT3 #(.INIT(8'hE8)) lut_n9651 (.I0(n9646), .I1(n9649), .I2(n9650), .O(n9651));
  LUT3 #(.INIT(8'h96)) lut_n9652 (.I0(n9623), .I1(n9631), .I2(n9632), .O(n9652));
  LUT3 #(.INIT(8'hE8)) lut_n9653 (.I0(n9643), .I1(n9651), .I2(n9652), .O(n9653));
  LUT3 #(.INIT(8'h96)) lut_n9654 (.I0(x582), .I1(x583), .I2(x584), .O(n9654));
  LUT5 #(.INIT(32'h96696996)) lut_n9655 (.I0(x573), .I1(x574), .I2(x575), .I3(n9647), .I4(n9648), .O(n9655));
  LUT5 #(.INIT(32'hFF969600)) lut_n9656 (.I0(x579), .I1(x580), .I2(x581), .I3(n9654), .I4(n9655), .O(n9656));
  LUT3 #(.INIT(8'h96)) lut_n9657 (.I0(x588), .I1(x589), .I2(x590), .O(n9657));
  LUT5 #(.INIT(32'h96696996)) lut_n9658 (.I0(x579), .I1(x580), .I2(x581), .I3(n9654), .I4(n9655), .O(n9658));
  LUT5 #(.INIT(32'hFF969600)) lut_n9659 (.I0(x585), .I1(x586), .I2(x587), .I3(n9657), .I4(n9658), .O(n9659));
  LUT3 #(.INIT(8'h96)) lut_n9660 (.I0(n9646), .I1(n9649), .I2(n9650), .O(n9660));
  LUT3 #(.INIT(8'hE8)) lut_n9661 (.I0(n9656), .I1(n9659), .I2(n9660), .O(n9661));
  LUT3 #(.INIT(8'h96)) lut_n9662 (.I0(x594), .I1(x595), .I2(x596), .O(n9662));
  LUT5 #(.INIT(32'h96696996)) lut_n9663 (.I0(x585), .I1(x586), .I2(x587), .I3(n9657), .I4(n9658), .O(n9663));
  LUT5 #(.INIT(32'hFF969600)) lut_n9664 (.I0(x591), .I1(x592), .I2(x593), .I3(n9662), .I4(n9663), .O(n9664));
  LUT3 #(.INIT(8'h96)) lut_n9665 (.I0(x600), .I1(x601), .I2(x602), .O(n9665));
  LUT5 #(.INIT(32'h96696996)) lut_n9666 (.I0(x591), .I1(x592), .I2(x593), .I3(n9662), .I4(n9663), .O(n9666));
  LUT5 #(.INIT(32'hFF969600)) lut_n9667 (.I0(x597), .I1(x598), .I2(x599), .I3(n9665), .I4(n9666), .O(n9667));
  LUT3 #(.INIT(8'h96)) lut_n9668 (.I0(n9656), .I1(n9659), .I2(n9660), .O(n9668));
  LUT3 #(.INIT(8'hE8)) lut_n9669 (.I0(n9664), .I1(n9667), .I2(n9668), .O(n9669));
  LUT3 #(.INIT(8'h96)) lut_n9670 (.I0(n9643), .I1(n9651), .I2(n9652), .O(n9670));
  LUT3 #(.INIT(8'hE8)) lut_n9671 (.I0(n9661), .I1(n9669), .I2(n9670), .O(n9671));
  LUT3 #(.INIT(8'h96)) lut_n9672 (.I0(n9615), .I1(n9633), .I2(n9634), .O(n9672));
  LUT3 #(.INIT(8'hE8)) lut_n9673 (.I0(n9653), .I1(n9671), .I2(n9672), .O(n9673));
  LUT3 #(.INIT(8'h96)) lut_n9674 (.I0(n9555), .I1(n9593), .I2(n9594), .O(n9674));
  LUT3 #(.INIT(8'hE8)) lut_n9675 (.I0(n9635), .I1(n9673), .I2(n9674), .O(n9675));
  LUT3 #(.INIT(8'h96)) lut_n9676 (.I0(x606), .I1(x607), .I2(x608), .O(n9676));
  LUT5 #(.INIT(32'h96696996)) lut_n9677 (.I0(x597), .I1(x598), .I2(x599), .I3(n9665), .I4(n9666), .O(n9677));
  LUT5 #(.INIT(32'hFF969600)) lut_n9678 (.I0(x603), .I1(x604), .I2(x605), .I3(n9676), .I4(n9677), .O(n9678));
  LUT3 #(.INIT(8'h96)) lut_n9679 (.I0(x612), .I1(x613), .I2(x614), .O(n9679));
  LUT5 #(.INIT(32'h96696996)) lut_n9680 (.I0(x603), .I1(x604), .I2(x605), .I3(n9676), .I4(n9677), .O(n9680));
  LUT5 #(.INIT(32'hFF969600)) lut_n9681 (.I0(x609), .I1(x610), .I2(x611), .I3(n9679), .I4(n9680), .O(n9681));
  LUT3 #(.INIT(8'h96)) lut_n9682 (.I0(n9664), .I1(n9667), .I2(n9668), .O(n9682));
  LUT3 #(.INIT(8'hE8)) lut_n9683 (.I0(n9678), .I1(n9681), .I2(n9682), .O(n9683));
  LUT3 #(.INIT(8'h96)) lut_n9684 (.I0(x618), .I1(x619), .I2(x620), .O(n9684));
  LUT5 #(.INIT(32'h96696996)) lut_n9685 (.I0(x609), .I1(x610), .I2(x611), .I3(n9679), .I4(n9680), .O(n9685));
  LUT5 #(.INIT(32'hFF969600)) lut_n9686 (.I0(x615), .I1(x616), .I2(x617), .I3(n9684), .I4(n9685), .O(n9686));
  LUT3 #(.INIT(8'h96)) lut_n9687 (.I0(x624), .I1(x625), .I2(x626), .O(n9687));
  LUT5 #(.INIT(32'h96696996)) lut_n9688 (.I0(x615), .I1(x616), .I2(x617), .I3(n9684), .I4(n9685), .O(n9688));
  LUT5 #(.INIT(32'hFF969600)) lut_n9689 (.I0(x621), .I1(x622), .I2(x623), .I3(n9687), .I4(n9688), .O(n9689));
  LUT3 #(.INIT(8'h96)) lut_n9690 (.I0(n9678), .I1(n9681), .I2(n9682), .O(n9690));
  LUT3 #(.INIT(8'hE8)) lut_n9691 (.I0(n9686), .I1(n9689), .I2(n9690), .O(n9691));
  LUT3 #(.INIT(8'h96)) lut_n9692 (.I0(n9661), .I1(n9669), .I2(n9670), .O(n9692));
  LUT3 #(.INIT(8'hE8)) lut_n9693 (.I0(n9683), .I1(n9691), .I2(n9692), .O(n9693));
  LUT3 #(.INIT(8'h96)) lut_n9694 (.I0(x630), .I1(x631), .I2(x632), .O(n9694));
  LUT5 #(.INIT(32'h96696996)) lut_n9695 (.I0(x621), .I1(x622), .I2(x623), .I3(n9687), .I4(n9688), .O(n9695));
  LUT5 #(.INIT(32'hFF969600)) lut_n9696 (.I0(x627), .I1(x628), .I2(x629), .I3(n9694), .I4(n9695), .O(n9696));
  LUT3 #(.INIT(8'h96)) lut_n9697 (.I0(x636), .I1(x637), .I2(x638), .O(n9697));
  LUT5 #(.INIT(32'h96696996)) lut_n9698 (.I0(x627), .I1(x628), .I2(x629), .I3(n9694), .I4(n9695), .O(n9698));
  LUT5 #(.INIT(32'hFF969600)) lut_n9699 (.I0(x633), .I1(x634), .I2(x635), .I3(n9697), .I4(n9698), .O(n9699));
  LUT3 #(.INIT(8'h96)) lut_n9700 (.I0(n9686), .I1(n9689), .I2(n9690), .O(n9700));
  LUT3 #(.INIT(8'hE8)) lut_n9701 (.I0(n9696), .I1(n9699), .I2(n9700), .O(n9701));
  LUT3 #(.INIT(8'h96)) lut_n9702 (.I0(x642), .I1(x643), .I2(x644), .O(n9702));
  LUT5 #(.INIT(32'h96696996)) lut_n9703 (.I0(x633), .I1(x634), .I2(x635), .I3(n9697), .I4(n9698), .O(n9703));
  LUT5 #(.INIT(32'hFF969600)) lut_n9704 (.I0(x639), .I1(x640), .I2(x641), .I3(n9702), .I4(n9703), .O(n9704));
  LUT3 #(.INIT(8'h96)) lut_n9705 (.I0(x648), .I1(x649), .I2(x650), .O(n9705));
  LUT5 #(.INIT(32'h96696996)) lut_n9706 (.I0(x639), .I1(x640), .I2(x641), .I3(n9702), .I4(n9703), .O(n9706));
  LUT5 #(.INIT(32'hFF969600)) lut_n9707 (.I0(x645), .I1(x646), .I2(x647), .I3(n9705), .I4(n9706), .O(n9707));
  LUT3 #(.INIT(8'h96)) lut_n9708 (.I0(n9696), .I1(n9699), .I2(n9700), .O(n9708));
  LUT3 #(.INIT(8'hE8)) lut_n9709 (.I0(n9704), .I1(n9707), .I2(n9708), .O(n9709));
  LUT3 #(.INIT(8'h96)) lut_n9710 (.I0(n9683), .I1(n9691), .I2(n9692), .O(n9710));
  LUT3 #(.INIT(8'hE8)) lut_n9711 (.I0(n9701), .I1(n9709), .I2(n9710), .O(n9711));
  LUT3 #(.INIT(8'h96)) lut_n9712 (.I0(n9653), .I1(n9671), .I2(n9672), .O(n9712));
  LUT3 #(.INIT(8'hE8)) lut_n9713 (.I0(n9693), .I1(n9711), .I2(n9712), .O(n9713));
  LUT3 #(.INIT(8'h96)) lut_n9714 (.I0(x654), .I1(x655), .I2(x656), .O(n9714));
  LUT5 #(.INIT(32'h96696996)) lut_n9715 (.I0(x645), .I1(x646), .I2(x647), .I3(n9705), .I4(n9706), .O(n9715));
  LUT5 #(.INIT(32'hFF969600)) lut_n9716 (.I0(x651), .I1(x652), .I2(x653), .I3(n9714), .I4(n9715), .O(n9716));
  LUT3 #(.INIT(8'h96)) lut_n9717 (.I0(x660), .I1(x661), .I2(x662), .O(n9717));
  LUT5 #(.INIT(32'h96696996)) lut_n9718 (.I0(x651), .I1(x652), .I2(x653), .I3(n9714), .I4(n9715), .O(n9718));
  LUT5 #(.INIT(32'hFF969600)) lut_n9719 (.I0(x657), .I1(x658), .I2(x659), .I3(n9717), .I4(n9718), .O(n9719));
  LUT3 #(.INIT(8'h96)) lut_n9720 (.I0(n9704), .I1(n9707), .I2(n9708), .O(n9720));
  LUT3 #(.INIT(8'hE8)) lut_n9721 (.I0(n9716), .I1(n9719), .I2(n9720), .O(n9721));
  LUT3 #(.INIT(8'h96)) lut_n9722 (.I0(x666), .I1(x667), .I2(x668), .O(n9722));
  LUT5 #(.INIT(32'h96696996)) lut_n9723 (.I0(x657), .I1(x658), .I2(x659), .I3(n9717), .I4(n9718), .O(n9723));
  LUT5 #(.INIT(32'hFF969600)) lut_n9724 (.I0(x663), .I1(x664), .I2(x665), .I3(n9722), .I4(n9723), .O(n9724));
  LUT3 #(.INIT(8'h96)) lut_n9725 (.I0(x672), .I1(x673), .I2(x674), .O(n9725));
  LUT5 #(.INIT(32'h96696996)) lut_n9726 (.I0(x663), .I1(x664), .I2(x665), .I3(n9722), .I4(n9723), .O(n9726));
  LUT5 #(.INIT(32'hFF969600)) lut_n9727 (.I0(x669), .I1(x670), .I2(x671), .I3(n9725), .I4(n9726), .O(n9727));
  LUT3 #(.INIT(8'h96)) lut_n9728 (.I0(n9716), .I1(n9719), .I2(n9720), .O(n9728));
  LUT3 #(.INIT(8'hE8)) lut_n9729 (.I0(n9724), .I1(n9727), .I2(n9728), .O(n9729));
  LUT3 #(.INIT(8'h96)) lut_n9730 (.I0(n9701), .I1(n9709), .I2(n9710), .O(n9730));
  LUT3 #(.INIT(8'hE8)) lut_n9731 (.I0(n9721), .I1(n9729), .I2(n9730), .O(n9731));
  LUT3 #(.INIT(8'h96)) lut_n9732 (.I0(x678), .I1(x679), .I2(x680), .O(n9732));
  LUT5 #(.INIT(32'h96696996)) lut_n9733 (.I0(x669), .I1(x670), .I2(x671), .I3(n9725), .I4(n9726), .O(n9733));
  LUT5 #(.INIT(32'hFF969600)) lut_n9734 (.I0(x675), .I1(x676), .I2(x677), .I3(n9732), .I4(n9733), .O(n9734));
  LUT3 #(.INIT(8'h96)) lut_n9735 (.I0(x684), .I1(x685), .I2(x686), .O(n9735));
  LUT5 #(.INIT(32'h96696996)) lut_n9736 (.I0(x675), .I1(x676), .I2(x677), .I3(n9732), .I4(n9733), .O(n9736));
  LUT5 #(.INIT(32'hFF969600)) lut_n9737 (.I0(x681), .I1(x682), .I2(x683), .I3(n9735), .I4(n9736), .O(n9737));
  LUT3 #(.INIT(8'h96)) lut_n9738 (.I0(n9724), .I1(n9727), .I2(n9728), .O(n9738));
  LUT3 #(.INIT(8'hE8)) lut_n9739 (.I0(n9734), .I1(n9737), .I2(n9738), .O(n9739));
  LUT3 #(.INIT(8'h96)) lut_n9740 (.I0(x690), .I1(x691), .I2(x692), .O(n9740));
  LUT5 #(.INIT(32'h96696996)) lut_n9741 (.I0(x681), .I1(x682), .I2(x683), .I3(n9735), .I4(n9736), .O(n9741));
  LUT5 #(.INIT(32'hFF969600)) lut_n9742 (.I0(x687), .I1(x688), .I2(x689), .I3(n9740), .I4(n9741), .O(n9742));
  LUT3 #(.INIT(8'h96)) lut_n9743 (.I0(x696), .I1(x697), .I2(x698), .O(n9743));
  LUT5 #(.INIT(32'h96696996)) lut_n9744 (.I0(x687), .I1(x688), .I2(x689), .I3(n9740), .I4(n9741), .O(n9744));
  LUT5 #(.INIT(32'hFF969600)) lut_n9745 (.I0(x693), .I1(x694), .I2(x695), .I3(n9743), .I4(n9744), .O(n9745));
  LUT3 #(.INIT(8'h96)) lut_n9746 (.I0(n9734), .I1(n9737), .I2(n9738), .O(n9746));
  LUT3 #(.INIT(8'hE8)) lut_n9747 (.I0(n9742), .I1(n9745), .I2(n9746), .O(n9747));
  LUT3 #(.INIT(8'h96)) lut_n9748 (.I0(n9721), .I1(n9729), .I2(n9730), .O(n9748));
  LUT3 #(.INIT(8'hE8)) lut_n9749 (.I0(n9739), .I1(n9747), .I2(n9748), .O(n9749));
  LUT3 #(.INIT(8'h96)) lut_n9750 (.I0(n9693), .I1(n9711), .I2(n9712), .O(n9750));
  LUT3 #(.INIT(8'hE8)) lut_n9751 (.I0(n9731), .I1(n9749), .I2(n9750), .O(n9751));
  LUT3 #(.INIT(8'h96)) lut_n9752 (.I0(n9635), .I1(n9673), .I2(n9674), .O(n9752));
  LUT3 #(.INIT(8'hE8)) lut_n9753 (.I0(n9713), .I1(n9751), .I2(n9752), .O(n9753));
  LUT3 #(.INIT(8'h96)) lut_n9754 (.I0(n9517), .I1(n9595), .I2(n9596), .O(n9754));
  LUT3 #(.INIT(8'hE8)) lut_n9755 (.I0(n9675), .I1(n9753), .I2(n9754), .O(n9755));
  LUT3 #(.INIT(8'h96)) lut_n9756 (.I0(n9279), .I1(n9437), .I2(n9438), .O(n9756));
  LUT3 #(.INIT(8'hE8)) lut_n9757 (.I0(n9597), .I1(n9755), .I2(n9756), .O(n9757));
  LUT3 #(.INIT(8'h96)) lut_n9758 (.I0(n8991), .I1(n9149), .I2(n9150), .O(n9758));
  LUT3 #(.INIT(8'hE8)) lut_n9759 (.I0(n9439), .I1(n9757), .I2(n9758), .O(n9759));
  LUT3 #(.INIT(8'h96)) lut_n9760 (.I0(n8511), .I1(n8829), .I2(n8830), .O(n9760));
  LUT3 #(.INIT(8'hE8)) lut_n9761 (.I0(n9151), .I1(n9759), .I2(n9760), .O(n9761));
  LUT3 #(.INIT(8'h96)) lut_n9762 (.I0(x702), .I1(x703), .I2(x704), .O(n9762));
  LUT5 #(.INIT(32'h96696996)) lut_n9763 (.I0(x693), .I1(x694), .I2(x695), .I3(n9743), .I4(n9744), .O(n9763));
  LUT5 #(.INIT(32'hFF969600)) lut_n9764 (.I0(x699), .I1(x700), .I2(x701), .I3(n9762), .I4(n9763), .O(n9764));
  LUT3 #(.INIT(8'h96)) lut_n9765 (.I0(x708), .I1(x709), .I2(x710), .O(n9765));
  LUT5 #(.INIT(32'h96696996)) lut_n9766 (.I0(x699), .I1(x700), .I2(x701), .I3(n9762), .I4(n9763), .O(n9766));
  LUT5 #(.INIT(32'hFF969600)) lut_n9767 (.I0(x705), .I1(x706), .I2(x707), .I3(n9765), .I4(n9766), .O(n9767));
  LUT3 #(.INIT(8'h96)) lut_n9768 (.I0(n9742), .I1(n9745), .I2(n9746), .O(n9768));
  LUT3 #(.INIT(8'hE8)) lut_n9769 (.I0(n9764), .I1(n9767), .I2(n9768), .O(n9769));
  LUT3 #(.INIT(8'h96)) lut_n9770 (.I0(x714), .I1(x715), .I2(x716), .O(n9770));
  LUT5 #(.INIT(32'h96696996)) lut_n9771 (.I0(x705), .I1(x706), .I2(x707), .I3(n9765), .I4(n9766), .O(n9771));
  LUT5 #(.INIT(32'hFF969600)) lut_n9772 (.I0(x711), .I1(x712), .I2(x713), .I3(n9770), .I4(n9771), .O(n9772));
  LUT3 #(.INIT(8'h96)) lut_n9773 (.I0(x720), .I1(x721), .I2(x722), .O(n9773));
  LUT5 #(.INIT(32'h96696996)) lut_n9774 (.I0(x711), .I1(x712), .I2(x713), .I3(n9770), .I4(n9771), .O(n9774));
  LUT5 #(.INIT(32'hFF969600)) lut_n9775 (.I0(x717), .I1(x718), .I2(x719), .I3(n9773), .I4(n9774), .O(n9775));
  LUT3 #(.INIT(8'h96)) lut_n9776 (.I0(n9764), .I1(n9767), .I2(n9768), .O(n9776));
  LUT3 #(.INIT(8'hE8)) lut_n9777 (.I0(n9772), .I1(n9775), .I2(n9776), .O(n9777));
  LUT3 #(.INIT(8'h96)) lut_n9778 (.I0(n9739), .I1(n9747), .I2(n9748), .O(n9778));
  LUT3 #(.INIT(8'hE8)) lut_n9779 (.I0(n9769), .I1(n9777), .I2(n9778), .O(n9779));
  LUT3 #(.INIT(8'h96)) lut_n9780 (.I0(x726), .I1(x727), .I2(x728), .O(n9780));
  LUT5 #(.INIT(32'h96696996)) lut_n9781 (.I0(x717), .I1(x718), .I2(x719), .I3(n9773), .I4(n9774), .O(n9781));
  LUT5 #(.INIT(32'hFF969600)) lut_n9782 (.I0(x723), .I1(x724), .I2(x725), .I3(n9780), .I4(n9781), .O(n9782));
  LUT3 #(.INIT(8'h96)) lut_n9783 (.I0(x732), .I1(x733), .I2(x734), .O(n9783));
  LUT5 #(.INIT(32'h96696996)) lut_n9784 (.I0(x723), .I1(x724), .I2(x725), .I3(n9780), .I4(n9781), .O(n9784));
  LUT5 #(.INIT(32'hFF969600)) lut_n9785 (.I0(x729), .I1(x730), .I2(x731), .I3(n9783), .I4(n9784), .O(n9785));
  LUT3 #(.INIT(8'h96)) lut_n9786 (.I0(n9772), .I1(n9775), .I2(n9776), .O(n9786));
  LUT3 #(.INIT(8'hE8)) lut_n9787 (.I0(n9782), .I1(n9785), .I2(n9786), .O(n9787));
  LUT3 #(.INIT(8'h96)) lut_n9788 (.I0(x738), .I1(x739), .I2(x740), .O(n9788));
  LUT5 #(.INIT(32'h96696996)) lut_n9789 (.I0(x729), .I1(x730), .I2(x731), .I3(n9783), .I4(n9784), .O(n9789));
  LUT5 #(.INIT(32'hFF969600)) lut_n9790 (.I0(x735), .I1(x736), .I2(x737), .I3(n9788), .I4(n9789), .O(n9790));
  LUT3 #(.INIT(8'h96)) lut_n9791 (.I0(x744), .I1(x745), .I2(x746), .O(n9791));
  LUT5 #(.INIT(32'h96696996)) lut_n9792 (.I0(x735), .I1(x736), .I2(x737), .I3(n9788), .I4(n9789), .O(n9792));
  LUT5 #(.INIT(32'hFF969600)) lut_n9793 (.I0(x741), .I1(x742), .I2(x743), .I3(n9791), .I4(n9792), .O(n9793));
  LUT3 #(.INIT(8'h96)) lut_n9794 (.I0(n9782), .I1(n9785), .I2(n9786), .O(n9794));
  LUT3 #(.INIT(8'hE8)) lut_n9795 (.I0(n9790), .I1(n9793), .I2(n9794), .O(n9795));
  LUT3 #(.INIT(8'h96)) lut_n9796 (.I0(n9769), .I1(n9777), .I2(n9778), .O(n9796));
  LUT3 #(.INIT(8'hE8)) lut_n9797 (.I0(n9787), .I1(n9795), .I2(n9796), .O(n9797));
  LUT3 #(.INIT(8'h96)) lut_n9798 (.I0(n9731), .I1(n9749), .I2(n9750), .O(n9798));
  LUT3 #(.INIT(8'hE8)) lut_n9799 (.I0(n9779), .I1(n9797), .I2(n9798), .O(n9799));
  LUT3 #(.INIT(8'h96)) lut_n9800 (.I0(x750), .I1(x751), .I2(x752), .O(n9800));
  LUT5 #(.INIT(32'h96696996)) lut_n9801 (.I0(x741), .I1(x742), .I2(x743), .I3(n9791), .I4(n9792), .O(n9801));
  LUT5 #(.INIT(32'hFF969600)) lut_n9802 (.I0(x747), .I1(x748), .I2(x749), .I3(n9800), .I4(n9801), .O(n9802));
  LUT3 #(.INIT(8'h96)) lut_n9803 (.I0(x756), .I1(x757), .I2(x758), .O(n9803));
  LUT5 #(.INIT(32'h96696996)) lut_n9804 (.I0(x747), .I1(x748), .I2(x749), .I3(n9800), .I4(n9801), .O(n9804));
  LUT5 #(.INIT(32'hFF969600)) lut_n9805 (.I0(x753), .I1(x754), .I2(x755), .I3(n9803), .I4(n9804), .O(n9805));
  LUT3 #(.INIT(8'h96)) lut_n9806 (.I0(n9790), .I1(n9793), .I2(n9794), .O(n9806));
  LUT3 #(.INIT(8'hE8)) lut_n9807 (.I0(n9802), .I1(n9805), .I2(n9806), .O(n9807));
  LUT3 #(.INIT(8'h96)) lut_n9808 (.I0(x762), .I1(x763), .I2(x764), .O(n9808));
  LUT5 #(.INIT(32'h96696996)) lut_n9809 (.I0(x753), .I1(x754), .I2(x755), .I3(n9803), .I4(n9804), .O(n9809));
  LUT5 #(.INIT(32'hFF969600)) lut_n9810 (.I0(x759), .I1(x760), .I2(x761), .I3(n9808), .I4(n9809), .O(n9810));
  LUT3 #(.INIT(8'h96)) lut_n9811 (.I0(x768), .I1(x769), .I2(x770), .O(n9811));
  LUT5 #(.INIT(32'h96696996)) lut_n9812 (.I0(x759), .I1(x760), .I2(x761), .I3(n9808), .I4(n9809), .O(n9812));
  LUT5 #(.INIT(32'hFF969600)) lut_n9813 (.I0(x765), .I1(x766), .I2(x767), .I3(n9811), .I4(n9812), .O(n9813));
  LUT3 #(.INIT(8'h96)) lut_n9814 (.I0(n9802), .I1(n9805), .I2(n9806), .O(n9814));
  LUT3 #(.INIT(8'hE8)) lut_n9815 (.I0(n9810), .I1(n9813), .I2(n9814), .O(n9815));
  LUT3 #(.INIT(8'h96)) lut_n9816 (.I0(n9787), .I1(n9795), .I2(n9796), .O(n9816));
  LUT3 #(.INIT(8'hE8)) lut_n9817 (.I0(n9807), .I1(n9815), .I2(n9816), .O(n9817));
  LUT3 #(.INIT(8'h96)) lut_n9818 (.I0(x774), .I1(x775), .I2(x776), .O(n9818));
  LUT5 #(.INIT(32'h96696996)) lut_n9819 (.I0(x765), .I1(x766), .I2(x767), .I3(n9811), .I4(n9812), .O(n9819));
  LUT5 #(.INIT(32'hFF969600)) lut_n9820 (.I0(x771), .I1(x772), .I2(x773), .I3(n9818), .I4(n9819), .O(n9820));
  LUT3 #(.INIT(8'h96)) lut_n9821 (.I0(x780), .I1(x781), .I2(x782), .O(n9821));
  LUT5 #(.INIT(32'h96696996)) lut_n9822 (.I0(x771), .I1(x772), .I2(x773), .I3(n9818), .I4(n9819), .O(n9822));
  LUT5 #(.INIT(32'hFF969600)) lut_n9823 (.I0(x777), .I1(x778), .I2(x779), .I3(n9821), .I4(n9822), .O(n9823));
  LUT3 #(.INIT(8'h96)) lut_n9824 (.I0(n9810), .I1(n9813), .I2(n9814), .O(n9824));
  LUT3 #(.INIT(8'hE8)) lut_n9825 (.I0(n9820), .I1(n9823), .I2(n9824), .O(n9825));
  LUT3 #(.INIT(8'h96)) lut_n9826 (.I0(x786), .I1(x787), .I2(x788), .O(n9826));
  LUT5 #(.INIT(32'h96696996)) lut_n9827 (.I0(x777), .I1(x778), .I2(x779), .I3(n9821), .I4(n9822), .O(n9827));
  LUT5 #(.INIT(32'hFF969600)) lut_n9828 (.I0(x783), .I1(x784), .I2(x785), .I3(n9826), .I4(n9827), .O(n9828));
  LUT3 #(.INIT(8'h96)) lut_n9829 (.I0(x792), .I1(x793), .I2(x794), .O(n9829));
  LUT5 #(.INIT(32'h96696996)) lut_n9830 (.I0(x783), .I1(x784), .I2(x785), .I3(n9826), .I4(n9827), .O(n9830));
  LUT5 #(.INIT(32'hFF969600)) lut_n9831 (.I0(x789), .I1(x790), .I2(x791), .I3(n9829), .I4(n9830), .O(n9831));
  LUT3 #(.INIT(8'h96)) lut_n9832 (.I0(n9820), .I1(n9823), .I2(n9824), .O(n9832));
  LUT3 #(.INIT(8'hE8)) lut_n9833 (.I0(n9828), .I1(n9831), .I2(n9832), .O(n9833));
  LUT3 #(.INIT(8'h96)) lut_n9834 (.I0(n9807), .I1(n9815), .I2(n9816), .O(n9834));
  LUT3 #(.INIT(8'hE8)) lut_n9835 (.I0(n9825), .I1(n9833), .I2(n9834), .O(n9835));
  LUT3 #(.INIT(8'h96)) lut_n9836 (.I0(n9779), .I1(n9797), .I2(n9798), .O(n9836));
  LUT3 #(.INIT(8'hE8)) lut_n9837 (.I0(n9817), .I1(n9835), .I2(n9836), .O(n9837));
  LUT3 #(.INIT(8'h96)) lut_n9838 (.I0(n9713), .I1(n9751), .I2(n9752), .O(n9838));
  LUT3 #(.INIT(8'hE8)) lut_n9839 (.I0(n9799), .I1(n9837), .I2(n9838), .O(n9839));
  LUT3 #(.INIT(8'h96)) lut_n9840 (.I0(x798), .I1(x799), .I2(x800), .O(n9840));
  LUT5 #(.INIT(32'h96696996)) lut_n9841 (.I0(x789), .I1(x790), .I2(x791), .I3(n9829), .I4(n9830), .O(n9841));
  LUT5 #(.INIT(32'hFF969600)) lut_n9842 (.I0(x795), .I1(x796), .I2(x797), .I3(n9840), .I4(n9841), .O(n9842));
  LUT3 #(.INIT(8'h96)) lut_n9843 (.I0(x804), .I1(x805), .I2(x806), .O(n9843));
  LUT5 #(.INIT(32'h96696996)) lut_n9844 (.I0(x795), .I1(x796), .I2(x797), .I3(n9840), .I4(n9841), .O(n9844));
  LUT5 #(.INIT(32'hFF969600)) lut_n9845 (.I0(x801), .I1(x802), .I2(x803), .I3(n9843), .I4(n9844), .O(n9845));
  LUT3 #(.INIT(8'h96)) lut_n9846 (.I0(n9828), .I1(n9831), .I2(n9832), .O(n9846));
  LUT3 #(.INIT(8'hE8)) lut_n9847 (.I0(n9842), .I1(n9845), .I2(n9846), .O(n9847));
  LUT3 #(.INIT(8'h96)) lut_n9848 (.I0(x810), .I1(x811), .I2(x812), .O(n9848));
  LUT5 #(.INIT(32'h96696996)) lut_n9849 (.I0(x801), .I1(x802), .I2(x803), .I3(n9843), .I4(n9844), .O(n9849));
  LUT5 #(.INIT(32'hFF969600)) lut_n9850 (.I0(x807), .I1(x808), .I2(x809), .I3(n9848), .I4(n9849), .O(n9850));
  LUT3 #(.INIT(8'h96)) lut_n9851 (.I0(x816), .I1(x817), .I2(x818), .O(n9851));
  LUT5 #(.INIT(32'h96696996)) lut_n9852 (.I0(x807), .I1(x808), .I2(x809), .I3(n9848), .I4(n9849), .O(n9852));
  LUT5 #(.INIT(32'hFF969600)) lut_n9853 (.I0(x813), .I1(x814), .I2(x815), .I3(n9851), .I4(n9852), .O(n9853));
  LUT3 #(.INIT(8'h96)) lut_n9854 (.I0(n9842), .I1(n9845), .I2(n9846), .O(n9854));
  LUT3 #(.INIT(8'hE8)) lut_n9855 (.I0(n9850), .I1(n9853), .I2(n9854), .O(n9855));
  LUT3 #(.INIT(8'h96)) lut_n9856 (.I0(n9825), .I1(n9833), .I2(n9834), .O(n9856));
  LUT3 #(.INIT(8'hE8)) lut_n9857 (.I0(n9847), .I1(n9855), .I2(n9856), .O(n9857));
  LUT3 #(.INIT(8'h96)) lut_n9858 (.I0(x822), .I1(x823), .I2(x824), .O(n9858));
  LUT5 #(.INIT(32'h96696996)) lut_n9859 (.I0(x813), .I1(x814), .I2(x815), .I3(n9851), .I4(n9852), .O(n9859));
  LUT5 #(.INIT(32'hFF969600)) lut_n9860 (.I0(x819), .I1(x820), .I2(x821), .I3(n9858), .I4(n9859), .O(n9860));
  LUT3 #(.INIT(8'h96)) lut_n9861 (.I0(x828), .I1(x829), .I2(x830), .O(n9861));
  LUT5 #(.INIT(32'h96696996)) lut_n9862 (.I0(x819), .I1(x820), .I2(x821), .I3(n9858), .I4(n9859), .O(n9862));
  LUT5 #(.INIT(32'hFF969600)) lut_n9863 (.I0(x825), .I1(x826), .I2(x827), .I3(n9861), .I4(n9862), .O(n9863));
  LUT3 #(.INIT(8'h96)) lut_n9864 (.I0(n9850), .I1(n9853), .I2(n9854), .O(n9864));
  LUT3 #(.INIT(8'hE8)) lut_n9865 (.I0(n9860), .I1(n9863), .I2(n9864), .O(n9865));
  LUT3 #(.INIT(8'h96)) lut_n9866 (.I0(x834), .I1(x835), .I2(x836), .O(n9866));
  LUT5 #(.INIT(32'h96696996)) lut_n9867 (.I0(x825), .I1(x826), .I2(x827), .I3(n9861), .I4(n9862), .O(n9867));
  LUT5 #(.INIT(32'hFF969600)) lut_n9868 (.I0(x831), .I1(x832), .I2(x833), .I3(n9866), .I4(n9867), .O(n9868));
  LUT3 #(.INIT(8'h96)) lut_n9869 (.I0(x840), .I1(x841), .I2(x842), .O(n9869));
  LUT5 #(.INIT(32'h96696996)) lut_n9870 (.I0(x831), .I1(x832), .I2(x833), .I3(n9866), .I4(n9867), .O(n9870));
  LUT5 #(.INIT(32'hFF969600)) lut_n9871 (.I0(x837), .I1(x838), .I2(x839), .I3(n9869), .I4(n9870), .O(n9871));
  LUT3 #(.INIT(8'h96)) lut_n9872 (.I0(n9860), .I1(n9863), .I2(n9864), .O(n9872));
  LUT3 #(.INIT(8'hE8)) lut_n9873 (.I0(n9868), .I1(n9871), .I2(n9872), .O(n9873));
  LUT3 #(.INIT(8'h96)) lut_n9874 (.I0(n9847), .I1(n9855), .I2(n9856), .O(n9874));
  LUT3 #(.INIT(8'hE8)) lut_n9875 (.I0(n9865), .I1(n9873), .I2(n9874), .O(n9875));
  LUT3 #(.INIT(8'h96)) lut_n9876 (.I0(n9817), .I1(n9835), .I2(n9836), .O(n9876));
  LUT3 #(.INIT(8'hE8)) lut_n9877 (.I0(n9857), .I1(n9875), .I2(n9876), .O(n9877));
  LUT3 #(.INIT(8'h96)) lut_n9878 (.I0(x846), .I1(x847), .I2(x848), .O(n9878));
  LUT5 #(.INIT(32'h96696996)) lut_n9879 (.I0(x837), .I1(x838), .I2(x839), .I3(n9869), .I4(n9870), .O(n9879));
  LUT5 #(.INIT(32'hFF969600)) lut_n9880 (.I0(x843), .I1(x844), .I2(x845), .I3(n9878), .I4(n9879), .O(n9880));
  LUT3 #(.INIT(8'h96)) lut_n9881 (.I0(x852), .I1(x853), .I2(x854), .O(n9881));
  LUT5 #(.INIT(32'h96696996)) lut_n9882 (.I0(x843), .I1(x844), .I2(x845), .I3(n9878), .I4(n9879), .O(n9882));
  LUT5 #(.INIT(32'hFF969600)) lut_n9883 (.I0(x849), .I1(x850), .I2(x851), .I3(n9881), .I4(n9882), .O(n9883));
  LUT3 #(.INIT(8'h96)) lut_n9884 (.I0(n9868), .I1(n9871), .I2(n9872), .O(n9884));
  LUT3 #(.INIT(8'hE8)) lut_n9885 (.I0(n9880), .I1(n9883), .I2(n9884), .O(n9885));
  LUT3 #(.INIT(8'h96)) lut_n9886 (.I0(x858), .I1(x859), .I2(x860), .O(n9886));
  LUT5 #(.INIT(32'h96696996)) lut_n9887 (.I0(x849), .I1(x850), .I2(x851), .I3(n9881), .I4(n9882), .O(n9887));
  LUT5 #(.INIT(32'hFF969600)) lut_n9888 (.I0(x855), .I1(x856), .I2(x857), .I3(n9886), .I4(n9887), .O(n9888));
  LUT3 #(.INIT(8'h96)) lut_n9889 (.I0(x864), .I1(x865), .I2(x866), .O(n9889));
  LUT5 #(.INIT(32'h96696996)) lut_n9890 (.I0(x855), .I1(x856), .I2(x857), .I3(n9886), .I4(n9887), .O(n9890));
  LUT5 #(.INIT(32'hFF969600)) lut_n9891 (.I0(x861), .I1(x862), .I2(x863), .I3(n9889), .I4(n9890), .O(n9891));
  LUT3 #(.INIT(8'h96)) lut_n9892 (.I0(n9880), .I1(n9883), .I2(n9884), .O(n9892));
  LUT3 #(.INIT(8'hE8)) lut_n9893 (.I0(n9888), .I1(n9891), .I2(n9892), .O(n9893));
  LUT3 #(.INIT(8'h96)) lut_n9894 (.I0(n9865), .I1(n9873), .I2(n9874), .O(n9894));
  LUT3 #(.INIT(8'hE8)) lut_n9895 (.I0(n9885), .I1(n9893), .I2(n9894), .O(n9895));
  LUT3 #(.INIT(8'h96)) lut_n9896 (.I0(x870), .I1(x871), .I2(x872), .O(n9896));
  LUT5 #(.INIT(32'h96696996)) lut_n9897 (.I0(x861), .I1(x862), .I2(x863), .I3(n9889), .I4(n9890), .O(n9897));
  LUT5 #(.INIT(32'hFF969600)) lut_n9898 (.I0(x867), .I1(x868), .I2(x869), .I3(n9896), .I4(n9897), .O(n9898));
  LUT3 #(.INIT(8'h96)) lut_n9899 (.I0(x876), .I1(x877), .I2(x878), .O(n9899));
  LUT5 #(.INIT(32'h96696996)) lut_n9900 (.I0(x867), .I1(x868), .I2(x869), .I3(n9896), .I4(n9897), .O(n9900));
  LUT5 #(.INIT(32'hFF969600)) lut_n9901 (.I0(x873), .I1(x874), .I2(x875), .I3(n9899), .I4(n9900), .O(n9901));
  LUT3 #(.INIT(8'h96)) lut_n9902 (.I0(n9888), .I1(n9891), .I2(n9892), .O(n9902));
  LUT3 #(.INIT(8'hE8)) lut_n9903 (.I0(n9898), .I1(n9901), .I2(n9902), .O(n9903));
  LUT3 #(.INIT(8'h96)) lut_n9904 (.I0(x882), .I1(x883), .I2(x884), .O(n9904));
  LUT5 #(.INIT(32'h96696996)) lut_n9905 (.I0(x873), .I1(x874), .I2(x875), .I3(n9899), .I4(n9900), .O(n9905));
  LUT5 #(.INIT(32'hFF969600)) lut_n9906 (.I0(x879), .I1(x880), .I2(x881), .I3(n9904), .I4(n9905), .O(n9906));
  LUT3 #(.INIT(8'h96)) lut_n9907 (.I0(x888), .I1(x889), .I2(x890), .O(n9907));
  LUT5 #(.INIT(32'h96696996)) lut_n9908 (.I0(x879), .I1(x880), .I2(x881), .I3(n9904), .I4(n9905), .O(n9908));
  LUT5 #(.INIT(32'hFF969600)) lut_n9909 (.I0(x885), .I1(x886), .I2(x887), .I3(n9907), .I4(n9908), .O(n9909));
  LUT3 #(.INIT(8'h96)) lut_n9910 (.I0(n9898), .I1(n9901), .I2(n9902), .O(n9910));
  LUT3 #(.INIT(8'hE8)) lut_n9911 (.I0(n9906), .I1(n9909), .I2(n9910), .O(n9911));
  LUT3 #(.INIT(8'h96)) lut_n9912 (.I0(n9885), .I1(n9893), .I2(n9894), .O(n9912));
  LUT3 #(.INIT(8'hE8)) lut_n9913 (.I0(n9903), .I1(n9911), .I2(n9912), .O(n9913));
  LUT3 #(.INIT(8'h96)) lut_n9914 (.I0(n9857), .I1(n9875), .I2(n9876), .O(n9914));
  LUT3 #(.INIT(8'hE8)) lut_n9915 (.I0(n9895), .I1(n9913), .I2(n9914), .O(n9915));
  LUT3 #(.INIT(8'h96)) lut_n9916 (.I0(n9799), .I1(n9837), .I2(n9838), .O(n9916));
  LUT3 #(.INIT(8'hE8)) lut_n9917 (.I0(n9877), .I1(n9915), .I2(n9916), .O(n9917));
  LUT3 #(.INIT(8'h96)) lut_n9918 (.I0(n9675), .I1(n9753), .I2(n9754), .O(n9918));
  LUT3 #(.INIT(8'hE8)) lut_n9919 (.I0(n9839), .I1(n9917), .I2(n9918), .O(n9919));
  LUT3 #(.INIT(8'h96)) lut_n9920 (.I0(x894), .I1(x895), .I2(x896), .O(n9920));
  LUT5 #(.INIT(32'h96696996)) lut_n9921 (.I0(x885), .I1(x886), .I2(x887), .I3(n9907), .I4(n9908), .O(n9921));
  LUT5 #(.INIT(32'hFF969600)) lut_n9922 (.I0(x891), .I1(x892), .I2(x893), .I3(n9920), .I4(n9921), .O(n9922));
  LUT3 #(.INIT(8'h96)) lut_n9923 (.I0(x900), .I1(x901), .I2(x902), .O(n9923));
  LUT5 #(.INIT(32'h96696996)) lut_n9924 (.I0(x891), .I1(x892), .I2(x893), .I3(n9920), .I4(n9921), .O(n9924));
  LUT5 #(.INIT(32'hFF969600)) lut_n9925 (.I0(x897), .I1(x898), .I2(x899), .I3(n9923), .I4(n9924), .O(n9925));
  LUT3 #(.INIT(8'h96)) lut_n9926 (.I0(n9906), .I1(n9909), .I2(n9910), .O(n9926));
  LUT3 #(.INIT(8'hE8)) lut_n9927 (.I0(n9922), .I1(n9925), .I2(n9926), .O(n9927));
  LUT3 #(.INIT(8'h96)) lut_n9928 (.I0(x906), .I1(x907), .I2(x908), .O(n9928));
  LUT5 #(.INIT(32'h96696996)) lut_n9929 (.I0(x897), .I1(x898), .I2(x899), .I3(n9923), .I4(n9924), .O(n9929));
  LUT5 #(.INIT(32'hFF969600)) lut_n9930 (.I0(x903), .I1(x904), .I2(x905), .I3(n9928), .I4(n9929), .O(n9930));
  LUT3 #(.INIT(8'h96)) lut_n9931 (.I0(x912), .I1(x913), .I2(x914), .O(n9931));
  LUT5 #(.INIT(32'h96696996)) lut_n9932 (.I0(x903), .I1(x904), .I2(x905), .I3(n9928), .I4(n9929), .O(n9932));
  LUT5 #(.INIT(32'hFF969600)) lut_n9933 (.I0(x909), .I1(x910), .I2(x911), .I3(n9931), .I4(n9932), .O(n9933));
  LUT3 #(.INIT(8'h96)) lut_n9934 (.I0(n9922), .I1(n9925), .I2(n9926), .O(n9934));
  LUT3 #(.INIT(8'hE8)) lut_n9935 (.I0(n9930), .I1(n9933), .I2(n9934), .O(n9935));
  LUT3 #(.INIT(8'h96)) lut_n9936 (.I0(n9903), .I1(n9911), .I2(n9912), .O(n9936));
  LUT3 #(.INIT(8'hE8)) lut_n9937 (.I0(n9927), .I1(n9935), .I2(n9936), .O(n9937));
  LUT3 #(.INIT(8'h96)) lut_n9938 (.I0(x918), .I1(x919), .I2(x920), .O(n9938));
  LUT5 #(.INIT(32'h96696996)) lut_n9939 (.I0(x909), .I1(x910), .I2(x911), .I3(n9931), .I4(n9932), .O(n9939));
  LUT5 #(.INIT(32'hFF969600)) lut_n9940 (.I0(x915), .I1(x916), .I2(x917), .I3(n9938), .I4(n9939), .O(n9940));
  LUT3 #(.INIT(8'h96)) lut_n9941 (.I0(x924), .I1(x925), .I2(x926), .O(n9941));
  LUT5 #(.INIT(32'h96696996)) lut_n9942 (.I0(x915), .I1(x916), .I2(x917), .I3(n9938), .I4(n9939), .O(n9942));
  LUT5 #(.INIT(32'hFF969600)) lut_n9943 (.I0(x921), .I1(x922), .I2(x923), .I3(n9941), .I4(n9942), .O(n9943));
  LUT3 #(.INIT(8'h96)) lut_n9944 (.I0(n9930), .I1(n9933), .I2(n9934), .O(n9944));
  LUT3 #(.INIT(8'hE8)) lut_n9945 (.I0(n9940), .I1(n9943), .I2(n9944), .O(n9945));
  LUT3 #(.INIT(8'h96)) lut_n9946 (.I0(x930), .I1(x931), .I2(x932), .O(n9946));
  LUT5 #(.INIT(32'h96696996)) lut_n9947 (.I0(x921), .I1(x922), .I2(x923), .I3(n9941), .I4(n9942), .O(n9947));
  LUT5 #(.INIT(32'hFF969600)) lut_n9948 (.I0(x927), .I1(x928), .I2(x929), .I3(n9946), .I4(n9947), .O(n9948));
  LUT3 #(.INIT(8'h96)) lut_n9949 (.I0(x936), .I1(x937), .I2(x938), .O(n9949));
  LUT5 #(.INIT(32'h96696996)) lut_n9950 (.I0(x927), .I1(x928), .I2(x929), .I3(n9946), .I4(n9947), .O(n9950));
  LUT5 #(.INIT(32'hFF969600)) lut_n9951 (.I0(x933), .I1(x934), .I2(x935), .I3(n9949), .I4(n9950), .O(n9951));
  LUT3 #(.INIT(8'h96)) lut_n9952 (.I0(n9940), .I1(n9943), .I2(n9944), .O(n9952));
  LUT3 #(.INIT(8'hE8)) lut_n9953 (.I0(n9948), .I1(n9951), .I2(n9952), .O(n9953));
  LUT3 #(.INIT(8'h96)) lut_n9954 (.I0(n9927), .I1(n9935), .I2(n9936), .O(n9954));
  LUT3 #(.INIT(8'hE8)) lut_n9955 (.I0(n9945), .I1(n9953), .I2(n9954), .O(n9955));
  LUT3 #(.INIT(8'h96)) lut_n9956 (.I0(n9895), .I1(n9913), .I2(n9914), .O(n9956));
  LUT3 #(.INIT(8'hE8)) lut_n9957 (.I0(n9937), .I1(n9955), .I2(n9956), .O(n9957));
  LUT3 #(.INIT(8'h96)) lut_n9958 (.I0(x942), .I1(x943), .I2(x944), .O(n9958));
  LUT5 #(.INIT(32'h96696996)) lut_n9959 (.I0(x933), .I1(x934), .I2(x935), .I3(n9949), .I4(n9950), .O(n9959));
  LUT5 #(.INIT(32'hFF969600)) lut_n9960 (.I0(x939), .I1(x940), .I2(x941), .I3(n9958), .I4(n9959), .O(n9960));
  LUT3 #(.INIT(8'h96)) lut_n9961 (.I0(x948), .I1(x949), .I2(x950), .O(n9961));
  LUT5 #(.INIT(32'h96696996)) lut_n9962 (.I0(x939), .I1(x940), .I2(x941), .I3(n9958), .I4(n9959), .O(n9962));
  LUT5 #(.INIT(32'hFF969600)) lut_n9963 (.I0(x945), .I1(x946), .I2(x947), .I3(n9961), .I4(n9962), .O(n9963));
  LUT3 #(.INIT(8'h96)) lut_n9964 (.I0(n9948), .I1(n9951), .I2(n9952), .O(n9964));
  LUT3 #(.INIT(8'hE8)) lut_n9965 (.I0(n9960), .I1(n9963), .I2(n9964), .O(n9965));
  LUT3 #(.INIT(8'h96)) lut_n9966 (.I0(x954), .I1(x955), .I2(x956), .O(n9966));
  LUT5 #(.INIT(32'h96696996)) lut_n9967 (.I0(x945), .I1(x946), .I2(x947), .I3(n9961), .I4(n9962), .O(n9967));
  LUT5 #(.INIT(32'hFF969600)) lut_n9968 (.I0(x951), .I1(x952), .I2(x953), .I3(n9966), .I4(n9967), .O(n9968));
  LUT3 #(.INIT(8'h96)) lut_n9969 (.I0(x960), .I1(x961), .I2(x962), .O(n9969));
  LUT5 #(.INIT(32'h96696996)) lut_n9970 (.I0(x951), .I1(x952), .I2(x953), .I3(n9966), .I4(n9967), .O(n9970));
  LUT5 #(.INIT(32'hFF969600)) lut_n9971 (.I0(x957), .I1(x958), .I2(x959), .I3(n9969), .I4(n9970), .O(n9971));
  LUT3 #(.INIT(8'h96)) lut_n9972 (.I0(n9960), .I1(n9963), .I2(n9964), .O(n9972));
  LUT3 #(.INIT(8'hE8)) lut_n9973 (.I0(n9968), .I1(n9971), .I2(n9972), .O(n9973));
  LUT3 #(.INIT(8'h96)) lut_n9974 (.I0(n9945), .I1(n9953), .I2(n9954), .O(n9974));
  LUT3 #(.INIT(8'hE8)) lut_n9975 (.I0(n9965), .I1(n9973), .I2(n9974), .O(n9975));
  LUT3 #(.INIT(8'h96)) lut_n9976 (.I0(x966), .I1(x967), .I2(x968), .O(n9976));
  LUT5 #(.INIT(32'h96696996)) lut_n9977 (.I0(x957), .I1(x958), .I2(x959), .I3(n9969), .I4(n9970), .O(n9977));
  LUT5 #(.INIT(32'hFF969600)) lut_n9978 (.I0(x963), .I1(x964), .I2(x965), .I3(n9976), .I4(n9977), .O(n9978));
  LUT3 #(.INIT(8'h96)) lut_n9979 (.I0(x972), .I1(x973), .I2(x974), .O(n9979));
  LUT5 #(.INIT(32'h96696996)) lut_n9980 (.I0(x963), .I1(x964), .I2(x965), .I3(n9976), .I4(n9977), .O(n9980));
  LUT5 #(.INIT(32'hFF969600)) lut_n9981 (.I0(x969), .I1(x970), .I2(x971), .I3(n9979), .I4(n9980), .O(n9981));
  LUT3 #(.INIT(8'h96)) lut_n9982 (.I0(n9968), .I1(n9971), .I2(n9972), .O(n9982));
  LUT3 #(.INIT(8'hE8)) lut_n9983 (.I0(n9978), .I1(n9981), .I2(n9982), .O(n9983));
  LUT3 #(.INIT(8'h96)) lut_n9984 (.I0(x978), .I1(x979), .I2(x980), .O(n9984));
  LUT5 #(.INIT(32'h96696996)) lut_n9985 (.I0(x969), .I1(x970), .I2(x971), .I3(n9979), .I4(n9980), .O(n9985));
  LUT5 #(.INIT(32'hFF969600)) lut_n9986 (.I0(x975), .I1(x976), .I2(x977), .I3(n9984), .I4(n9985), .O(n9986));
  LUT3 #(.INIT(8'h96)) lut_n9987 (.I0(x984), .I1(x985), .I2(x986), .O(n9987));
  LUT5 #(.INIT(32'h96696996)) lut_n9988 (.I0(x975), .I1(x976), .I2(x977), .I3(n9984), .I4(n9985), .O(n9988));
  LUT5 #(.INIT(32'hFF969600)) lut_n9989 (.I0(x981), .I1(x982), .I2(x983), .I3(n9987), .I4(n9988), .O(n9989));
  LUT3 #(.INIT(8'h96)) lut_n9990 (.I0(n9978), .I1(n9981), .I2(n9982), .O(n9990));
  LUT3 #(.INIT(8'hE8)) lut_n9991 (.I0(n9986), .I1(n9989), .I2(n9990), .O(n9991));
  LUT3 #(.INIT(8'h96)) lut_n9992 (.I0(n9965), .I1(n9973), .I2(n9974), .O(n9992));
  LUT3 #(.INIT(8'hE8)) lut_n9993 (.I0(n9983), .I1(n9991), .I2(n9992), .O(n9993));
  LUT3 #(.INIT(8'h96)) lut_n9994 (.I0(n9937), .I1(n9955), .I2(n9956), .O(n9994));
  LUT3 #(.INIT(8'hE8)) lut_n9995 (.I0(n9975), .I1(n9993), .I2(n9994), .O(n9995));
  LUT3 #(.INIT(8'h96)) lut_n9996 (.I0(n9877), .I1(n9915), .I2(n9916), .O(n9996));
  LUT3 #(.INIT(8'hE8)) lut_n9997 (.I0(n9957), .I1(n9995), .I2(n9996), .O(n9997));
  LUT3 #(.INIT(8'h96)) lut_n9998 (.I0(x990), .I1(x991), .I2(x992), .O(n9998));
  LUT5 #(.INIT(32'h96696996)) lut_n9999 (.I0(x981), .I1(x982), .I2(x983), .I3(n9987), .I4(n9988), .O(n9999));
  LUT5 #(.INIT(32'hFF969600)) lut_n10000 (.I0(x987), .I1(x988), .I2(x989), .I3(n9998), .I4(n9999), .O(n10000));
  LUT3 #(.INIT(8'h96)) lut_n10001 (.I0(x996), .I1(x997), .I2(x998), .O(n10001));
  LUT5 #(.INIT(32'h96696996)) lut_n10002 (.I0(x987), .I1(x988), .I2(x989), .I3(n9998), .I4(n9999), .O(n10002));
  LUT5 #(.INIT(32'hFF969600)) lut_n10003 (.I0(x993), .I1(x994), .I2(x995), .I3(n10001), .I4(n10002), .O(n10003));
  LUT3 #(.INIT(8'h96)) lut_n10004 (.I0(n9986), .I1(n9989), .I2(n9990), .O(n10004));
  LUT3 #(.INIT(8'hE8)) lut_n10005 (.I0(n10000), .I1(n10003), .I2(n10004), .O(n10005));
  LUT3 #(.INIT(8'h96)) lut_n10006 (.I0(x1002), .I1(x1003), .I2(x1004), .O(n10006));
  LUT5 #(.INIT(32'h96696996)) lut_n10007 (.I0(x993), .I1(x994), .I2(x995), .I3(n10001), .I4(n10002), .O(n10007));
  LUT5 #(.INIT(32'hFF969600)) lut_n10008 (.I0(x999), .I1(x1000), .I2(x1001), .I3(n10006), .I4(n10007), .O(n10008));
  LUT3 #(.INIT(8'h96)) lut_n10009 (.I0(x1008), .I1(x1009), .I2(x1010), .O(n10009));
  LUT5 #(.INIT(32'h96696996)) lut_n10010 (.I0(x999), .I1(x1000), .I2(x1001), .I3(n10006), .I4(n10007), .O(n10010));
  LUT5 #(.INIT(32'hFF969600)) lut_n10011 (.I0(x1005), .I1(x1006), .I2(x1007), .I3(n10009), .I4(n10010), .O(n10011));
  LUT3 #(.INIT(8'h96)) lut_n10012 (.I0(n10000), .I1(n10003), .I2(n10004), .O(n10012));
  LUT3 #(.INIT(8'hE8)) lut_n10013 (.I0(n10008), .I1(n10011), .I2(n10012), .O(n10013));
  LUT3 #(.INIT(8'h96)) lut_n10014 (.I0(n9983), .I1(n9991), .I2(n9992), .O(n10014));
  LUT3 #(.INIT(8'hE8)) lut_n10015 (.I0(n10005), .I1(n10013), .I2(n10014), .O(n10015));
  LUT3 #(.INIT(8'h96)) lut_n10016 (.I0(x1014), .I1(x1015), .I2(x1016), .O(n10016));
  LUT5 #(.INIT(32'h96696996)) lut_n10017 (.I0(x1005), .I1(x1006), .I2(x1007), .I3(n10009), .I4(n10010), .O(n10017));
  LUT5 #(.INIT(32'hFF969600)) lut_n10018 (.I0(x1011), .I1(x1012), .I2(x1013), .I3(n10016), .I4(n10017), .O(n10018));
  LUT3 #(.INIT(8'h96)) lut_n10019 (.I0(x1020), .I1(x1021), .I2(x1022), .O(n10019));
  LUT5 #(.INIT(32'h96696996)) lut_n10020 (.I0(x1011), .I1(x1012), .I2(x1013), .I3(n10016), .I4(n10017), .O(n10020));
  LUT5 #(.INIT(32'hFF969600)) lut_n10021 (.I0(x1017), .I1(x1018), .I2(x1019), .I3(n10019), .I4(n10020), .O(n10021));
  LUT3 #(.INIT(8'h96)) lut_n10022 (.I0(n10008), .I1(n10011), .I2(n10012), .O(n10022));
  LUT3 #(.INIT(8'hE8)) lut_n10023 (.I0(n10018), .I1(n10021), .I2(n10022), .O(n10023));
  LUT3 #(.INIT(8'h96)) lut_n10024 (.I0(x1026), .I1(x1027), .I2(x1028), .O(n10024));
  LUT5 #(.INIT(32'h96696996)) lut_n10025 (.I0(x1017), .I1(x1018), .I2(x1019), .I3(n10019), .I4(n10020), .O(n10025));
  LUT5 #(.INIT(32'hFF969600)) lut_n10026 (.I0(x1023), .I1(x1024), .I2(x1025), .I3(n10024), .I4(n10025), .O(n10026));
  LUT3 #(.INIT(8'h96)) lut_n10027 (.I0(x1032), .I1(x1033), .I2(x1034), .O(n10027));
  LUT5 #(.INIT(32'h96696996)) lut_n10028 (.I0(x1023), .I1(x1024), .I2(x1025), .I3(n10024), .I4(n10025), .O(n10028));
  LUT5 #(.INIT(32'hFF969600)) lut_n10029 (.I0(x1029), .I1(x1030), .I2(x1031), .I3(n10027), .I4(n10028), .O(n10029));
  LUT3 #(.INIT(8'h96)) lut_n10030 (.I0(n10018), .I1(n10021), .I2(n10022), .O(n10030));
  LUT3 #(.INIT(8'hE8)) lut_n10031 (.I0(n10026), .I1(n10029), .I2(n10030), .O(n10031));
  LUT3 #(.INIT(8'h96)) lut_n10032 (.I0(n10005), .I1(n10013), .I2(n10014), .O(n10032));
  LUT3 #(.INIT(8'hE8)) lut_n10033 (.I0(n10023), .I1(n10031), .I2(n10032), .O(n10033));
  LUT3 #(.INIT(8'h96)) lut_n10034 (.I0(n9975), .I1(n9993), .I2(n9994), .O(n10034));
  LUT3 #(.INIT(8'hE8)) lut_n10035 (.I0(n10015), .I1(n10033), .I2(n10034), .O(n10035));
  LUT3 #(.INIT(8'h96)) lut_n10036 (.I0(x1038), .I1(x1039), .I2(x1040), .O(n10036));
  LUT5 #(.INIT(32'h96696996)) lut_n10037 (.I0(x1029), .I1(x1030), .I2(x1031), .I3(n10027), .I4(n10028), .O(n10037));
  LUT5 #(.INIT(32'hFF969600)) lut_n10038 (.I0(x1035), .I1(x1036), .I2(x1037), .I3(n10036), .I4(n10037), .O(n10038));
  LUT3 #(.INIT(8'h96)) lut_n10039 (.I0(x1044), .I1(x1045), .I2(x1046), .O(n10039));
  LUT5 #(.INIT(32'h96696996)) lut_n10040 (.I0(x1035), .I1(x1036), .I2(x1037), .I3(n10036), .I4(n10037), .O(n10040));
  LUT5 #(.INIT(32'hFF969600)) lut_n10041 (.I0(x1041), .I1(x1042), .I2(x1043), .I3(n10039), .I4(n10040), .O(n10041));
  LUT3 #(.INIT(8'h96)) lut_n10042 (.I0(n10026), .I1(n10029), .I2(n10030), .O(n10042));
  LUT3 #(.INIT(8'hE8)) lut_n10043 (.I0(n10038), .I1(n10041), .I2(n10042), .O(n10043));
  LUT3 #(.INIT(8'h96)) lut_n10044 (.I0(x1050), .I1(x1051), .I2(x1052), .O(n10044));
  LUT5 #(.INIT(32'h96696996)) lut_n10045 (.I0(x1041), .I1(x1042), .I2(x1043), .I3(n10039), .I4(n10040), .O(n10045));
  LUT5 #(.INIT(32'hFF969600)) lut_n10046 (.I0(x1047), .I1(x1048), .I2(x1049), .I3(n10044), .I4(n10045), .O(n10046));
  LUT3 #(.INIT(8'h96)) lut_n10047 (.I0(x1056), .I1(x1057), .I2(x1058), .O(n10047));
  LUT5 #(.INIT(32'h96696996)) lut_n10048 (.I0(x1047), .I1(x1048), .I2(x1049), .I3(n10044), .I4(n10045), .O(n10048));
  LUT5 #(.INIT(32'hFF969600)) lut_n10049 (.I0(x1053), .I1(x1054), .I2(x1055), .I3(n10047), .I4(n10048), .O(n10049));
  LUT3 #(.INIT(8'h96)) lut_n10050 (.I0(n10038), .I1(n10041), .I2(n10042), .O(n10050));
  LUT3 #(.INIT(8'hE8)) lut_n10051 (.I0(n10046), .I1(n10049), .I2(n10050), .O(n10051));
  LUT3 #(.INIT(8'h96)) lut_n10052 (.I0(n10023), .I1(n10031), .I2(n10032), .O(n10052));
  LUT3 #(.INIT(8'hE8)) lut_n10053 (.I0(n10043), .I1(n10051), .I2(n10052), .O(n10053));
  LUT3 #(.INIT(8'h96)) lut_n10054 (.I0(x1062), .I1(x1063), .I2(x1064), .O(n10054));
  LUT5 #(.INIT(32'h96696996)) lut_n10055 (.I0(x1053), .I1(x1054), .I2(x1055), .I3(n10047), .I4(n10048), .O(n10055));
  LUT5 #(.INIT(32'hFF969600)) lut_n10056 (.I0(x1059), .I1(x1060), .I2(x1061), .I3(n10054), .I4(n10055), .O(n10056));
  LUT3 #(.INIT(8'h96)) lut_n10057 (.I0(x1068), .I1(x1069), .I2(x1070), .O(n10057));
  LUT5 #(.INIT(32'h96696996)) lut_n10058 (.I0(x1059), .I1(x1060), .I2(x1061), .I3(n10054), .I4(n10055), .O(n10058));
  LUT5 #(.INIT(32'hFF969600)) lut_n10059 (.I0(x1065), .I1(x1066), .I2(x1067), .I3(n10057), .I4(n10058), .O(n10059));
  LUT3 #(.INIT(8'h96)) lut_n10060 (.I0(n10046), .I1(n10049), .I2(n10050), .O(n10060));
  LUT3 #(.INIT(8'hE8)) lut_n10061 (.I0(n10056), .I1(n10059), .I2(n10060), .O(n10061));
  LUT3 #(.INIT(8'h96)) lut_n10062 (.I0(x1074), .I1(x1075), .I2(x1076), .O(n10062));
  LUT5 #(.INIT(32'h96696996)) lut_n10063 (.I0(x1065), .I1(x1066), .I2(x1067), .I3(n10057), .I4(n10058), .O(n10063));
  LUT5 #(.INIT(32'hFF969600)) lut_n10064 (.I0(x1071), .I1(x1072), .I2(x1073), .I3(n10062), .I4(n10063), .O(n10064));
  LUT3 #(.INIT(8'h96)) lut_n10065 (.I0(x1080), .I1(x1081), .I2(x1082), .O(n10065));
  LUT5 #(.INIT(32'h96696996)) lut_n10066 (.I0(x1071), .I1(x1072), .I2(x1073), .I3(n10062), .I4(n10063), .O(n10066));
  LUT5 #(.INIT(32'hFF969600)) lut_n10067 (.I0(x1077), .I1(x1078), .I2(x1079), .I3(n10065), .I4(n10066), .O(n10067));
  LUT3 #(.INIT(8'h96)) lut_n10068 (.I0(n10056), .I1(n10059), .I2(n10060), .O(n10068));
  LUT3 #(.INIT(8'hE8)) lut_n10069 (.I0(n10064), .I1(n10067), .I2(n10068), .O(n10069));
  LUT3 #(.INIT(8'h96)) lut_n10070 (.I0(n10043), .I1(n10051), .I2(n10052), .O(n10070));
  LUT3 #(.INIT(8'hE8)) lut_n10071 (.I0(n10061), .I1(n10069), .I2(n10070), .O(n10071));
  LUT3 #(.INIT(8'h96)) lut_n10072 (.I0(n10015), .I1(n10033), .I2(n10034), .O(n10072));
  LUT3 #(.INIT(8'hE8)) lut_n10073 (.I0(n10053), .I1(n10071), .I2(n10072), .O(n10073));
  LUT3 #(.INIT(8'h96)) lut_n10074 (.I0(n9957), .I1(n9995), .I2(n9996), .O(n10074));
  LUT3 #(.INIT(8'hE8)) lut_n10075 (.I0(n10035), .I1(n10073), .I2(n10074), .O(n10075));
  LUT3 #(.INIT(8'h96)) lut_n10076 (.I0(n9839), .I1(n9917), .I2(n9918), .O(n10076));
  LUT3 #(.INIT(8'hE8)) lut_n10077 (.I0(n9997), .I1(n10075), .I2(n10076), .O(n10077));
  LUT3 #(.INIT(8'h96)) lut_n10078 (.I0(n9597), .I1(n9755), .I2(n9756), .O(n10078));
  LUT3 #(.INIT(8'hE8)) lut_n10079 (.I0(n9919), .I1(n10077), .I2(n10078), .O(n10079));
  LUT3 #(.INIT(8'h96)) lut_n10080 (.I0(x1086), .I1(x1087), .I2(x1088), .O(n10080));
  LUT5 #(.INIT(32'h96696996)) lut_n10081 (.I0(x1077), .I1(x1078), .I2(x1079), .I3(n10065), .I4(n10066), .O(n10081));
  LUT5 #(.INIT(32'hFF969600)) lut_n10082 (.I0(x1083), .I1(x1084), .I2(x1085), .I3(n10080), .I4(n10081), .O(n10082));
  LUT3 #(.INIT(8'h96)) lut_n10083 (.I0(x1092), .I1(x1093), .I2(x1094), .O(n10083));
  LUT5 #(.INIT(32'h96696996)) lut_n10084 (.I0(x1083), .I1(x1084), .I2(x1085), .I3(n10080), .I4(n10081), .O(n10084));
  LUT5 #(.INIT(32'hFF969600)) lut_n10085 (.I0(x1089), .I1(x1090), .I2(x1091), .I3(n10083), .I4(n10084), .O(n10085));
  LUT3 #(.INIT(8'h96)) lut_n10086 (.I0(n10064), .I1(n10067), .I2(n10068), .O(n10086));
  LUT3 #(.INIT(8'hE8)) lut_n10087 (.I0(n10082), .I1(n10085), .I2(n10086), .O(n10087));
  LUT3 #(.INIT(8'h96)) lut_n10088 (.I0(x1098), .I1(x1099), .I2(x1100), .O(n10088));
  LUT5 #(.INIT(32'h96696996)) lut_n10089 (.I0(x1089), .I1(x1090), .I2(x1091), .I3(n10083), .I4(n10084), .O(n10089));
  LUT5 #(.INIT(32'hFF969600)) lut_n10090 (.I0(x1095), .I1(x1096), .I2(x1097), .I3(n10088), .I4(n10089), .O(n10090));
  LUT3 #(.INIT(8'h96)) lut_n10091 (.I0(x1104), .I1(x1105), .I2(x1106), .O(n10091));
  LUT5 #(.INIT(32'h96696996)) lut_n10092 (.I0(x1095), .I1(x1096), .I2(x1097), .I3(n10088), .I4(n10089), .O(n10092));
  LUT5 #(.INIT(32'hFF969600)) lut_n10093 (.I0(x1101), .I1(x1102), .I2(x1103), .I3(n10091), .I4(n10092), .O(n10093));
  LUT3 #(.INIT(8'h96)) lut_n10094 (.I0(n10082), .I1(n10085), .I2(n10086), .O(n10094));
  LUT3 #(.INIT(8'hE8)) lut_n10095 (.I0(n10090), .I1(n10093), .I2(n10094), .O(n10095));
  LUT3 #(.INIT(8'h96)) lut_n10096 (.I0(n10061), .I1(n10069), .I2(n10070), .O(n10096));
  LUT3 #(.INIT(8'hE8)) lut_n10097 (.I0(n10087), .I1(n10095), .I2(n10096), .O(n10097));
  LUT3 #(.INIT(8'h96)) lut_n10098 (.I0(x1110), .I1(x1111), .I2(x1112), .O(n10098));
  LUT5 #(.INIT(32'h96696996)) lut_n10099 (.I0(x1101), .I1(x1102), .I2(x1103), .I3(n10091), .I4(n10092), .O(n10099));
  LUT5 #(.INIT(32'hFF969600)) lut_n10100 (.I0(x1107), .I1(x1108), .I2(x1109), .I3(n10098), .I4(n10099), .O(n10100));
  LUT3 #(.INIT(8'h96)) lut_n10101 (.I0(x1116), .I1(x1117), .I2(x1118), .O(n10101));
  LUT5 #(.INIT(32'h96696996)) lut_n10102 (.I0(x1107), .I1(x1108), .I2(x1109), .I3(n10098), .I4(n10099), .O(n10102));
  LUT5 #(.INIT(32'hFF969600)) lut_n10103 (.I0(x1113), .I1(x1114), .I2(x1115), .I3(n10101), .I4(n10102), .O(n10103));
  LUT3 #(.INIT(8'h96)) lut_n10104 (.I0(n10090), .I1(n10093), .I2(n10094), .O(n10104));
  LUT3 #(.INIT(8'hE8)) lut_n10105 (.I0(n10100), .I1(n10103), .I2(n10104), .O(n10105));
  LUT3 #(.INIT(8'h96)) lut_n10106 (.I0(x1122), .I1(x1123), .I2(x1124), .O(n10106));
  LUT5 #(.INIT(32'h96696996)) lut_n10107 (.I0(x1113), .I1(x1114), .I2(x1115), .I3(n10101), .I4(n10102), .O(n10107));
  LUT5 #(.INIT(32'hFF969600)) lut_n10108 (.I0(x1119), .I1(x1120), .I2(x1121), .I3(n10106), .I4(n10107), .O(n10108));
  LUT3 #(.INIT(8'h96)) lut_n10109 (.I0(x1128), .I1(x1129), .I2(x1130), .O(n10109));
  LUT5 #(.INIT(32'h96696996)) lut_n10110 (.I0(x1119), .I1(x1120), .I2(x1121), .I3(n10106), .I4(n10107), .O(n10110));
  LUT5 #(.INIT(32'hFF969600)) lut_n10111 (.I0(x1125), .I1(x1126), .I2(x1127), .I3(n10109), .I4(n10110), .O(n10111));
  LUT3 #(.INIT(8'h96)) lut_n10112 (.I0(n10100), .I1(n10103), .I2(n10104), .O(n10112));
  LUT3 #(.INIT(8'hE8)) lut_n10113 (.I0(n10108), .I1(n10111), .I2(n10112), .O(n10113));
  LUT3 #(.INIT(8'h96)) lut_n10114 (.I0(n10087), .I1(n10095), .I2(n10096), .O(n10114));
  LUT3 #(.INIT(8'hE8)) lut_n10115 (.I0(n10105), .I1(n10113), .I2(n10114), .O(n10115));
  LUT3 #(.INIT(8'h96)) lut_n10116 (.I0(n10053), .I1(n10071), .I2(n10072), .O(n10116));
  LUT3 #(.INIT(8'hE8)) lut_n10117 (.I0(n10097), .I1(n10115), .I2(n10116), .O(n10117));
  LUT3 #(.INIT(8'h96)) lut_n10118 (.I0(x1134), .I1(x1135), .I2(x1136), .O(n10118));
  LUT5 #(.INIT(32'h96696996)) lut_n10119 (.I0(x1125), .I1(x1126), .I2(x1127), .I3(n10109), .I4(n10110), .O(n10119));
  LUT5 #(.INIT(32'hFF969600)) lut_n10120 (.I0(x1131), .I1(x1132), .I2(x1133), .I3(n10118), .I4(n10119), .O(n10120));
  LUT3 #(.INIT(8'h96)) lut_n10121 (.I0(x1140), .I1(x1141), .I2(x1142), .O(n10121));
  LUT5 #(.INIT(32'h96696996)) lut_n10122 (.I0(x1131), .I1(x1132), .I2(x1133), .I3(n10118), .I4(n10119), .O(n10122));
  LUT5 #(.INIT(32'hFF969600)) lut_n10123 (.I0(x1137), .I1(x1138), .I2(x1139), .I3(n10121), .I4(n10122), .O(n10123));
  LUT3 #(.INIT(8'h96)) lut_n10124 (.I0(n10108), .I1(n10111), .I2(n10112), .O(n10124));
  LUT3 #(.INIT(8'hE8)) lut_n10125 (.I0(n10120), .I1(n10123), .I2(n10124), .O(n10125));
  LUT3 #(.INIT(8'h96)) lut_n10126 (.I0(x1146), .I1(x1147), .I2(x1148), .O(n10126));
  LUT5 #(.INIT(32'h96696996)) lut_n10127 (.I0(x1137), .I1(x1138), .I2(x1139), .I3(n10121), .I4(n10122), .O(n10127));
  LUT5 #(.INIT(32'hFF969600)) lut_n10128 (.I0(x1143), .I1(x1144), .I2(x1145), .I3(n10126), .I4(n10127), .O(n10128));
  LUT3 #(.INIT(8'h96)) lut_n10129 (.I0(x1152), .I1(x1153), .I2(x1154), .O(n10129));
  LUT5 #(.INIT(32'h96696996)) lut_n10130 (.I0(x1143), .I1(x1144), .I2(x1145), .I3(n10126), .I4(n10127), .O(n10130));
  LUT5 #(.INIT(32'hFF969600)) lut_n10131 (.I0(x1149), .I1(x1150), .I2(x1151), .I3(n10129), .I4(n10130), .O(n10131));
  LUT3 #(.INIT(8'h96)) lut_n10132 (.I0(n10120), .I1(n10123), .I2(n10124), .O(n10132));
  LUT3 #(.INIT(8'hE8)) lut_n10133 (.I0(n10128), .I1(n10131), .I2(n10132), .O(n10133));
  LUT3 #(.INIT(8'h96)) lut_n10134 (.I0(n10105), .I1(n10113), .I2(n10114), .O(n10134));
  LUT3 #(.INIT(8'hE8)) lut_n10135 (.I0(n10125), .I1(n10133), .I2(n10134), .O(n10135));
  LUT3 #(.INIT(8'h96)) lut_n10136 (.I0(x1158), .I1(x1159), .I2(x1160), .O(n10136));
  LUT5 #(.INIT(32'h96696996)) lut_n10137 (.I0(x1149), .I1(x1150), .I2(x1151), .I3(n10129), .I4(n10130), .O(n10137));
  LUT5 #(.INIT(32'hFF969600)) lut_n10138 (.I0(x1155), .I1(x1156), .I2(x1157), .I3(n10136), .I4(n10137), .O(n10138));
  LUT3 #(.INIT(8'h96)) lut_n10139 (.I0(x1164), .I1(x1165), .I2(x1166), .O(n10139));
  LUT5 #(.INIT(32'h96696996)) lut_n10140 (.I0(x1155), .I1(x1156), .I2(x1157), .I3(n10136), .I4(n10137), .O(n10140));
  LUT5 #(.INIT(32'hFF969600)) lut_n10141 (.I0(x1161), .I1(x1162), .I2(x1163), .I3(n10139), .I4(n10140), .O(n10141));
  LUT3 #(.INIT(8'h96)) lut_n10142 (.I0(n10128), .I1(n10131), .I2(n10132), .O(n10142));
  LUT3 #(.INIT(8'hE8)) lut_n10143 (.I0(n10138), .I1(n10141), .I2(n10142), .O(n10143));
  LUT3 #(.INIT(8'h96)) lut_n10144 (.I0(x1170), .I1(x1171), .I2(x1172), .O(n10144));
  LUT5 #(.INIT(32'h96696996)) lut_n10145 (.I0(x1161), .I1(x1162), .I2(x1163), .I3(n10139), .I4(n10140), .O(n10145));
  LUT5 #(.INIT(32'hFF969600)) lut_n10146 (.I0(x1167), .I1(x1168), .I2(x1169), .I3(n10144), .I4(n10145), .O(n10146));
  LUT3 #(.INIT(8'h96)) lut_n10147 (.I0(x1176), .I1(x1177), .I2(x1178), .O(n10147));
  LUT5 #(.INIT(32'h96696996)) lut_n10148 (.I0(x1167), .I1(x1168), .I2(x1169), .I3(n10144), .I4(n10145), .O(n10148));
  LUT5 #(.INIT(32'hFF969600)) lut_n10149 (.I0(x1173), .I1(x1174), .I2(x1175), .I3(n10147), .I4(n10148), .O(n10149));
  LUT3 #(.INIT(8'h96)) lut_n10150 (.I0(n10138), .I1(n10141), .I2(n10142), .O(n10150));
  LUT3 #(.INIT(8'hE8)) lut_n10151 (.I0(n10146), .I1(n10149), .I2(n10150), .O(n10151));
  LUT3 #(.INIT(8'h96)) lut_n10152 (.I0(n10125), .I1(n10133), .I2(n10134), .O(n10152));
  LUT3 #(.INIT(8'hE8)) lut_n10153 (.I0(n10143), .I1(n10151), .I2(n10152), .O(n10153));
  LUT3 #(.INIT(8'h96)) lut_n10154 (.I0(n10097), .I1(n10115), .I2(n10116), .O(n10154));
  LUT3 #(.INIT(8'hE8)) lut_n10155 (.I0(n10135), .I1(n10153), .I2(n10154), .O(n10155));
  LUT3 #(.INIT(8'h96)) lut_n10156 (.I0(n10035), .I1(n10073), .I2(n10074), .O(n10156));
  LUT3 #(.INIT(8'hE8)) lut_n10157 (.I0(n10117), .I1(n10155), .I2(n10156), .O(n10157));
  LUT3 #(.INIT(8'h96)) lut_n10158 (.I0(x1182), .I1(x1183), .I2(x1184), .O(n10158));
  LUT5 #(.INIT(32'h96696996)) lut_n10159 (.I0(x1173), .I1(x1174), .I2(x1175), .I3(n10147), .I4(n10148), .O(n10159));
  LUT5 #(.INIT(32'hFF969600)) lut_n10160 (.I0(x1179), .I1(x1180), .I2(x1181), .I3(n10158), .I4(n10159), .O(n10160));
  LUT3 #(.INIT(8'h96)) lut_n10161 (.I0(x1188), .I1(x1189), .I2(x1190), .O(n10161));
  LUT5 #(.INIT(32'h96696996)) lut_n10162 (.I0(x1179), .I1(x1180), .I2(x1181), .I3(n10158), .I4(n10159), .O(n10162));
  LUT5 #(.INIT(32'hFF969600)) lut_n10163 (.I0(x1185), .I1(x1186), .I2(x1187), .I3(n10161), .I4(n10162), .O(n10163));
  LUT3 #(.INIT(8'h96)) lut_n10164 (.I0(n10146), .I1(n10149), .I2(n10150), .O(n10164));
  LUT3 #(.INIT(8'hE8)) lut_n10165 (.I0(n10160), .I1(n10163), .I2(n10164), .O(n10165));
  LUT3 #(.INIT(8'h96)) lut_n10166 (.I0(x1194), .I1(x1195), .I2(x1196), .O(n10166));
  LUT5 #(.INIT(32'h96696996)) lut_n10167 (.I0(x1185), .I1(x1186), .I2(x1187), .I3(n10161), .I4(n10162), .O(n10167));
  LUT5 #(.INIT(32'hFF969600)) lut_n10168 (.I0(x1191), .I1(x1192), .I2(x1193), .I3(n10166), .I4(n10167), .O(n10168));
  LUT3 #(.INIT(8'h96)) lut_n10169 (.I0(x1200), .I1(x1201), .I2(x1202), .O(n10169));
  LUT5 #(.INIT(32'h96696996)) lut_n10170 (.I0(x1191), .I1(x1192), .I2(x1193), .I3(n10166), .I4(n10167), .O(n10170));
  LUT5 #(.INIT(32'hFF969600)) lut_n10171 (.I0(x1197), .I1(x1198), .I2(x1199), .I3(n10169), .I4(n10170), .O(n10171));
  LUT3 #(.INIT(8'h96)) lut_n10172 (.I0(n10160), .I1(n10163), .I2(n10164), .O(n10172));
  LUT3 #(.INIT(8'hE8)) lut_n10173 (.I0(n10168), .I1(n10171), .I2(n10172), .O(n10173));
  LUT3 #(.INIT(8'h96)) lut_n10174 (.I0(n10143), .I1(n10151), .I2(n10152), .O(n10174));
  LUT3 #(.INIT(8'hE8)) lut_n10175 (.I0(n10165), .I1(n10173), .I2(n10174), .O(n10175));
  LUT3 #(.INIT(8'h96)) lut_n10176 (.I0(x1206), .I1(x1207), .I2(x1208), .O(n10176));
  LUT5 #(.INIT(32'h96696996)) lut_n10177 (.I0(x1197), .I1(x1198), .I2(x1199), .I3(n10169), .I4(n10170), .O(n10177));
  LUT5 #(.INIT(32'hFF969600)) lut_n10178 (.I0(x1203), .I1(x1204), .I2(x1205), .I3(n10176), .I4(n10177), .O(n10178));
  LUT3 #(.INIT(8'h96)) lut_n10179 (.I0(x1212), .I1(x1213), .I2(x1214), .O(n10179));
  LUT5 #(.INIT(32'h96696996)) lut_n10180 (.I0(x1203), .I1(x1204), .I2(x1205), .I3(n10176), .I4(n10177), .O(n10180));
  LUT5 #(.INIT(32'hFF969600)) lut_n10181 (.I0(x1209), .I1(x1210), .I2(x1211), .I3(n10179), .I4(n10180), .O(n10181));
  LUT3 #(.INIT(8'h96)) lut_n10182 (.I0(n10168), .I1(n10171), .I2(n10172), .O(n10182));
  LUT3 #(.INIT(8'hE8)) lut_n10183 (.I0(n10178), .I1(n10181), .I2(n10182), .O(n10183));
  LUT3 #(.INIT(8'h96)) lut_n10184 (.I0(x1218), .I1(x1219), .I2(x1220), .O(n10184));
  LUT5 #(.INIT(32'h96696996)) lut_n10185 (.I0(x1209), .I1(x1210), .I2(x1211), .I3(n10179), .I4(n10180), .O(n10185));
  LUT5 #(.INIT(32'hFF969600)) lut_n10186 (.I0(x1215), .I1(x1216), .I2(x1217), .I3(n10184), .I4(n10185), .O(n10186));
  LUT3 #(.INIT(8'h96)) lut_n10187 (.I0(x1224), .I1(x1225), .I2(x1226), .O(n10187));
  LUT5 #(.INIT(32'h96696996)) lut_n10188 (.I0(x1215), .I1(x1216), .I2(x1217), .I3(n10184), .I4(n10185), .O(n10188));
  LUT5 #(.INIT(32'hFF969600)) lut_n10189 (.I0(x1221), .I1(x1222), .I2(x1223), .I3(n10187), .I4(n10188), .O(n10189));
  LUT3 #(.INIT(8'h96)) lut_n10190 (.I0(n10178), .I1(n10181), .I2(n10182), .O(n10190));
  LUT3 #(.INIT(8'hE8)) lut_n10191 (.I0(n10186), .I1(n10189), .I2(n10190), .O(n10191));
  LUT3 #(.INIT(8'h96)) lut_n10192 (.I0(n10165), .I1(n10173), .I2(n10174), .O(n10192));
  LUT3 #(.INIT(8'hE8)) lut_n10193 (.I0(n10183), .I1(n10191), .I2(n10192), .O(n10193));
  LUT3 #(.INIT(8'h96)) lut_n10194 (.I0(n10135), .I1(n10153), .I2(n10154), .O(n10194));
  LUT3 #(.INIT(8'hE8)) lut_n10195 (.I0(n10175), .I1(n10193), .I2(n10194), .O(n10195));
  LUT3 #(.INIT(8'h96)) lut_n10196 (.I0(x1230), .I1(x1231), .I2(x1232), .O(n10196));
  LUT5 #(.INIT(32'h96696996)) lut_n10197 (.I0(x1221), .I1(x1222), .I2(x1223), .I3(n10187), .I4(n10188), .O(n10197));
  LUT5 #(.INIT(32'hFF969600)) lut_n10198 (.I0(x1227), .I1(x1228), .I2(x1229), .I3(n10196), .I4(n10197), .O(n10198));
  LUT3 #(.INIT(8'h96)) lut_n10199 (.I0(x1236), .I1(x1237), .I2(x1238), .O(n10199));
  LUT5 #(.INIT(32'h96696996)) lut_n10200 (.I0(x1227), .I1(x1228), .I2(x1229), .I3(n10196), .I4(n10197), .O(n10200));
  LUT5 #(.INIT(32'hFF969600)) lut_n10201 (.I0(x1233), .I1(x1234), .I2(x1235), .I3(n10199), .I4(n10200), .O(n10201));
  LUT3 #(.INIT(8'h96)) lut_n10202 (.I0(n10186), .I1(n10189), .I2(n10190), .O(n10202));
  LUT3 #(.INIT(8'hE8)) lut_n10203 (.I0(n10198), .I1(n10201), .I2(n10202), .O(n10203));
  LUT3 #(.INIT(8'h96)) lut_n10204 (.I0(x1242), .I1(x1243), .I2(x1244), .O(n10204));
  LUT5 #(.INIT(32'h96696996)) lut_n10205 (.I0(x1233), .I1(x1234), .I2(x1235), .I3(n10199), .I4(n10200), .O(n10205));
  LUT5 #(.INIT(32'hFF969600)) lut_n10206 (.I0(x1239), .I1(x1240), .I2(x1241), .I3(n10204), .I4(n10205), .O(n10206));
  LUT3 #(.INIT(8'h96)) lut_n10207 (.I0(x1248), .I1(x1249), .I2(x1250), .O(n10207));
  LUT5 #(.INIT(32'h96696996)) lut_n10208 (.I0(x1239), .I1(x1240), .I2(x1241), .I3(n10204), .I4(n10205), .O(n10208));
  LUT5 #(.INIT(32'hFF969600)) lut_n10209 (.I0(x1245), .I1(x1246), .I2(x1247), .I3(n10207), .I4(n10208), .O(n10209));
  LUT3 #(.INIT(8'h96)) lut_n10210 (.I0(n10198), .I1(n10201), .I2(n10202), .O(n10210));
  LUT3 #(.INIT(8'hE8)) lut_n10211 (.I0(n10206), .I1(n10209), .I2(n10210), .O(n10211));
  LUT3 #(.INIT(8'h96)) lut_n10212 (.I0(n10183), .I1(n10191), .I2(n10192), .O(n10212));
  LUT3 #(.INIT(8'hE8)) lut_n10213 (.I0(n10203), .I1(n10211), .I2(n10212), .O(n10213));
  LUT3 #(.INIT(8'h96)) lut_n10214 (.I0(x1254), .I1(x1255), .I2(x1256), .O(n10214));
  LUT5 #(.INIT(32'h96696996)) lut_n10215 (.I0(x1245), .I1(x1246), .I2(x1247), .I3(n10207), .I4(n10208), .O(n10215));
  LUT5 #(.INIT(32'hFF969600)) lut_n10216 (.I0(x1251), .I1(x1252), .I2(x1253), .I3(n10214), .I4(n10215), .O(n10216));
  LUT3 #(.INIT(8'h96)) lut_n10217 (.I0(x1260), .I1(x1261), .I2(x1262), .O(n10217));
  LUT5 #(.INIT(32'h96696996)) lut_n10218 (.I0(x1251), .I1(x1252), .I2(x1253), .I3(n10214), .I4(n10215), .O(n10218));
  LUT5 #(.INIT(32'hFF969600)) lut_n10219 (.I0(x1257), .I1(x1258), .I2(x1259), .I3(n10217), .I4(n10218), .O(n10219));
  LUT3 #(.INIT(8'h96)) lut_n10220 (.I0(n10206), .I1(n10209), .I2(n10210), .O(n10220));
  LUT3 #(.INIT(8'hE8)) lut_n10221 (.I0(n10216), .I1(n10219), .I2(n10220), .O(n10221));
  LUT3 #(.INIT(8'h96)) lut_n10222 (.I0(x1266), .I1(x1267), .I2(x1268), .O(n10222));
  LUT5 #(.INIT(32'h96696996)) lut_n10223 (.I0(x1257), .I1(x1258), .I2(x1259), .I3(n10217), .I4(n10218), .O(n10223));
  LUT5 #(.INIT(32'hFF969600)) lut_n10224 (.I0(x1263), .I1(x1264), .I2(x1265), .I3(n10222), .I4(n10223), .O(n10224));
  LUT3 #(.INIT(8'h96)) lut_n10225 (.I0(x1272), .I1(x1273), .I2(x1274), .O(n10225));
  LUT5 #(.INIT(32'h96696996)) lut_n10226 (.I0(x1263), .I1(x1264), .I2(x1265), .I3(n10222), .I4(n10223), .O(n10226));
  LUT5 #(.INIT(32'hFF969600)) lut_n10227 (.I0(x1269), .I1(x1270), .I2(x1271), .I3(n10225), .I4(n10226), .O(n10227));
  LUT3 #(.INIT(8'h96)) lut_n10228 (.I0(n10216), .I1(n10219), .I2(n10220), .O(n10228));
  LUT3 #(.INIT(8'hE8)) lut_n10229 (.I0(n10224), .I1(n10227), .I2(n10228), .O(n10229));
  LUT3 #(.INIT(8'h96)) lut_n10230 (.I0(n10203), .I1(n10211), .I2(n10212), .O(n10230));
  LUT3 #(.INIT(8'hE8)) lut_n10231 (.I0(n10221), .I1(n10229), .I2(n10230), .O(n10231));
  LUT3 #(.INIT(8'h96)) lut_n10232 (.I0(n10175), .I1(n10193), .I2(n10194), .O(n10232));
  LUT3 #(.INIT(8'hE8)) lut_n10233 (.I0(n10213), .I1(n10231), .I2(n10232), .O(n10233));
  LUT3 #(.INIT(8'h96)) lut_n10234 (.I0(n10117), .I1(n10155), .I2(n10156), .O(n10234));
  LUT3 #(.INIT(8'hE8)) lut_n10235 (.I0(n10195), .I1(n10233), .I2(n10234), .O(n10235));
  LUT3 #(.INIT(8'h96)) lut_n10236 (.I0(n9997), .I1(n10075), .I2(n10076), .O(n10236));
  LUT3 #(.INIT(8'hE8)) lut_n10237 (.I0(n10157), .I1(n10235), .I2(n10236), .O(n10237));
  LUT3 #(.INIT(8'h96)) lut_n10238 (.I0(x1278), .I1(x1279), .I2(x1280), .O(n10238));
  LUT5 #(.INIT(32'h96696996)) lut_n10239 (.I0(x1269), .I1(x1270), .I2(x1271), .I3(n10225), .I4(n10226), .O(n10239));
  LUT5 #(.INIT(32'hFF969600)) lut_n10240 (.I0(x1275), .I1(x1276), .I2(x1277), .I3(n10238), .I4(n10239), .O(n10240));
  LUT3 #(.INIT(8'h96)) lut_n10241 (.I0(x1284), .I1(x1285), .I2(x1286), .O(n10241));
  LUT5 #(.INIT(32'h96696996)) lut_n10242 (.I0(x1275), .I1(x1276), .I2(x1277), .I3(n10238), .I4(n10239), .O(n10242));
  LUT5 #(.INIT(32'hFF969600)) lut_n10243 (.I0(x1281), .I1(x1282), .I2(x1283), .I3(n10241), .I4(n10242), .O(n10243));
  LUT3 #(.INIT(8'h96)) lut_n10244 (.I0(n10224), .I1(n10227), .I2(n10228), .O(n10244));
  LUT3 #(.INIT(8'hE8)) lut_n10245 (.I0(n10240), .I1(n10243), .I2(n10244), .O(n10245));
  LUT3 #(.INIT(8'h96)) lut_n10246 (.I0(x1290), .I1(x1291), .I2(x1292), .O(n10246));
  LUT5 #(.INIT(32'h96696996)) lut_n10247 (.I0(x1281), .I1(x1282), .I2(x1283), .I3(n10241), .I4(n10242), .O(n10247));
  LUT5 #(.INIT(32'hFF969600)) lut_n10248 (.I0(x1287), .I1(x1288), .I2(x1289), .I3(n10246), .I4(n10247), .O(n10248));
  LUT3 #(.INIT(8'h96)) lut_n10249 (.I0(x1296), .I1(x1297), .I2(x1298), .O(n10249));
  LUT5 #(.INIT(32'h96696996)) lut_n10250 (.I0(x1287), .I1(x1288), .I2(x1289), .I3(n10246), .I4(n10247), .O(n10250));
  LUT5 #(.INIT(32'hFF969600)) lut_n10251 (.I0(x1293), .I1(x1294), .I2(x1295), .I3(n10249), .I4(n10250), .O(n10251));
  LUT3 #(.INIT(8'h96)) lut_n10252 (.I0(n10240), .I1(n10243), .I2(n10244), .O(n10252));
  LUT3 #(.INIT(8'hE8)) lut_n10253 (.I0(n10248), .I1(n10251), .I2(n10252), .O(n10253));
  LUT3 #(.INIT(8'h96)) lut_n10254 (.I0(n10221), .I1(n10229), .I2(n10230), .O(n10254));
  LUT3 #(.INIT(8'hE8)) lut_n10255 (.I0(n10245), .I1(n10253), .I2(n10254), .O(n10255));
  LUT3 #(.INIT(8'h96)) lut_n10256 (.I0(x1302), .I1(x1303), .I2(x1304), .O(n10256));
  LUT5 #(.INIT(32'h96696996)) lut_n10257 (.I0(x1293), .I1(x1294), .I2(x1295), .I3(n10249), .I4(n10250), .O(n10257));
  LUT5 #(.INIT(32'hFF969600)) lut_n10258 (.I0(x1299), .I1(x1300), .I2(x1301), .I3(n10256), .I4(n10257), .O(n10258));
  LUT3 #(.INIT(8'h96)) lut_n10259 (.I0(x1308), .I1(x1309), .I2(x1310), .O(n10259));
  LUT5 #(.INIT(32'h96696996)) lut_n10260 (.I0(x1299), .I1(x1300), .I2(x1301), .I3(n10256), .I4(n10257), .O(n10260));
  LUT5 #(.INIT(32'hFF969600)) lut_n10261 (.I0(x1305), .I1(x1306), .I2(x1307), .I3(n10259), .I4(n10260), .O(n10261));
  LUT3 #(.INIT(8'h96)) lut_n10262 (.I0(n10248), .I1(n10251), .I2(n10252), .O(n10262));
  LUT3 #(.INIT(8'hE8)) lut_n10263 (.I0(n10258), .I1(n10261), .I2(n10262), .O(n10263));
  LUT3 #(.INIT(8'h96)) lut_n10264 (.I0(x1314), .I1(x1315), .I2(x1316), .O(n10264));
  LUT5 #(.INIT(32'h96696996)) lut_n10265 (.I0(x1305), .I1(x1306), .I2(x1307), .I3(n10259), .I4(n10260), .O(n10265));
  LUT5 #(.INIT(32'hFF969600)) lut_n10266 (.I0(x1311), .I1(x1312), .I2(x1313), .I3(n10264), .I4(n10265), .O(n10266));
  LUT3 #(.INIT(8'h96)) lut_n10267 (.I0(x1320), .I1(x1321), .I2(x1322), .O(n10267));
  LUT5 #(.INIT(32'h96696996)) lut_n10268 (.I0(x1311), .I1(x1312), .I2(x1313), .I3(n10264), .I4(n10265), .O(n10268));
  LUT5 #(.INIT(32'hFF969600)) lut_n10269 (.I0(x1317), .I1(x1318), .I2(x1319), .I3(n10267), .I4(n10268), .O(n10269));
  LUT3 #(.INIT(8'h96)) lut_n10270 (.I0(n10258), .I1(n10261), .I2(n10262), .O(n10270));
  LUT3 #(.INIT(8'hE8)) lut_n10271 (.I0(n10266), .I1(n10269), .I2(n10270), .O(n10271));
  LUT3 #(.INIT(8'h96)) lut_n10272 (.I0(n10245), .I1(n10253), .I2(n10254), .O(n10272));
  LUT3 #(.INIT(8'hE8)) lut_n10273 (.I0(n10263), .I1(n10271), .I2(n10272), .O(n10273));
  LUT3 #(.INIT(8'h96)) lut_n10274 (.I0(n10213), .I1(n10231), .I2(n10232), .O(n10274));
  LUT3 #(.INIT(8'hE8)) lut_n10275 (.I0(n10255), .I1(n10273), .I2(n10274), .O(n10275));
  LUT3 #(.INIT(8'h96)) lut_n10276 (.I0(x1326), .I1(x1327), .I2(x1328), .O(n10276));
  LUT5 #(.INIT(32'h96696996)) lut_n10277 (.I0(x1317), .I1(x1318), .I2(x1319), .I3(n10267), .I4(n10268), .O(n10277));
  LUT5 #(.INIT(32'hFF969600)) lut_n10278 (.I0(x1323), .I1(x1324), .I2(x1325), .I3(n10276), .I4(n10277), .O(n10278));
  LUT3 #(.INIT(8'h96)) lut_n10279 (.I0(x1332), .I1(x1333), .I2(x1334), .O(n10279));
  LUT5 #(.INIT(32'h96696996)) lut_n10280 (.I0(x1323), .I1(x1324), .I2(x1325), .I3(n10276), .I4(n10277), .O(n10280));
  LUT5 #(.INIT(32'hFF969600)) lut_n10281 (.I0(x1329), .I1(x1330), .I2(x1331), .I3(n10279), .I4(n10280), .O(n10281));
  LUT3 #(.INIT(8'h96)) lut_n10282 (.I0(n10266), .I1(n10269), .I2(n10270), .O(n10282));
  LUT3 #(.INIT(8'hE8)) lut_n10283 (.I0(n10278), .I1(n10281), .I2(n10282), .O(n10283));
  LUT3 #(.INIT(8'h96)) lut_n10284 (.I0(x1338), .I1(x1339), .I2(x1340), .O(n10284));
  LUT5 #(.INIT(32'h96696996)) lut_n10285 (.I0(x1329), .I1(x1330), .I2(x1331), .I3(n10279), .I4(n10280), .O(n10285));
  LUT5 #(.INIT(32'hFF969600)) lut_n10286 (.I0(x1335), .I1(x1336), .I2(x1337), .I3(n10284), .I4(n10285), .O(n10286));
  LUT3 #(.INIT(8'h96)) lut_n10287 (.I0(x1344), .I1(x1345), .I2(x1346), .O(n10287));
  LUT5 #(.INIT(32'h96696996)) lut_n10288 (.I0(x1335), .I1(x1336), .I2(x1337), .I3(n10284), .I4(n10285), .O(n10288));
  LUT5 #(.INIT(32'hFF969600)) lut_n10289 (.I0(x1341), .I1(x1342), .I2(x1343), .I3(n10287), .I4(n10288), .O(n10289));
  LUT3 #(.INIT(8'h96)) lut_n10290 (.I0(n10278), .I1(n10281), .I2(n10282), .O(n10290));
  LUT3 #(.INIT(8'hE8)) lut_n10291 (.I0(n10286), .I1(n10289), .I2(n10290), .O(n10291));
  LUT3 #(.INIT(8'h96)) lut_n10292 (.I0(n10263), .I1(n10271), .I2(n10272), .O(n10292));
  LUT3 #(.INIT(8'hE8)) lut_n10293 (.I0(n10283), .I1(n10291), .I2(n10292), .O(n10293));
  LUT3 #(.INIT(8'h96)) lut_n10294 (.I0(x1350), .I1(x1351), .I2(x1352), .O(n10294));
  LUT5 #(.INIT(32'h96696996)) lut_n10295 (.I0(x1341), .I1(x1342), .I2(x1343), .I3(n10287), .I4(n10288), .O(n10295));
  LUT5 #(.INIT(32'hFF969600)) lut_n10296 (.I0(x1347), .I1(x1348), .I2(x1349), .I3(n10294), .I4(n10295), .O(n10296));
  LUT3 #(.INIT(8'h96)) lut_n10297 (.I0(x1356), .I1(x1357), .I2(x1358), .O(n10297));
  LUT5 #(.INIT(32'h96696996)) lut_n10298 (.I0(x1347), .I1(x1348), .I2(x1349), .I3(n10294), .I4(n10295), .O(n10298));
  LUT5 #(.INIT(32'hFF969600)) lut_n10299 (.I0(x1353), .I1(x1354), .I2(x1355), .I3(n10297), .I4(n10298), .O(n10299));
  LUT3 #(.INIT(8'h96)) lut_n10300 (.I0(n10286), .I1(n10289), .I2(n10290), .O(n10300));
  LUT3 #(.INIT(8'hE8)) lut_n10301 (.I0(n10296), .I1(n10299), .I2(n10300), .O(n10301));
  LUT3 #(.INIT(8'h96)) lut_n10302 (.I0(x1362), .I1(x1363), .I2(x1364), .O(n10302));
  LUT5 #(.INIT(32'h96696996)) lut_n10303 (.I0(x1353), .I1(x1354), .I2(x1355), .I3(n10297), .I4(n10298), .O(n10303));
  LUT5 #(.INIT(32'hFF969600)) lut_n10304 (.I0(x1359), .I1(x1360), .I2(x1361), .I3(n10302), .I4(n10303), .O(n10304));
  LUT3 #(.INIT(8'h96)) lut_n10305 (.I0(x1368), .I1(x1369), .I2(x1370), .O(n10305));
  LUT5 #(.INIT(32'h96696996)) lut_n10306 (.I0(x1359), .I1(x1360), .I2(x1361), .I3(n10302), .I4(n10303), .O(n10306));
  LUT5 #(.INIT(32'hFF969600)) lut_n10307 (.I0(x1365), .I1(x1366), .I2(x1367), .I3(n10305), .I4(n10306), .O(n10307));
  LUT3 #(.INIT(8'h96)) lut_n10308 (.I0(n10296), .I1(n10299), .I2(n10300), .O(n10308));
  LUT3 #(.INIT(8'hE8)) lut_n10309 (.I0(n10304), .I1(n10307), .I2(n10308), .O(n10309));
  LUT3 #(.INIT(8'h96)) lut_n10310 (.I0(n10283), .I1(n10291), .I2(n10292), .O(n10310));
  LUT3 #(.INIT(8'hE8)) lut_n10311 (.I0(n10301), .I1(n10309), .I2(n10310), .O(n10311));
  LUT3 #(.INIT(8'h96)) lut_n10312 (.I0(n10255), .I1(n10273), .I2(n10274), .O(n10312));
  LUT3 #(.INIT(8'hE8)) lut_n10313 (.I0(n10293), .I1(n10311), .I2(n10312), .O(n10313));
  LUT3 #(.INIT(8'h96)) lut_n10314 (.I0(n10195), .I1(n10233), .I2(n10234), .O(n10314));
  LUT3 #(.INIT(8'hE8)) lut_n10315 (.I0(n10275), .I1(n10313), .I2(n10314), .O(n10315));
  LUT3 #(.INIT(8'h96)) lut_n10316 (.I0(x1374), .I1(x1375), .I2(x1376), .O(n10316));
  LUT5 #(.INIT(32'h96696996)) lut_n10317 (.I0(x1365), .I1(x1366), .I2(x1367), .I3(n10305), .I4(n10306), .O(n10317));
  LUT5 #(.INIT(32'hFF969600)) lut_n10318 (.I0(x1371), .I1(x1372), .I2(x1373), .I3(n10316), .I4(n10317), .O(n10318));
  LUT3 #(.INIT(8'h96)) lut_n10319 (.I0(x1380), .I1(x1381), .I2(x1382), .O(n10319));
  LUT5 #(.INIT(32'h96696996)) lut_n10320 (.I0(x1371), .I1(x1372), .I2(x1373), .I3(n10316), .I4(n10317), .O(n10320));
  LUT5 #(.INIT(32'hFF969600)) lut_n10321 (.I0(x1377), .I1(x1378), .I2(x1379), .I3(n10319), .I4(n10320), .O(n10321));
  LUT3 #(.INIT(8'h96)) lut_n10322 (.I0(n10304), .I1(n10307), .I2(n10308), .O(n10322));
  LUT3 #(.INIT(8'hE8)) lut_n10323 (.I0(n10318), .I1(n10321), .I2(n10322), .O(n10323));
  LUT3 #(.INIT(8'h96)) lut_n10324 (.I0(x1386), .I1(x1387), .I2(x1388), .O(n10324));
  LUT5 #(.INIT(32'h96696996)) lut_n10325 (.I0(x1377), .I1(x1378), .I2(x1379), .I3(n10319), .I4(n10320), .O(n10325));
  LUT5 #(.INIT(32'hFF969600)) lut_n10326 (.I0(x1383), .I1(x1384), .I2(x1385), .I3(n10324), .I4(n10325), .O(n10326));
  LUT3 #(.INIT(8'h96)) lut_n10327 (.I0(x1392), .I1(x1393), .I2(x1394), .O(n10327));
  LUT5 #(.INIT(32'h96696996)) lut_n10328 (.I0(x1383), .I1(x1384), .I2(x1385), .I3(n10324), .I4(n10325), .O(n10328));
  LUT5 #(.INIT(32'hFF969600)) lut_n10329 (.I0(x1389), .I1(x1390), .I2(x1391), .I3(n10327), .I4(n10328), .O(n10329));
  LUT3 #(.INIT(8'h96)) lut_n10330 (.I0(n10318), .I1(n10321), .I2(n10322), .O(n10330));
  LUT3 #(.INIT(8'hE8)) lut_n10331 (.I0(n10326), .I1(n10329), .I2(n10330), .O(n10331));
  LUT3 #(.INIT(8'h96)) lut_n10332 (.I0(n10301), .I1(n10309), .I2(n10310), .O(n10332));
  LUT3 #(.INIT(8'hE8)) lut_n10333 (.I0(n10323), .I1(n10331), .I2(n10332), .O(n10333));
  LUT3 #(.INIT(8'h96)) lut_n10334 (.I0(x1398), .I1(x1399), .I2(x1400), .O(n10334));
  LUT5 #(.INIT(32'h96696996)) lut_n10335 (.I0(x1389), .I1(x1390), .I2(x1391), .I3(n10327), .I4(n10328), .O(n10335));
  LUT5 #(.INIT(32'hFF969600)) lut_n10336 (.I0(x1395), .I1(x1396), .I2(x1397), .I3(n10334), .I4(n10335), .O(n10336));
  LUT3 #(.INIT(8'h96)) lut_n10337 (.I0(x1404), .I1(x1405), .I2(x1406), .O(n10337));
  LUT5 #(.INIT(32'h96696996)) lut_n10338 (.I0(x1395), .I1(x1396), .I2(x1397), .I3(n10334), .I4(n10335), .O(n10338));
  LUT5 #(.INIT(32'hFF969600)) lut_n10339 (.I0(x1401), .I1(x1402), .I2(x1403), .I3(n10337), .I4(n10338), .O(n10339));
  LUT3 #(.INIT(8'h96)) lut_n10340 (.I0(n10326), .I1(n10329), .I2(n10330), .O(n10340));
  LUT3 #(.INIT(8'hE8)) lut_n10341 (.I0(n10336), .I1(n10339), .I2(n10340), .O(n10341));
  LUT3 #(.INIT(8'h96)) lut_n10342 (.I0(x1410), .I1(x1411), .I2(x1412), .O(n10342));
  LUT5 #(.INIT(32'h96696996)) lut_n10343 (.I0(x1401), .I1(x1402), .I2(x1403), .I3(n10337), .I4(n10338), .O(n10343));
  LUT5 #(.INIT(32'hFF969600)) lut_n10344 (.I0(x1407), .I1(x1408), .I2(x1409), .I3(n10342), .I4(n10343), .O(n10344));
  LUT3 #(.INIT(8'h96)) lut_n10345 (.I0(x1416), .I1(x1417), .I2(x1418), .O(n10345));
  LUT5 #(.INIT(32'h96696996)) lut_n10346 (.I0(x1407), .I1(x1408), .I2(x1409), .I3(n10342), .I4(n10343), .O(n10346));
  LUT5 #(.INIT(32'hFF969600)) lut_n10347 (.I0(x1413), .I1(x1414), .I2(x1415), .I3(n10345), .I4(n10346), .O(n10347));
  LUT3 #(.INIT(8'h96)) lut_n10348 (.I0(n10336), .I1(n10339), .I2(n10340), .O(n10348));
  LUT3 #(.INIT(8'hE8)) lut_n10349 (.I0(n10344), .I1(n10347), .I2(n10348), .O(n10349));
  LUT3 #(.INIT(8'h96)) lut_n10350 (.I0(n10323), .I1(n10331), .I2(n10332), .O(n10350));
  LUT3 #(.INIT(8'hE8)) lut_n10351 (.I0(n10341), .I1(n10349), .I2(n10350), .O(n10351));
  LUT3 #(.INIT(8'h96)) lut_n10352 (.I0(n10293), .I1(n10311), .I2(n10312), .O(n10352));
  LUT3 #(.INIT(8'hE8)) lut_n10353 (.I0(n10333), .I1(n10351), .I2(n10352), .O(n10353));
  LUT3 #(.INIT(8'h96)) lut_n10354 (.I0(x1422), .I1(x1423), .I2(x1424), .O(n10354));
  LUT5 #(.INIT(32'h96696996)) lut_n10355 (.I0(x1413), .I1(x1414), .I2(x1415), .I3(n10345), .I4(n10346), .O(n10355));
  LUT5 #(.INIT(32'hFF969600)) lut_n10356 (.I0(x1419), .I1(x1420), .I2(x1421), .I3(n10354), .I4(n10355), .O(n10356));
  LUT3 #(.INIT(8'h96)) lut_n10357 (.I0(x1428), .I1(x1429), .I2(x1430), .O(n10357));
  LUT5 #(.INIT(32'h96696996)) lut_n10358 (.I0(x1419), .I1(x1420), .I2(x1421), .I3(n10354), .I4(n10355), .O(n10358));
  LUT5 #(.INIT(32'hFF969600)) lut_n10359 (.I0(x1425), .I1(x1426), .I2(x1427), .I3(n10357), .I4(n10358), .O(n10359));
  LUT3 #(.INIT(8'h96)) lut_n10360 (.I0(n10344), .I1(n10347), .I2(n10348), .O(n10360));
  LUT3 #(.INIT(8'hE8)) lut_n10361 (.I0(n10356), .I1(n10359), .I2(n10360), .O(n10361));
  LUT3 #(.INIT(8'h96)) lut_n10362 (.I0(x1434), .I1(x1435), .I2(x1436), .O(n10362));
  LUT5 #(.INIT(32'h96696996)) lut_n10363 (.I0(x1425), .I1(x1426), .I2(x1427), .I3(n10357), .I4(n10358), .O(n10363));
  LUT5 #(.INIT(32'hFF969600)) lut_n10364 (.I0(x1431), .I1(x1432), .I2(x1433), .I3(n10362), .I4(n10363), .O(n10364));
  LUT3 #(.INIT(8'h96)) lut_n10365 (.I0(x1440), .I1(x1441), .I2(x1442), .O(n10365));
  LUT5 #(.INIT(32'h96696996)) lut_n10366 (.I0(x1431), .I1(x1432), .I2(x1433), .I3(n10362), .I4(n10363), .O(n10366));
  LUT5 #(.INIT(32'hFF969600)) lut_n10367 (.I0(x1437), .I1(x1438), .I2(x1439), .I3(n10365), .I4(n10366), .O(n10367));
  LUT3 #(.INIT(8'h96)) lut_n10368 (.I0(n10356), .I1(n10359), .I2(n10360), .O(n10368));
  LUT3 #(.INIT(8'hE8)) lut_n10369 (.I0(n10364), .I1(n10367), .I2(n10368), .O(n10369));
  LUT3 #(.INIT(8'h96)) lut_n10370 (.I0(n10341), .I1(n10349), .I2(n10350), .O(n10370));
  LUT3 #(.INIT(8'hE8)) lut_n10371 (.I0(n10361), .I1(n10369), .I2(n10370), .O(n10371));
  LUT3 #(.INIT(8'h96)) lut_n10372 (.I0(x1446), .I1(x1447), .I2(x1448), .O(n10372));
  LUT5 #(.INIT(32'h96696996)) lut_n10373 (.I0(x1437), .I1(x1438), .I2(x1439), .I3(n10365), .I4(n10366), .O(n10373));
  LUT5 #(.INIT(32'hFF969600)) lut_n10374 (.I0(x1443), .I1(x1444), .I2(x1445), .I3(n10372), .I4(n10373), .O(n10374));
  LUT3 #(.INIT(8'h96)) lut_n10375 (.I0(x1452), .I1(x1453), .I2(x1454), .O(n10375));
  LUT5 #(.INIT(32'h96696996)) lut_n10376 (.I0(x1443), .I1(x1444), .I2(x1445), .I3(n10372), .I4(n10373), .O(n10376));
  LUT5 #(.INIT(32'hFF969600)) lut_n10377 (.I0(x1449), .I1(x1450), .I2(x1451), .I3(n10375), .I4(n10376), .O(n10377));
  LUT3 #(.INIT(8'h96)) lut_n10378 (.I0(n10364), .I1(n10367), .I2(n10368), .O(n10378));
  LUT3 #(.INIT(8'hE8)) lut_n10379 (.I0(n10374), .I1(n10377), .I2(n10378), .O(n10379));
  LUT3 #(.INIT(8'h96)) lut_n10380 (.I0(x1458), .I1(x1459), .I2(x1460), .O(n10380));
  LUT5 #(.INIT(32'h96696996)) lut_n10381 (.I0(x1449), .I1(x1450), .I2(x1451), .I3(n10375), .I4(n10376), .O(n10381));
  LUT5 #(.INIT(32'hFF969600)) lut_n10382 (.I0(x1455), .I1(x1456), .I2(x1457), .I3(n10380), .I4(n10381), .O(n10382));
  LUT3 #(.INIT(8'h96)) lut_n10383 (.I0(x1464), .I1(x1465), .I2(x1466), .O(n10383));
  LUT5 #(.INIT(32'h96696996)) lut_n10384 (.I0(x1455), .I1(x1456), .I2(x1457), .I3(n10380), .I4(n10381), .O(n10384));
  LUT5 #(.INIT(32'hFF969600)) lut_n10385 (.I0(x1461), .I1(x1462), .I2(x1463), .I3(n10383), .I4(n10384), .O(n10385));
  LUT3 #(.INIT(8'h96)) lut_n10386 (.I0(n10374), .I1(n10377), .I2(n10378), .O(n10386));
  LUT3 #(.INIT(8'hE8)) lut_n10387 (.I0(n10382), .I1(n10385), .I2(n10386), .O(n10387));
  LUT3 #(.INIT(8'h96)) lut_n10388 (.I0(n10361), .I1(n10369), .I2(n10370), .O(n10388));
  LUT3 #(.INIT(8'hE8)) lut_n10389 (.I0(n10379), .I1(n10387), .I2(n10388), .O(n10389));
  LUT3 #(.INIT(8'h96)) lut_n10390 (.I0(n10333), .I1(n10351), .I2(n10352), .O(n10390));
  LUT3 #(.INIT(8'hE8)) lut_n10391 (.I0(n10371), .I1(n10389), .I2(n10390), .O(n10391));
  LUT3 #(.INIT(8'h96)) lut_n10392 (.I0(n10275), .I1(n10313), .I2(n10314), .O(n10392));
  LUT3 #(.INIT(8'hE8)) lut_n10393 (.I0(n10353), .I1(n10391), .I2(n10392), .O(n10393));
  LUT3 #(.INIT(8'h96)) lut_n10394 (.I0(n10157), .I1(n10235), .I2(n10236), .O(n10394));
  LUT3 #(.INIT(8'hE8)) lut_n10395 (.I0(n10315), .I1(n10393), .I2(n10394), .O(n10395));
  LUT3 #(.INIT(8'h96)) lut_n10396 (.I0(n9919), .I1(n10077), .I2(n10078), .O(n10396));
  LUT3 #(.INIT(8'hE8)) lut_n10397 (.I0(n10237), .I1(n10395), .I2(n10396), .O(n10397));
  LUT3 #(.INIT(8'h96)) lut_n10398 (.I0(n9439), .I1(n9757), .I2(n9758), .O(n10398));
  LUT3 #(.INIT(8'hE8)) lut_n10399 (.I0(n10079), .I1(n10397), .I2(n10398), .O(n10399));
  LUT3 #(.INIT(8'h96)) lut_n10400 (.I0(x1470), .I1(x1471), .I2(x1472), .O(n10400));
  LUT5 #(.INIT(32'h96696996)) lut_n10401 (.I0(x1461), .I1(x1462), .I2(x1463), .I3(n10383), .I4(n10384), .O(n10401));
  LUT5 #(.INIT(32'hFF969600)) lut_n10402 (.I0(x1467), .I1(x1468), .I2(x1469), .I3(n10400), .I4(n10401), .O(n10402));
  LUT3 #(.INIT(8'h96)) lut_n10403 (.I0(x1476), .I1(x1477), .I2(x1478), .O(n10403));
  LUT5 #(.INIT(32'h96696996)) lut_n10404 (.I0(x1467), .I1(x1468), .I2(x1469), .I3(n10400), .I4(n10401), .O(n10404));
  LUT5 #(.INIT(32'hFF969600)) lut_n10405 (.I0(x1473), .I1(x1474), .I2(x1475), .I3(n10403), .I4(n10404), .O(n10405));
  LUT3 #(.INIT(8'h96)) lut_n10406 (.I0(n10382), .I1(n10385), .I2(n10386), .O(n10406));
  LUT3 #(.INIT(8'hE8)) lut_n10407 (.I0(n10402), .I1(n10405), .I2(n10406), .O(n10407));
  LUT3 #(.INIT(8'h96)) lut_n10408 (.I0(x1482), .I1(x1483), .I2(x1484), .O(n10408));
  LUT5 #(.INIT(32'h96696996)) lut_n10409 (.I0(x1473), .I1(x1474), .I2(x1475), .I3(n10403), .I4(n10404), .O(n10409));
  LUT5 #(.INIT(32'hFF969600)) lut_n10410 (.I0(x1479), .I1(x1480), .I2(x1481), .I3(n10408), .I4(n10409), .O(n10410));
  LUT3 #(.INIT(8'h96)) lut_n10411 (.I0(x1488), .I1(x1489), .I2(x1490), .O(n10411));
  LUT5 #(.INIT(32'h96696996)) lut_n10412 (.I0(x1479), .I1(x1480), .I2(x1481), .I3(n10408), .I4(n10409), .O(n10412));
  LUT5 #(.INIT(32'hFF969600)) lut_n10413 (.I0(x1485), .I1(x1486), .I2(x1487), .I3(n10411), .I4(n10412), .O(n10413));
  LUT3 #(.INIT(8'h96)) lut_n10414 (.I0(n10402), .I1(n10405), .I2(n10406), .O(n10414));
  LUT3 #(.INIT(8'hE8)) lut_n10415 (.I0(n10410), .I1(n10413), .I2(n10414), .O(n10415));
  LUT3 #(.INIT(8'h96)) lut_n10416 (.I0(n10379), .I1(n10387), .I2(n10388), .O(n10416));
  LUT3 #(.INIT(8'hE8)) lut_n10417 (.I0(n10407), .I1(n10415), .I2(n10416), .O(n10417));
  LUT3 #(.INIT(8'h96)) lut_n10418 (.I0(x1494), .I1(x1495), .I2(x1496), .O(n10418));
  LUT5 #(.INIT(32'h96696996)) lut_n10419 (.I0(x1485), .I1(x1486), .I2(x1487), .I3(n10411), .I4(n10412), .O(n10419));
  LUT5 #(.INIT(32'hFF969600)) lut_n10420 (.I0(x1491), .I1(x1492), .I2(x1493), .I3(n10418), .I4(n10419), .O(n10420));
  LUT3 #(.INIT(8'h96)) lut_n10421 (.I0(x1500), .I1(x1501), .I2(x1502), .O(n10421));
  LUT5 #(.INIT(32'h96696996)) lut_n10422 (.I0(x1491), .I1(x1492), .I2(x1493), .I3(n10418), .I4(n10419), .O(n10422));
  LUT5 #(.INIT(32'hFF969600)) lut_n10423 (.I0(x1497), .I1(x1498), .I2(x1499), .I3(n10421), .I4(n10422), .O(n10423));
  LUT3 #(.INIT(8'h96)) lut_n10424 (.I0(n10410), .I1(n10413), .I2(n10414), .O(n10424));
  LUT3 #(.INIT(8'hE8)) lut_n10425 (.I0(n10420), .I1(n10423), .I2(n10424), .O(n10425));
  LUT3 #(.INIT(8'h96)) lut_n10426 (.I0(x1506), .I1(x1507), .I2(x1508), .O(n10426));
  LUT5 #(.INIT(32'h96696996)) lut_n10427 (.I0(x1497), .I1(x1498), .I2(x1499), .I3(n10421), .I4(n10422), .O(n10427));
  LUT5 #(.INIT(32'hFF969600)) lut_n10428 (.I0(x1503), .I1(x1504), .I2(x1505), .I3(n10426), .I4(n10427), .O(n10428));
  LUT3 #(.INIT(8'h96)) lut_n10429 (.I0(x1512), .I1(x1513), .I2(x1514), .O(n10429));
  LUT5 #(.INIT(32'h96696996)) lut_n10430 (.I0(x1503), .I1(x1504), .I2(x1505), .I3(n10426), .I4(n10427), .O(n10430));
  LUT5 #(.INIT(32'hFF969600)) lut_n10431 (.I0(x1509), .I1(x1510), .I2(x1511), .I3(n10429), .I4(n10430), .O(n10431));
  LUT3 #(.INIT(8'h96)) lut_n10432 (.I0(n10420), .I1(n10423), .I2(n10424), .O(n10432));
  LUT3 #(.INIT(8'hE8)) lut_n10433 (.I0(n10428), .I1(n10431), .I2(n10432), .O(n10433));
  LUT3 #(.INIT(8'h96)) lut_n10434 (.I0(n10407), .I1(n10415), .I2(n10416), .O(n10434));
  LUT3 #(.INIT(8'hE8)) lut_n10435 (.I0(n10425), .I1(n10433), .I2(n10434), .O(n10435));
  LUT3 #(.INIT(8'h96)) lut_n10436 (.I0(n10371), .I1(n10389), .I2(n10390), .O(n10436));
  LUT3 #(.INIT(8'hE8)) lut_n10437 (.I0(n10417), .I1(n10435), .I2(n10436), .O(n10437));
  LUT3 #(.INIT(8'h96)) lut_n10438 (.I0(x1518), .I1(x1519), .I2(x1520), .O(n10438));
  LUT5 #(.INIT(32'h96696996)) lut_n10439 (.I0(x1509), .I1(x1510), .I2(x1511), .I3(n10429), .I4(n10430), .O(n10439));
  LUT5 #(.INIT(32'hFF969600)) lut_n10440 (.I0(x1515), .I1(x1516), .I2(x1517), .I3(n10438), .I4(n10439), .O(n10440));
  LUT3 #(.INIT(8'h96)) lut_n10441 (.I0(x1524), .I1(x1525), .I2(x1526), .O(n10441));
  LUT5 #(.INIT(32'h96696996)) lut_n10442 (.I0(x1515), .I1(x1516), .I2(x1517), .I3(n10438), .I4(n10439), .O(n10442));
  LUT5 #(.INIT(32'hFF969600)) lut_n10443 (.I0(x1521), .I1(x1522), .I2(x1523), .I3(n10441), .I4(n10442), .O(n10443));
  LUT3 #(.INIT(8'h96)) lut_n10444 (.I0(n10428), .I1(n10431), .I2(n10432), .O(n10444));
  LUT3 #(.INIT(8'hE8)) lut_n10445 (.I0(n10440), .I1(n10443), .I2(n10444), .O(n10445));
  LUT3 #(.INIT(8'h96)) lut_n10446 (.I0(x1530), .I1(x1531), .I2(x1532), .O(n10446));
  LUT5 #(.INIT(32'h96696996)) lut_n10447 (.I0(x1521), .I1(x1522), .I2(x1523), .I3(n10441), .I4(n10442), .O(n10447));
  LUT5 #(.INIT(32'hFF969600)) lut_n10448 (.I0(x1527), .I1(x1528), .I2(x1529), .I3(n10446), .I4(n10447), .O(n10448));
  LUT3 #(.INIT(8'h96)) lut_n10449 (.I0(x1536), .I1(x1537), .I2(x1538), .O(n10449));
  LUT5 #(.INIT(32'h96696996)) lut_n10450 (.I0(x1527), .I1(x1528), .I2(x1529), .I3(n10446), .I4(n10447), .O(n10450));
  LUT5 #(.INIT(32'hFF969600)) lut_n10451 (.I0(x1533), .I1(x1534), .I2(x1535), .I3(n10449), .I4(n10450), .O(n10451));
  LUT3 #(.INIT(8'h96)) lut_n10452 (.I0(n10440), .I1(n10443), .I2(n10444), .O(n10452));
  LUT3 #(.INIT(8'hE8)) lut_n10453 (.I0(n10448), .I1(n10451), .I2(n10452), .O(n10453));
  LUT3 #(.INIT(8'h96)) lut_n10454 (.I0(n10425), .I1(n10433), .I2(n10434), .O(n10454));
  LUT3 #(.INIT(8'hE8)) lut_n10455 (.I0(n10445), .I1(n10453), .I2(n10454), .O(n10455));
  LUT3 #(.INIT(8'h96)) lut_n10456 (.I0(x1542), .I1(x1543), .I2(x1544), .O(n10456));
  LUT5 #(.INIT(32'h96696996)) lut_n10457 (.I0(x1533), .I1(x1534), .I2(x1535), .I3(n10449), .I4(n10450), .O(n10457));
  LUT5 #(.INIT(32'hFF969600)) lut_n10458 (.I0(x1539), .I1(x1540), .I2(x1541), .I3(n10456), .I4(n10457), .O(n10458));
  LUT3 #(.INIT(8'h96)) lut_n10459 (.I0(x1548), .I1(x1549), .I2(x1550), .O(n10459));
  LUT5 #(.INIT(32'h96696996)) lut_n10460 (.I0(x1539), .I1(x1540), .I2(x1541), .I3(n10456), .I4(n10457), .O(n10460));
  LUT5 #(.INIT(32'hFF969600)) lut_n10461 (.I0(x1545), .I1(x1546), .I2(x1547), .I3(n10459), .I4(n10460), .O(n10461));
  LUT3 #(.INIT(8'h96)) lut_n10462 (.I0(n10448), .I1(n10451), .I2(n10452), .O(n10462));
  LUT3 #(.INIT(8'hE8)) lut_n10463 (.I0(n10458), .I1(n10461), .I2(n10462), .O(n10463));
  LUT3 #(.INIT(8'h96)) lut_n10464 (.I0(x1554), .I1(x1555), .I2(x1556), .O(n10464));
  LUT5 #(.INIT(32'h96696996)) lut_n10465 (.I0(x1545), .I1(x1546), .I2(x1547), .I3(n10459), .I4(n10460), .O(n10465));
  LUT5 #(.INIT(32'hFF969600)) lut_n10466 (.I0(x1551), .I1(x1552), .I2(x1553), .I3(n10464), .I4(n10465), .O(n10466));
  LUT3 #(.INIT(8'h96)) lut_n10467 (.I0(x1560), .I1(x1561), .I2(x1562), .O(n10467));
  LUT5 #(.INIT(32'h96696996)) lut_n10468 (.I0(x1551), .I1(x1552), .I2(x1553), .I3(n10464), .I4(n10465), .O(n10468));
  LUT5 #(.INIT(32'hFF969600)) lut_n10469 (.I0(x1557), .I1(x1558), .I2(x1559), .I3(n10467), .I4(n10468), .O(n10469));
  LUT3 #(.INIT(8'h96)) lut_n10470 (.I0(n10458), .I1(n10461), .I2(n10462), .O(n10470));
  LUT3 #(.INIT(8'hE8)) lut_n10471 (.I0(n10466), .I1(n10469), .I2(n10470), .O(n10471));
  LUT3 #(.INIT(8'h96)) lut_n10472 (.I0(n10445), .I1(n10453), .I2(n10454), .O(n10472));
  LUT3 #(.INIT(8'hE8)) lut_n10473 (.I0(n10463), .I1(n10471), .I2(n10472), .O(n10473));
  LUT3 #(.INIT(8'h96)) lut_n10474 (.I0(n10417), .I1(n10435), .I2(n10436), .O(n10474));
  LUT3 #(.INIT(8'hE8)) lut_n10475 (.I0(n10455), .I1(n10473), .I2(n10474), .O(n10475));
  LUT3 #(.INIT(8'h96)) lut_n10476 (.I0(n10353), .I1(n10391), .I2(n10392), .O(n10476));
  LUT3 #(.INIT(8'hE8)) lut_n10477 (.I0(n10437), .I1(n10475), .I2(n10476), .O(n10477));
  LUT3 #(.INIT(8'h96)) lut_n10478 (.I0(x1566), .I1(x1567), .I2(x1568), .O(n10478));
  LUT5 #(.INIT(32'h96696996)) lut_n10479 (.I0(x1557), .I1(x1558), .I2(x1559), .I3(n10467), .I4(n10468), .O(n10479));
  LUT5 #(.INIT(32'hFF969600)) lut_n10480 (.I0(x1563), .I1(x1564), .I2(x1565), .I3(n10478), .I4(n10479), .O(n10480));
  LUT3 #(.INIT(8'h96)) lut_n10481 (.I0(x1572), .I1(x1573), .I2(x1574), .O(n10481));
  LUT5 #(.INIT(32'h96696996)) lut_n10482 (.I0(x1563), .I1(x1564), .I2(x1565), .I3(n10478), .I4(n10479), .O(n10482));
  LUT5 #(.INIT(32'hFF969600)) lut_n10483 (.I0(x1569), .I1(x1570), .I2(x1571), .I3(n10481), .I4(n10482), .O(n10483));
  LUT3 #(.INIT(8'h96)) lut_n10484 (.I0(n10466), .I1(n10469), .I2(n10470), .O(n10484));
  LUT3 #(.INIT(8'hE8)) lut_n10485 (.I0(n10480), .I1(n10483), .I2(n10484), .O(n10485));
  LUT3 #(.INIT(8'h96)) lut_n10486 (.I0(x1578), .I1(x1579), .I2(x1580), .O(n10486));
  LUT5 #(.INIT(32'h96696996)) lut_n10487 (.I0(x1569), .I1(x1570), .I2(x1571), .I3(n10481), .I4(n10482), .O(n10487));
  LUT5 #(.INIT(32'hFF969600)) lut_n10488 (.I0(x1575), .I1(x1576), .I2(x1577), .I3(n10486), .I4(n10487), .O(n10488));
  LUT3 #(.INIT(8'h96)) lut_n10489 (.I0(x1584), .I1(x1585), .I2(x1586), .O(n10489));
  LUT5 #(.INIT(32'h96696996)) lut_n10490 (.I0(x1575), .I1(x1576), .I2(x1577), .I3(n10486), .I4(n10487), .O(n10490));
  LUT5 #(.INIT(32'hFF969600)) lut_n10491 (.I0(x1581), .I1(x1582), .I2(x1583), .I3(n10489), .I4(n10490), .O(n10491));
  LUT3 #(.INIT(8'h96)) lut_n10492 (.I0(n10480), .I1(n10483), .I2(n10484), .O(n10492));
  LUT3 #(.INIT(8'hE8)) lut_n10493 (.I0(n10488), .I1(n10491), .I2(n10492), .O(n10493));
  LUT3 #(.INIT(8'h96)) lut_n10494 (.I0(n10463), .I1(n10471), .I2(n10472), .O(n10494));
  LUT3 #(.INIT(8'hE8)) lut_n10495 (.I0(n10485), .I1(n10493), .I2(n10494), .O(n10495));
  LUT3 #(.INIT(8'h96)) lut_n10496 (.I0(x1590), .I1(x1591), .I2(x1592), .O(n10496));
  LUT5 #(.INIT(32'h96696996)) lut_n10497 (.I0(x1581), .I1(x1582), .I2(x1583), .I3(n10489), .I4(n10490), .O(n10497));
  LUT5 #(.INIT(32'hFF969600)) lut_n10498 (.I0(x1587), .I1(x1588), .I2(x1589), .I3(n10496), .I4(n10497), .O(n10498));
  LUT3 #(.INIT(8'h96)) lut_n10499 (.I0(x1596), .I1(x1597), .I2(x1598), .O(n10499));
  LUT5 #(.INIT(32'h96696996)) lut_n10500 (.I0(x1587), .I1(x1588), .I2(x1589), .I3(n10496), .I4(n10497), .O(n10500));
  LUT5 #(.INIT(32'hFF969600)) lut_n10501 (.I0(x1593), .I1(x1594), .I2(x1595), .I3(n10499), .I4(n10500), .O(n10501));
  LUT3 #(.INIT(8'h96)) lut_n10502 (.I0(n10488), .I1(n10491), .I2(n10492), .O(n10502));
  LUT3 #(.INIT(8'hE8)) lut_n10503 (.I0(n10498), .I1(n10501), .I2(n10502), .O(n10503));
  LUT3 #(.INIT(8'h96)) lut_n10504 (.I0(x1602), .I1(x1603), .I2(x1604), .O(n10504));
  LUT5 #(.INIT(32'h96696996)) lut_n10505 (.I0(x1593), .I1(x1594), .I2(x1595), .I3(n10499), .I4(n10500), .O(n10505));
  LUT5 #(.INIT(32'hFF969600)) lut_n10506 (.I0(x1599), .I1(x1600), .I2(x1601), .I3(n10504), .I4(n10505), .O(n10506));
  LUT3 #(.INIT(8'h96)) lut_n10507 (.I0(x1608), .I1(x1609), .I2(x1610), .O(n10507));
  LUT5 #(.INIT(32'h96696996)) lut_n10508 (.I0(x1599), .I1(x1600), .I2(x1601), .I3(n10504), .I4(n10505), .O(n10508));
  LUT5 #(.INIT(32'hFF969600)) lut_n10509 (.I0(x1605), .I1(x1606), .I2(x1607), .I3(n10507), .I4(n10508), .O(n10509));
  LUT3 #(.INIT(8'h96)) lut_n10510 (.I0(n10498), .I1(n10501), .I2(n10502), .O(n10510));
  LUT3 #(.INIT(8'hE8)) lut_n10511 (.I0(n10506), .I1(n10509), .I2(n10510), .O(n10511));
  LUT3 #(.INIT(8'h96)) lut_n10512 (.I0(n10485), .I1(n10493), .I2(n10494), .O(n10512));
  LUT3 #(.INIT(8'hE8)) lut_n10513 (.I0(n10503), .I1(n10511), .I2(n10512), .O(n10513));
  LUT3 #(.INIT(8'h96)) lut_n10514 (.I0(n10455), .I1(n10473), .I2(n10474), .O(n10514));
  LUT3 #(.INIT(8'hE8)) lut_n10515 (.I0(n10495), .I1(n10513), .I2(n10514), .O(n10515));
  LUT3 #(.INIT(8'h96)) lut_n10516 (.I0(x1614), .I1(x1615), .I2(x1616), .O(n10516));
  LUT5 #(.INIT(32'h96696996)) lut_n10517 (.I0(x1605), .I1(x1606), .I2(x1607), .I3(n10507), .I4(n10508), .O(n10517));
  LUT5 #(.INIT(32'hFF969600)) lut_n10518 (.I0(x1611), .I1(x1612), .I2(x1613), .I3(n10516), .I4(n10517), .O(n10518));
  LUT3 #(.INIT(8'h96)) lut_n10519 (.I0(x1620), .I1(x1621), .I2(x1622), .O(n10519));
  LUT5 #(.INIT(32'h96696996)) lut_n10520 (.I0(x1611), .I1(x1612), .I2(x1613), .I3(n10516), .I4(n10517), .O(n10520));
  LUT5 #(.INIT(32'hFF969600)) lut_n10521 (.I0(x1617), .I1(x1618), .I2(x1619), .I3(n10519), .I4(n10520), .O(n10521));
  LUT3 #(.INIT(8'h96)) lut_n10522 (.I0(n10506), .I1(n10509), .I2(n10510), .O(n10522));
  LUT3 #(.INIT(8'hE8)) lut_n10523 (.I0(n10518), .I1(n10521), .I2(n10522), .O(n10523));
  LUT3 #(.INIT(8'h96)) lut_n10524 (.I0(x1626), .I1(x1627), .I2(x1628), .O(n10524));
  LUT5 #(.INIT(32'h96696996)) lut_n10525 (.I0(x1617), .I1(x1618), .I2(x1619), .I3(n10519), .I4(n10520), .O(n10525));
  LUT5 #(.INIT(32'hFF969600)) lut_n10526 (.I0(x1623), .I1(x1624), .I2(x1625), .I3(n10524), .I4(n10525), .O(n10526));
  LUT3 #(.INIT(8'h96)) lut_n10527 (.I0(x1632), .I1(x1633), .I2(x1634), .O(n10527));
  LUT5 #(.INIT(32'h96696996)) lut_n10528 (.I0(x1623), .I1(x1624), .I2(x1625), .I3(n10524), .I4(n10525), .O(n10528));
  LUT5 #(.INIT(32'hFF969600)) lut_n10529 (.I0(x1629), .I1(x1630), .I2(x1631), .I3(n10527), .I4(n10528), .O(n10529));
  LUT3 #(.INIT(8'h96)) lut_n10530 (.I0(n10518), .I1(n10521), .I2(n10522), .O(n10530));
  LUT3 #(.INIT(8'hE8)) lut_n10531 (.I0(n10526), .I1(n10529), .I2(n10530), .O(n10531));
  LUT3 #(.INIT(8'h96)) lut_n10532 (.I0(n10503), .I1(n10511), .I2(n10512), .O(n10532));
  LUT3 #(.INIT(8'hE8)) lut_n10533 (.I0(n10523), .I1(n10531), .I2(n10532), .O(n10533));
  LUT3 #(.INIT(8'h96)) lut_n10534 (.I0(x1638), .I1(x1639), .I2(x1640), .O(n10534));
  LUT5 #(.INIT(32'h96696996)) lut_n10535 (.I0(x1629), .I1(x1630), .I2(x1631), .I3(n10527), .I4(n10528), .O(n10535));
  LUT5 #(.INIT(32'hFF969600)) lut_n10536 (.I0(x1635), .I1(x1636), .I2(x1637), .I3(n10534), .I4(n10535), .O(n10536));
  LUT3 #(.INIT(8'h96)) lut_n10537 (.I0(x1644), .I1(x1645), .I2(x1646), .O(n10537));
  LUT5 #(.INIT(32'h96696996)) lut_n10538 (.I0(x1635), .I1(x1636), .I2(x1637), .I3(n10534), .I4(n10535), .O(n10538));
  LUT5 #(.INIT(32'hFF969600)) lut_n10539 (.I0(x1641), .I1(x1642), .I2(x1643), .I3(n10537), .I4(n10538), .O(n10539));
  LUT3 #(.INIT(8'h96)) lut_n10540 (.I0(n10526), .I1(n10529), .I2(n10530), .O(n10540));
  LUT3 #(.INIT(8'hE8)) lut_n10541 (.I0(n10536), .I1(n10539), .I2(n10540), .O(n10541));
  LUT3 #(.INIT(8'h96)) lut_n10542 (.I0(x1650), .I1(x1651), .I2(x1652), .O(n10542));
  LUT5 #(.INIT(32'h96696996)) lut_n10543 (.I0(x1641), .I1(x1642), .I2(x1643), .I3(n10537), .I4(n10538), .O(n10543));
  LUT5 #(.INIT(32'hFF969600)) lut_n10544 (.I0(x1647), .I1(x1648), .I2(x1649), .I3(n10542), .I4(n10543), .O(n10544));
  LUT3 #(.INIT(8'h96)) lut_n10545 (.I0(x1656), .I1(x1657), .I2(x1658), .O(n10545));
  LUT5 #(.INIT(32'h96696996)) lut_n10546 (.I0(x1647), .I1(x1648), .I2(x1649), .I3(n10542), .I4(n10543), .O(n10546));
  LUT5 #(.INIT(32'hFF969600)) lut_n10547 (.I0(x1653), .I1(x1654), .I2(x1655), .I3(n10545), .I4(n10546), .O(n10547));
  LUT3 #(.INIT(8'h96)) lut_n10548 (.I0(n10536), .I1(n10539), .I2(n10540), .O(n10548));
  LUT3 #(.INIT(8'hE8)) lut_n10549 (.I0(n10544), .I1(n10547), .I2(n10548), .O(n10549));
  LUT3 #(.INIT(8'h96)) lut_n10550 (.I0(n10523), .I1(n10531), .I2(n10532), .O(n10550));
  LUT3 #(.INIT(8'hE8)) lut_n10551 (.I0(n10541), .I1(n10549), .I2(n10550), .O(n10551));
  LUT3 #(.INIT(8'h96)) lut_n10552 (.I0(n10495), .I1(n10513), .I2(n10514), .O(n10552));
  LUT3 #(.INIT(8'hE8)) lut_n10553 (.I0(n10533), .I1(n10551), .I2(n10552), .O(n10553));
  LUT3 #(.INIT(8'h96)) lut_n10554 (.I0(n10437), .I1(n10475), .I2(n10476), .O(n10554));
  LUT3 #(.INIT(8'hE8)) lut_n10555 (.I0(n10515), .I1(n10553), .I2(n10554), .O(n10555));
  LUT3 #(.INIT(8'h96)) lut_n10556 (.I0(n10315), .I1(n10393), .I2(n10394), .O(n10556));
  LUT3 #(.INIT(8'hE8)) lut_n10557 (.I0(n10477), .I1(n10555), .I2(n10556), .O(n10557));
  LUT3 #(.INIT(8'h96)) lut_n10558 (.I0(x1662), .I1(x1663), .I2(x1664), .O(n10558));
  LUT5 #(.INIT(32'h96696996)) lut_n10559 (.I0(x1653), .I1(x1654), .I2(x1655), .I3(n10545), .I4(n10546), .O(n10559));
  LUT5 #(.INIT(32'hFF969600)) lut_n10560 (.I0(x1659), .I1(x1660), .I2(x1661), .I3(n10558), .I4(n10559), .O(n10560));
  LUT3 #(.INIT(8'h96)) lut_n10561 (.I0(x1668), .I1(x1669), .I2(x1670), .O(n10561));
  LUT5 #(.INIT(32'h96696996)) lut_n10562 (.I0(x1659), .I1(x1660), .I2(x1661), .I3(n10558), .I4(n10559), .O(n10562));
  LUT5 #(.INIT(32'hFF969600)) lut_n10563 (.I0(x1665), .I1(x1666), .I2(x1667), .I3(n10561), .I4(n10562), .O(n10563));
  LUT3 #(.INIT(8'h96)) lut_n10564 (.I0(n10544), .I1(n10547), .I2(n10548), .O(n10564));
  LUT3 #(.INIT(8'hE8)) lut_n10565 (.I0(n10560), .I1(n10563), .I2(n10564), .O(n10565));
  LUT3 #(.INIT(8'h96)) lut_n10566 (.I0(x1674), .I1(x1675), .I2(x1676), .O(n10566));
  LUT5 #(.INIT(32'h96696996)) lut_n10567 (.I0(x1665), .I1(x1666), .I2(x1667), .I3(n10561), .I4(n10562), .O(n10567));
  LUT5 #(.INIT(32'hFF969600)) lut_n10568 (.I0(x1671), .I1(x1672), .I2(x1673), .I3(n10566), .I4(n10567), .O(n10568));
  LUT3 #(.INIT(8'h96)) lut_n10569 (.I0(x1680), .I1(x1681), .I2(x1682), .O(n10569));
  LUT5 #(.INIT(32'h96696996)) lut_n10570 (.I0(x1671), .I1(x1672), .I2(x1673), .I3(n10566), .I4(n10567), .O(n10570));
  LUT5 #(.INIT(32'hFF969600)) lut_n10571 (.I0(x1677), .I1(x1678), .I2(x1679), .I3(n10569), .I4(n10570), .O(n10571));
  LUT3 #(.INIT(8'h96)) lut_n10572 (.I0(n10560), .I1(n10563), .I2(n10564), .O(n10572));
  LUT3 #(.INIT(8'hE8)) lut_n10573 (.I0(n10568), .I1(n10571), .I2(n10572), .O(n10573));
  LUT3 #(.INIT(8'h96)) lut_n10574 (.I0(n10541), .I1(n10549), .I2(n10550), .O(n10574));
  LUT3 #(.INIT(8'hE8)) lut_n10575 (.I0(n10565), .I1(n10573), .I2(n10574), .O(n10575));
  LUT3 #(.INIT(8'h96)) lut_n10576 (.I0(x1686), .I1(x1687), .I2(x1688), .O(n10576));
  LUT5 #(.INIT(32'h96696996)) lut_n10577 (.I0(x1677), .I1(x1678), .I2(x1679), .I3(n10569), .I4(n10570), .O(n10577));
  LUT5 #(.INIT(32'hFF969600)) lut_n10578 (.I0(x1683), .I1(x1684), .I2(x1685), .I3(n10576), .I4(n10577), .O(n10578));
  LUT3 #(.INIT(8'h96)) lut_n10579 (.I0(x1692), .I1(x1693), .I2(x1694), .O(n10579));
  LUT5 #(.INIT(32'h96696996)) lut_n10580 (.I0(x1683), .I1(x1684), .I2(x1685), .I3(n10576), .I4(n10577), .O(n10580));
  LUT5 #(.INIT(32'hFF969600)) lut_n10581 (.I0(x1689), .I1(x1690), .I2(x1691), .I3(n10579), .I4(n10580), .O(n10581));
  LUT3 #(.INIT(8'h96)) lut_n10582 (.I0(n10568), .I1(n10571), .I2(n10572), .O(n10582));
  LUT3 #(.INIT(8'hE8)) lut_n10583 (.I0(n10578), .I1(n10581), .I2(n10582), .O(n10583));
  LUT3 #(.INIT(8'h96)) lut_n10584 (.I0(x1698), .I1(x1699), .I2(x1700), .O(n10584));
  LUT5 #(.INIT(32'h96696996)) lut_n10585 (.I0(x1689), .I1(x1690), .I2(x1691), .I3(n10579), .I4(n10580), .O(n10585));
  LUT5 #(.INIT(32'hFF969600)) lut_n10586 (.I0(x1695), .I1(x1696), .I2(x1697), .I3(n10584), .I4(n10585), .O(n10586));
  LUT3 #(.INIT(8'h96)) lut_n10587 (.I0(x1704), .I1(x1705), .I2(x1706), .O(n10587));
  LUT5 #(.INIT(32'h96696996)) lut_n10588 (.I0(x1695), .I1(x1696), .I2(x1697), .I3(n10584), .I4(n10585), .O(n10588));
  LUT5 #(.INIT(32'hFF969600)) lut_n10589 (.I0(x1701), .I1(x1702), .I2(x1703), .I3(n10587), .I4(n10588), .O(n10589));
  LUT3 #(.INIT(8'h96)) lut_n10590 (.I0(n10578), .I1(n10581), .I2(n10582), .O(n10590));
  LUT3 #(.INIT(8'hE8)) lut_n10591 (.I0(n10586), .I1(n10589), .I2(n10590), .O(n10591));
  LUT3 #(.INIT(8'h96)) lut_n10592 (.I0(n10565), .I1(n10573), .I2(n10574), .O(n10592));
  LUT3 #(.INIT(8'hE8)) lut_n10593 (.I0(n10583), .I1(n10591), .I2(n10592), .O(n10593));
  LUT3 #(.INIT(8'h96)) lut_n10594 (.I0(n10533), .I1(n10551), .I2(n10552), .O(n10594));
  LUT3 #(.INIT(8'hE8)) lut_n10595 (.I0(n10575), .I1(n10593), .I2(n10594), .O(n10595));
  LUT3 #(.INIT(8'h96)) lut_n10596 (.I0(x1710), .I1(x1711), .I2(x1712), .O(n10596));
  LUT5 #(.INIT(32'h96696996)) lut_n10597 (.I0(x1701), .I1(x1702), .I2(x1703), .I3(n10587), .I4(n10588), .O(n10597));
  LUT5 #(.INIT(32'hFF969600)) lut_n10598 (.I0(x1707), .I1(x1708), .I2(x1709), .I3(n10596), .I4(n10597), .O(n10598));
  LUT3 #(.INIT(8'h96)) lut_n10599 (.I0(x1716), .I1(x1717), .I2(x1718), .O(n10599));
  LUT5 #(.INIT(32'h96696996)) lut_n10600 (.I0(x1707), .I1(x1708), .I2(x1709), .I3(n10596), .I4(n10597), .O(n10600));
  LUT5 #(.INIT(32'hFF969600)) lut_n10601 (.I0(x1713), .I1(x1714), .I2(x1715), .I3(n10599), .I4(n10600), .O(n10601));
  LUT3 #(.INIT(8'h96)) lut_n10602 (.I0(n10586), .I1(n10589), .I2(n10590), .O(n10602));
  LUT3 #(.INIT(8'hE8)) lut_n10603 (.I0(n10598), .I1(n10601), .I2(n10602), .O(n10603));
  LUT3 #(.INIT(8'h96)) lut_n10604 (.I0(x1722), .I1(x1723), .I2(x1724), .O(n10604));
  LUT5 #(.INIT(32'h96696996)) lut_n10605 (.I0(x1713), .I1(x1714), .I2(x1715), .I3(n10599), .I4(n10600), .O(n10605));
  LUT5 #(.INIT(32'hFF969600)) lut_n10606 (.I0(x1719), .I1(x1720), .I2(x1721), .I3(n10604), .I4(n10605), .O(n10606));
  LUT3 #(.INIT(8'h96)) lut_n10607 (.I0(x1728), .I1(x1729), .I2(x1730), .O(n10607));
  LUT5 #(.INIT(32'h96696996)) lut_n10608 (.I0(x1719), .I1(x1720), .I2(x1721), .I3(n10604), .I4(n10605), .O(n10608));
  LUT5 #(.INIT(32'hFF969600)) lut_n10609 (.I0(x1725), .I1(x1726), .I2(x1727), .I3(n10607), .I4(n10608), .O(n10609));
  LUT3 #(.INIT(8'h96)) lut_n10610 (.I0(n10598), .I1(n10601), .I2(n10602), .O(n10610));
  LUT3 #(.INIT(8'hE8)) lut_n10611 (.I0(n10606), .I1(n10609), .I2(n10610), .O(n10611));
  LUT3 #(.INIT(8'h96)) lut_n10612 (.I0(n10583), .I1(n10591), .I2(n10592), .O(n10612));
  LUT3 #(.INIT(8'hE8)) lut_n10613 (.I0(n10603), .I1(n10611), .I2(n10612), .O(n10613));
  LUT3 #(.INIT(8'h96)) lut_n10614 (.I0(x1734), .I1(x1735), .I2(x1736), .O(n10614));
  LUT5 #(.INIT(32'h96696996)) lut_n10615 (.I0(x1725), .I1(x1726), .I2(x1727), .I3(n10607), .I4(n10608), .O(n10615));
  LUT5 #(.INIT(32'hFF969600)) lut_n10616 (.I0(x1731), .I1(x1732), .I2(x1733), .I3(n10614), .I4(n10615), .O(n10616));
  LUT3 #(.INIT(8'h96)) lut_n10617 (.I0(x1740), .I1(x1741), .I2(x1742), .O(n10617));
  LUT5 #(.INIT(32'h96696996)) lut_n10618 (.I0(x1731), .I1(x1732), .I2(x1733), .I3(n10614), .I4(n10615), .O(n10618));
  LUT5 #(.INIT(32'hFF969600)) lut_n10619 (.I0(x1737), .I1(x1738), .I2(x1739), .I3(n10617), .I4(n10618), .O(n10619));
  LUT3 #(.INIT(8'h96)) lut_n10620 (.I0(n10606), .I1(n10609), .I2(n10610), .O(n10620));
  LUT3 #(.INIT(8'hE8)) lut_n10621 (.I0(n10616), .I1(n10619), .I2(n10620), .O(n10621));
  LUT3 #(.INIT(8'h96)) lut_n10622 (.I0(x1746), .I1(x1747), .I2(x1748), .O(n10622));
  LUT5 #(.INIT(32'h96696996)) lut_n10623 (.I0(x1737), .I1(x1738), .I2(x1739), .I3(n10617), .I4(n10618), .O(n10623));
  LUT5 #(.INIT(32'hFF969600)) lut_n10624 (.I0(x1743), .I1(x1744), .I2(x1745), .I3(n10622), .I4(n10623), .O(n10624));
  LUT3 #(.INIT(8'h96)) lut_n10625 (.I0(x1752), .I1(x1753), .I2(x1754), .O(n10625));
  LUT5 #(.INIT(32'h96696996)) lut_n10626 (.I0(x1743), .I1(x1744), .I2(x1745), .I3(n10622), .I4(n10623), .O(n10626));
  LUT5 #(.INIT(32'hFF969600)) lut_n10627 (.I0(x1749), .I1(x1750), .I2(x1751), .I3(n10625), .I4(n10626), .O(n10627));
  LUT3 #(.INIT(8'h96)) lut_n10628 (.I0(n10616), .I1(n10619), .I2(n10620), .O(n10628));
  LUT3 #(.INIT(8'hE8)) lut_n10629 (.I0(n10624), .I1(n10627), .I2(n10628), .O(n10629));
  LUT3 #(.INIT(8'h96)) lut_n10630 (.I0(n10603), .I1(n10611), .I2(n10612), .O(n10630));
  LUT3 #(.INIT(8'hE8)) lut_n10631 (.I0(n10621), .I1(n10629), .I2(n10630), .O(n10631));
  LUT3 #(.INIT(8'h96)) lut_n10632 (.I0(n10575), .I1(n10593), .I2(n10594), .O(n10632));
  LUT3 #(.INIT(8'hE8)) lut_n10633 (.I0(n10613), .I1(n10631), .I2(n10632), .O(n10633));
  LUT3 #(.INIT(8'h96)) lut_n10634 (.I0(n10515), .I1(n10553), .I2(n10554), .O(n10634));
  LUT3 #(.INIT(8'hE8)) lut_n10635 (.I0(n10595), .I1(n10633), .I2(n10634), .O(n10635));
  LUT3 #(.INIT(8'h96)) lut_n10636 (.I0(x1758), .I1(x1759), .I2(x1760), .O(n10636));
  LUT5 #(.INIT(32'h96696996)) lut_n10637 (.I0(x1749), .I1(x1750), .I2(x1751), .I3(n10625), .I4(n10626), .O(n10637));
  LUT5 #(.INIT(32'hFF969600)) lut_n10638 (.I0(x1755), .I1(x1756), .I2(x1757), .I3(n10636), .I4(n10637), .O(n10638));
  LUT3 #(.INIT(8'h96)) lut_n10639 (.I0(x1764), .I1(x1765), .I2(x1766), .O(n10639));
  LUT5 #(.INIT(32'h96696996)) lut_n10640 (.I0(x1755), .I1(x1756), .I2(x1757), .I3(n10636), .I4(n10637), .O(n10640));
  LUT5 #(.INIT(32'hFF969600)) lut_n10641 (.I0(x1761), .I1(x1762), .I2(x1763), .I3(n10639), .I4(n10640), .O(n10641));
  LUT3 #(.INIT(8'h96)) lut_n10642 (.I0(n10624), .I1(n10627), .I2(n10628), .O(n10642));
  LUT3 #(.INIT(8'hE8)) lut_n10643 (.I0(n10638), .I1(n10641), .I2(n10642), .O(n10643));
  LUT3 #(.INIT(8'h96)) lut_n10644 (.I0(x1770), .I1(x1771), .I2(x1772), .O(n10644));
  LUT5 #(.INIT(32'h96696996)) lut_n10645 (.I0(x1761), .I1(x1762), .I2(x1763), .I3(n10639), .I4(n10640), .O(n10645));
  LUT5 #(.INIT(32'hFF969600)) lut_n10646 (.I0(x1767), .I1(x1768), .I2(x1769), .I3(n10644), .I4(n10645), .O(n10646));
  LUT3 #(.INIT(8'h96)) lut_n10647 (.I0(x1776), .I1(x1777), .I2(x1778), .O(n10647));
  LUT5 #(.INIT(32'h96696996)) lut_n10648 (.I0(x1767), .I1(x1768), .I2(x1769), .I3(n10644), .I4(n10645), .O(n10648));
  LUT5 #(.INIT(32'hFF969600)) lut_n10649 (.I0(x1773), .I1(x1774), .I2(x1775), .I3(n10647), .I4(n10648), .O(n10649));
  LUT3 #(.INIT(8'h96)) lut_n10650 (.I0(n10638), .I1(n10641), .I2(n10642), .O(n10650));
  LUT3 #(.INIT(8'hE8)) lut_n10651 (.I0(n10646), .I1(n10649), .I2(n10650), .O(n10651));
  LUT3 #(.INIT(8'h96)) lut_n10652 (.I0(n10621), .I1(n10629), .I2(n10630), .O(n10652));
  LUT3 #(.INIT(8'hE8)) lut_n10653 (.I0(n10643), .I1(n10651), .I2(n10652), .O(n10653));
  LUT3 #(.INIT(8'h96)) lut_n10654 (.I0(x1782), .I1(x1783), .I2(x1784), .O(n10654));
  LUT5 #(.INIT(32'h96696996)) lut_n10655 (.I0(x1773), .I1(x1774), .I2(x1775), .I3(n10647), .I4(n10648), .O(n10655));
  LUT5 #(.INIT(32'hFF969600)) lut_n10656 (.I0(x1779), .I1(x1780), .I2(x1781), .I3(n10654), .I4(n10655), .O(n10656));
  LUT3 #(.INIT(8'h96)) lut_n10657 (.I0(x1788), .I1(x1789), .I2(x1790), .O(n10657));
  LUT5 #(.INIT(32'h96696996)) lut_n10658 (.I0(x1779), .I1(x1780), .I2(x1781), .I3(n10654), .I4(n10655), .O(n10658));
  LUT5 #(.INIT(32'hFF969600)) lut_n10659 (.I0(x1785), .I1(x1786), .I2(x1787), .I3(n10657), .I4(n10658), .O(n10659));
  LUT3 #(.INIT(8'h96)) lut_n10660 (.I0(n10646), .I1(n10649), .I2(n10650), .O(n10660));
  LUT3 #(.INIT(8'hE8)) lut_n10661 (.I0(n10656), .I1(n10659), .I2(n10660), .O(n10661));
  LUT3 #(.INIT(8'h96)) lut_n10662 (.I0(x1794), .I1(x1795), .I2(x1796), .O(n10662));
  LUT5 #(.INIT(32'h96696996)) lut_n10663 (.I0(x1785), .I1(x1786), .I2(x1787), .I3(n10657), .I4(n10658), .O(n10663));
  LUT5 #(.INIT(32'hFF969600)) lut_n10664 (.I0(x1791), .I1(x1792), .I2(x1793), .I3(n10662), .I4(n10663), .O(n10664));
  LUT3 #(.INIT(8'h96)) lut_n10665 (.I0(x1800), .I1(x1801), .I2(x1802), .O(n10665));
  LUT5 #(.INIT(32'h96696996)) lut_n10666 (.I0(x1791), .I1(x1792), .I2(x1793), .I3(n10662), .I4(n10663), .O(n10666));
  LUT5 #(.INIT(32'hFF969600)) lut_n10667 (.I0(x1797), .I1(x1798), .I2(x1799), .I3(n10665), .I4(n10666), .O(n10667));
  LUT3 #(.INIT(8'h96)) lut_n10668 (.I0(n10656), .I1(n10659), .I2(n10660), .O(n10668));
  LUT3 #(.INIT(8'hE8)) lut_n10669 (.I0(n10664), .I1(n10667), .I2(n10668), .O(n10669));
  LUT3 #(.INIT(8'h96)) lut_n10670 (.I0(n10643), .I1(n10651), .I2(n10652), .O(n10670));
  LUT3 #(.INIT(8'hE8)) lut_n10671 (.I0(n10661), .I1(n10669), .I2(n10670), .O(n10671));
  LUT3 #(.INIT(8'h96)) lut_n10672 (.I0(n10613), .I1(n10631), .I2(n10632), .O(n10672));
  LUT3 #(.INIT(8'hE8)) lut_n10673 (.I0(n10653), .I1(n10671), .I2(n10672), .O(n10673));
  LUT3 #(.INIT(8'h96)) lut_n10674 (.I0(x1806), .I1(x1807), .I2(x1808), .O(n10674));
  LUT5 #(.INIT(32'h96696996)) lut_n10675 (.I0(x1797), .I1(x1798), .I2(x1799), .I3(n10665), .I4(n10666), .O(n10675));
  LUT5 #(.INIT(32'hFF969600)) lut_n10676 (.I0(x1803), .I1(x1804), .I2(x1805), .I3(n10674), .I4(n10675), .O(n10676));
  LUT3 #(.INIT(8'h96)) lut_n10677 (.I0(x1812), .I1(x1813), .I2(x1814), .O(n10677));
  LUT5 #(.INIT(32'h96696996)) lut_n10678 (.I0(x1803), .I1(x1804), .I2(x1805), .I3(n10674), .I4(n10675), .O(n10678));
  LUT5 #(.INIT(32'hFF969600)) lut_n10679 (.I0(x1809), .I1(x1810), .I2(x1811), .I3(n10677), .I4(n10678), .O(n10679));
  LUT3 #(.INIT(8'h96)) lut_n10680 (.I0(n10664), .I1(n10667), .I2(n10668), .O(n10680));
  LUT3 #(.INIT(8'hE8)) lut_n10681 (.I0(n10676), .I1(n10679), .I2(n10680), .O(n10681));
  LUT3 #(.INIT(8'h96)) lut_n10682 (.I0(x1818), .I1(x1819), .I2(x1820), .O(n10682));
  LUT5 #(.INIT(32'h96696996)) lut_n10683 (.I0(x1809), .I1(x1810), .I2(x1811), .I3(n10677), .I4(n10678), .O(n10683));
  LUT5 #(.INIT(32'hFF969600)) lut_n10684 (.I0(x1815), .I1(x1816), .I2(x1817), .I3(n10682), .I4(n10683), .O(n10684));
  LUT3 #(.INIT(8'h96)) lut_n10685 (.I0(x1824), .I1(x1825), .I2(x1826), .O(n10685));
  LUT5 #(.INIT(32'h96696996)) lut_n10686 (.I0(x1815), .I1(x1816), .I2(x1817), .I3(n10682), .I4(n10683), .O(n10686));
  LUT5 #(.INIT(32'hFF969600)) lut_n10687 (.I0(x1821), .I1(x1822), .I2(x1823), .I3(n10685), .I4(n10686), .O(n10687));
  LUT3 #(.INIT(8'h96)) lut_n10688 (.I0(n10676), .I1(n10679), .I2(n10680), .O(n10688));
  LUT3 #(.INIT(8'hE8)) lut_n10689 (.I0(n10684), .I1(n10687), .I2(n10688), .O(n10689));
  LUT3 #(.INIT(8'h96)) lut_n10690 (.I0(n10661), .I1(n10669), .I2(n10670), .O(n10690));
  LUT3 #(.INIT(8'hE8)) lut_n10691 (.I0(n10681), .I1(n10689), .I2(n10690), .O(n10691));
  LUT3 #(.INIT(8'h96)) lut_n10692 (.I0(x1830), .I1(x1831), .I2(x1832), .O(n10692));
  LUT5 #(.INIT(32'h96696996)) lut_n10693 (.I0(x1821), .I1(x1822), .I2(x1823), .I3(n10685), .I4(n10686), .O(n10693));
  LUT5 #(.INIT(32'hFF969600)) lut_n10694 (.I0(x1827), .I1(x1828), .I2(x1829), .I3(n10692), .I4(n10693), .O(n10694));
  LUT3 #(.INIT(8'h96)) lut_n10695 (.I0(x1836), .I1(x1837), .I2(x1838), .O(n10695));
  LUT5 #(.INIT(32'h96696996)) lut_n10696 (.I0(x1827), .I1(x1828), .I2(x1829), .I3(n10692), .I4(n10693), .O(n10696));
  LUT5 #(.INIT(32'hFF969600)) lut_n10697 (.I0(x1833), .I1(x1834), .I2(x1835), .I3(n10695), .I4(n10696), .O(n10697));
  LUT3 #(.INIT(8'h96)) lut_n10698 (.I0(n10684), .I1(n10687), .I2(n10688), .O(n10698));
  LUT3 #(.INIT(8'hE8)) lut_n10699 (.I0(n10694), .I1(n10697), .I2(n10698), .O(n10699));
  LUT3 #(.INIT(8'h96)) lut_n10700 (.I0(x1842), .I1(x1843), .I2(x1844), .O(n10700));
  LUT5 #(.INIT(32'h96696996)) lut_n10701 (.I0(x1833), .I1(x1834), .I2(x1835), .I3(n10695), .I4(n10696), .O(n10701));
  LUT5 #(.INIT(32'hFF969600)) lut_n10702 (.I0(x1839), .I1(x1840), .I2(x1841), .I3(n10700), .I4(n10701), .O(n10702));
  LUT3 #(.INIT(8'h96)) lut_n10703 (.I0(x1848), .I1(x1849), .I2(x1850), .O(n10703));
  LUT5 #(.INIT(32'h96696996)) lut_n10704 (.I0(x1839), .I1(x1840), .I2(x1841), .I3(n10700), .I4(n10701), .O(n10704));
  LUT5 #(.INIT(32'hFF969600)) lut_n10705 (.I0(x1845), .I1(x1846), .I2(x1847), .I3(n10703), .I4(n10704), .O(n10705));
  LUT3 #(.INIT(8'h96)) lut_n10706 (.I0(n10694), .I1(n10697), .I2(n10698), .O(n10706));
  LUT3 #(.INIT(8'hE8)) lut_n10707 (.I0(n10702), .I1(n10705), .I2(n10706), .O(n10707));
  LUT3 #(.INIT(8'h96)) lut_n10708 (.I0(n10681), .I1(n10689), .I2(n10690), .O(n10708));
  LUT3 #(.INIT(8'hE8)) lut_n10709 (.I0(n10699), .I1(n10707), .I2(n10708), .O(n10709));
  LUT3 #(.INIT(8'h96)) lut_n10710 (.I0(n10653), .I1(n10671), .I2(n10672), .O(n10710));
  LUT3 #(.INIT(8'hE8)) lut_n10711 (.I0(n10691), .I1(n10709), .I2(n10710), .O(n10711));
  LUT3 #(.INIT(8'h96)) lut_n10712 (.I0(n10595), .I1(n10633), .I2(n10634), .O(n10712));
  LUT3 #(.INIT(8'hE8)) lut_n10713 (.I0(n10673), .I1(n10711), .I2(n10712), .O(n10713));
  LUT3 #(.INIT(8'h96)) lut_n10714 (.I0(n10477), .I1(n10555), .I2(n10556), .O(n10714));
  LUT3 #(.INIT(8'hE8)) lut_n10715 (.I0(n10635), .I1(n10713), .I2(n10714), .O(n10715));
  LUT3 #(.INIT(8'h96)) lut_n10716 (.I0(n10237), .I1(n10395), .I2(n10396), .O(n10716));
  LUT3 #(.INIT(8'hE8)) lut_n10717 (.I0(n10557), .I1(n10715), .I2(n10716), .O(n10717));
  LUT3 #(.INIT(8'h96)) lut_n10718 (.I0(x1854), .I1(x1855), .I2(x1856), .O(n10718));
  LUT5 #(.INIT(32'h96696996)) lut_n10719 (.I0(x1845), .I1(x1846), .I2(x1847), .I3(n10703), .I4(n10704), .O(n10719));
  LUT5 #(.INIT(32'hFF969600)) lut_n10720 (.I0(x1851), .I1(x1852), .I2(x1853), .I3(n10718), .I4(n10719), .O(n10720));
  LUT3 #(.INIT(8'h96)) lut_n10721 (.I0(x1860), .I1(x1861), .I2(x1862), .O(n10721));
  LUT5 #(.INIT(32'h96696996)) lut_n10722 (.I0(x1851), .I1(x1852), .I2(x1853), .I3(n10718), .I4(n10719), .O(n10722));
  LUT5 #(.INIT(32'hFF969600)) lut_n10723 (.I0(x1857), .I1(x1858), .I2(x1859), .I3(n10721), .I4(n10722), .O(n10723));
  LUT3 #(.INIT(8'h96)) lut_n10724 (.I0(n10702), .I1(n10705), .I2(n10706), .O(n10724));
  LUT3 #(.INIT(8'hE8)) lut_n10725 (.I0(n10720), .I1(n10723), .I2(n10724), .O(n10725));
  LUT3 #(.INIT(8'h96)) lut_n10726 (.I0(x1866), .I1(x1867), .I2(x1868), .O(n10726));
  LUT5 #(.INIT(32'h96696996)) lut_n10727 (.I0(x1857), .I1(x1858), .I2(x1859), .I3(n10721), .I4(n10722), .O(n10727));
  LUT5 #(.INIT(32'hFF969600)) lut_n10728 (.I0(x1863), .I1(x1864), .I2(x1865), .I3(n10726), .I4(n10727), .O(n10728));
  LUT3 #(.INIT(8'h96)) lut_n10729 (.I0(x1872), .I1(x1873), .I2(x1874), .O(n10729));
  LUT5 #(.INIT(32'h96696996)) lut_n10730 (.I0(x1863), .I1(x1864), .I2(x1865), .I3(n10726), .I4(n10727), .O(n10730));
  LUT5 #(.INIT(32'hFF969600)) lut_n10731 (.I0(x1869), .I1(x1870), .I2(x1871), .I3(n10729), .I4(n10730), .O(n10731));
  LUT3 #(.INIT(8'h96)) lut_n10732 (.I0(n10720), .I1(n10723), .I2(n10724), .O(n10732));
  LUT3 #(.INIT(8'hE8)) lut_n10733 (.I0(n10728), .I1(n10731), .I2(n10732), .O(n10733));
  LUT3 #(.INIT(8'h96)) lut_n10734 (.I0(n10699), .I1(n10707), .I2(n10708), .O(n10734));
  LUT3 #(.INIT(8'hE8)) lut_n10735 (.I0(n10725), .I1(n10733), .I2(n10734), .O(n10735));
  LUT3 #(.INIT(8'h96)) lut_n10736 (.I0(x1878), .I1(x1879), .I2(x1880), .O(n10736));
  LUT5 #(.INIT(32'h96696996)) lut_n10737 (.I0(x1869), .I1(x1870), .I2(x1871), .I3(n10729), .I4(n10730), .O(n10737));
  LUT5 #(.INIT(32'hFF969600)) lut_n10738 (.I0(x1875), .I1(x1876), .I2(x1877), .I3(n10736), .I4(n10737), .O(n10738));
  LUT3 #(.INIT(8'h96)) lut_n10739 (.I0(x1884), .I1(x1885), .I2(x1886), .O(n10739));
  LUT5 #(.INIT(32'h96696996)) lut_n10740 (.I0(x1875), .I1(x1876), .I2(x1877), .I3(n10736), .I4(n10737), .O(n10740));
  LUT5 #(.INIT(32'hFF969600)) lut_n10741 (.I0(x1881), .I1(x1882), .I2(x1883), .I3(n10739), .I4(n10740), .O(n10741));
  LUT3 #(.INIT(8'h96)) lut_n10742 (.I0(n10728), .I1(n10731), .I2(n10732), .O(n10742));
  LUT3 #(.INIT(8'hE8)) lut_n10743 (.I0(n10738), .I1(n10741), .I2(n10742), .O(n10743));
  LUT3 #(.INIT(8'h96)) lut_n10744 (.I0(x1890), .I1(x1891), .I2(x1892), .O(n10744));
  LUT5 #(.INIT(32'h96696996)) lut_n10745 (.I0(x1881), .I1(x1882), .I2(x1883), .I3(n10739), .I4(n10740), .O(n10745));
  LUT5 #(.INIT(32'hFF969600)) lut_n10746 (.I0(x1887), .I1(x1888), .I2(x1889), .I3(n10744), .I4(n10745), .O(n10746));
  LUT3 #(.INIT(8'h96)) lut_n10747 (.I0(x1896), .I1(x1897), .I2(x1898), .O(n10747));
  LUT5 #(.INIT(32'h96696996)) lut_n10748 (.I0(x1887), .I1(x1888), .I2(x1889), .I3(n10744), .I4(n10745), .O(n10748));
  LUT5 #(.INIT(32'hFF969600)) lut_n10749 (.I0(x1893), .I1(x1894), .I2(x1895), .I3(n10747), .I4(n10748), .O(n10749));
  LUT3 #(.INIT(8'h96)) lut_n10750 (.I0(n10738), .I1(n10741), .I2(n10742), .O(n10750));
  LUT3 #(.INIT(8'hE8)) lut_n10751 (.I0(n10746), .I1(n10749), .I2(n10750), .O(n10751));
  LUT3 #(.INIT(8'h96)) lut_n10752 (.I0(n10725), .I1(n10733), .I2(n10734), .O(n10752));
  LUT3 #(.INIT(8'hE8)) lut_n10753 (.I0(n10743), .I1(n10751), .I2(n10752), .O(n10753));
  LUT3 #(.INIT(8'h96)) lut_n10754 (.I0(n10691), .I1(n10709), .I2(n10710), .O(n10754));
  LUT3 #(.INIT(8'hE8)) lut_n10755 (.I0(n10735), .I1(n10753), .I2(n10754), .O(n10755));
  LUT3 #(.INIT(8'h96)) lut_n10756 (.I0(x1902), .I1(x1903), .I2(x1904), .O(n10756));
  LUT5 #(.INIT(32'h96696996)) lut_n10757 (.I0(x1893), .I1(x1894), .I2(x1895), .I3(n10747), .I4(n10748), .O(n10757));
  LUT5 #(.INIT(32'hFF969600)) lut_n10758 (.I0(x1899), .I1(x1900), .I2(x1901), .I3(n10756), .I4(n10757), .O(n10758));
  LUT3 #(.INIT(8'h96)) lut_n10759 (.I0(x1908), .I1(x1909), .I2(x1910), .O(n10759));
  LUT5 #(.INIT(32'h96696996)) lut_n10760 (.I0(x1899), .I1(x1900), .I2(x1901), .I3(n10756), .I4(n10757), .O(n10760));
  LUT5 #(.INIT(32'hFF969600)) lut_n10761 (.I0(x1905), .I1(x1906), .I2(x1907), .I3(n10759), .I4(n10760), .O(n10761));
  LUT3 #(.INIT(8'h96)) lut_n10762 (.I0(n10746), .I1(n10749), .I2(n10750), .O(n10762));
  LUT3 #(.INIT(8'hE8)) lut_n10763 (.I0(n10758), .I1(n10761), .I2(n10762), .O(n10763));
  LUT3 #(.INIT(8'h96)) lut_n10764 (.I0(x1914), .I1(x1915), .I2(x1916), .O(n10764));
  LUT5 #(.INIT(32'h96696996)) lut_n10765 (.I0(x1905), .I1(x1906), .I2(x1907), .I3(n10759), .I4(n10760), .O(n10765));
  LUT5 #(.INIT(32'hFF969600)) lut_n10766 (.I0(x1911), .I1(x1912), .I2(x1913), .I3(n10764), .I4(n10765), .O(n10766));
  LUT3 #(.INIT(8'h96)) lut_n10767 (.I0(x1920), .I1(x1921), .I2(x1922), .O(n10767));
  LUT5 #(.INIT(32'h96696996)) lut_n10768 (.I0(x1911), .I1(x1912), .I2(x1913), .I3(n10764), .I4(n10765), .O(n10768));
  LUT5 #(.INIT(32'hFF969600)) lut_n10769 (.I0(x1917), .I1(x1918), .I2(x1919), .I3(n10767), .I4(n10768), .O(n10769));
  LUT3 #(.INIT(8'h96)) lut_n10770 (.I0(n10758), .I1(n10761), .I2(n10762), .O(n10770));
  LUT3 #(.INIT(8'hE8)) lut_n10771 (.I0(n10766), .I1(n10769), .I2(n10770), .O(n10771));
  LUT3 #(.INIT(8'h96)) lut_n10772 (.I0(n10743), .I1(n10751), .I2(n10752), .O(n10772));
  LUT3 #(.INIT(8'hE8)) lut_n10773 (.I0(n10763), .I1(n10771), .I2(n10772), .O(n10773));
  LUT3 #(.INIT(8'h96)) lut_n10774 (.I0(x1926), .I1(x1927), .I2(x1928), .O(n10774));
  LUT5 #(.INIT(32'h96696996)) lut_n10775 (.I0(x1917), .I1(x1918), .I2(x1919), .I3(n10767), .I4(n10768), .O(n10775));
  LUT5 #(.INIT(32'hFF969600)) lut_n10776 (.I0(x1923), .I1(x1924), .I2(x1925), .I3(n10774), .I4(n10775), .O(n10776));
  LUT3 #(.INIT(8'h96)) lut_n10777 (.I0(x1932), .I1(x1933), .I2(x1934), .O(n10777));
  LUT5 #(.INIT(32'h96696996)) lut_n10778 (.I0(x1923), .I1(x1924), .I2(x1925), .I3(n10774), .I4(n10775), .O(n10778));
  LUT5 #(.INIT(32'hFF969600)) lut_n10779 (.I0(x1929), .I1(x1930), .I2(x1931), .I3(n10777), .I4(n10778), .O(n10779));
  LUT3 #(.INIT(8'h96)) lut_n10780 (.I0(n10766), .I1(n10769), .I2(n10770), .O(n10780));
  LUT3 #(.INIT(8'hE8)) lut_n10781 (.I0(n10776), .I1(n10779), .I2(n10780), .O(n10781));
  LUT3 #(.INIT(8'h96)) lut_n10782 (.I0(x1938), .I1(x1939), .I2(x1940), .O(n10782));
  LUT5 #(.INIT(32'h96696996)) lut_n10783 (.I0(x1929), .I1(x1930), .I2(x1931), .I3(n10777), .I4(n10778), .O(n10783));
  LUT5 #(.INIT(32'hFF969600)) lut_n10784 (.I0(x1935), .I1(x1936), .I2(x1937), .I3(n10782), .I4(n10783), .O(n10784));
  LUT3 #(.INIT(8'h96)) lut_n10785 (.I0(x1944), .I1(x1945), .I2(x1946), .O(n10785));
  LUT5 #(.INIT(32'h96696996)) lut_n10786 (.I0(x1935), .I1(x1936), .I2(x1937), .I3(n10782), .I4(n10783), .O(n10786));
  LUT5 #(.INIT(32'hFF969600)) lut_n10787 (.I0(x1941), .I1(x1942), .I2(x1943), .I3(n10785), .I4(n10786), .O(n10787));
  LUT3 #(.INIT(8'h96)) lut_n10788 (.I0(n10776), .I1(n10779), .I2(n10780), .O(n10788));
  LUT3 #(.INIT(8'hE8)) lut_n10789 (.I0(n10784), .I1(n10787), .I2(n10788), .O(n10789));
  LUT3 #(.INIT(8'h96)) lut_n10790 (.I0(n10763), .I1(n10771), .I2(n10772), .O(n10790));
  LUT3 #(.INIT(8'hE8)) lut_n10791 (.I0(n10781), .I1(n10789), .I2(n10790), .O(n10791));
  LUT3 #(.INIT(8'h96)) lut_n10792 (.I0(n10735), .I1(n10753), .I2(n10754), .O(n10792));
  LUT3 #(.INIT(8'hE8)) lut_n10793 (.I0(n10773), .I1(n10791), .I2(n10792), .O(n10793));
  LUT3 #(.INIT(8'h96)) lut_n10794 (.I0(n10673), .I1(n10711), .I2(n10712), .O(n10794));
  LUT3 #(.INIT(8'hE8)) lut_n10795 (.I0(n10755), .I1(n10793), .I2(n10794), .O(n10795));
  LUT3 #(.INIT(8'h96)) lut_n10796 (.I0(x1950), .I1(x1951), .I2(x1952), .O(n10796));
  LUT5 #(.INIT(32'h96696996)) lut_n10797 (.I0(x1941), .I1(x1942), .I2(x1943), .I3(n10785), .I4(n10786), .O(n10797));
  LUT5 #(.INIT(32'hFF969600)) lut_n10798 (.I0(x1947), .I1(x1948), .I2(x1949), .I3(n10796), .I4(n10797), .O(n10798));
  LUT3 #(.INIT(8'h96)) lut_n10799 (.I0(x1956), .I1(x1957), .I2(x1958), .O(n10799));
  LUT5 #(.INIT(32'h96696996)) lut_n10800 (.I0(x1947), .I1(x1948), .I2(x1949), .I3(n10796), .I4(n10797), .O(n10800));
  LUT5 #(.INIT(32'hFF969600)) lut_n10801 (.I0(x1953), .I1(x1954), .I2(x1955), .I3(n10799), .I4(n10800), .O(n10801));
  LUT3 #(.INIT(8'h96)) lut_n10802 (.I0(n10784), .I1(n10787), .I2(n10788), .O(n10802));
  LUT3 #(.INIT(8'hE8)) lut_n10803 (.I0(n10798), .I1(n10801), .I2(n10802), .O(n10803));
  LUT3 #(.INIT(8'h96)) lut_n10804 (.I0(x1962), .I1(x1963), .I2(x1964), .O(n10804));
  LUT5 #(.INIT(32'h96696996)) lut_n10805 (.I0(x1953), .I1(x1954), .I2(x1955), .I3(n10799), .I4(n10800), .O(n10805));
  LUT5 #(.INIT(32'hFF969600)) lut_n10806 (.I0(x1959), .I1(x1960), .I2(x1961), .I3(n10804), .I4(n10805), .O(n10806));
  LUT3 #(.INIT(8'h96)) lut_n10807 (.I0(x1968), .I1(x1969), .I2(x1970), .O(n10807));
  LUT5 #(.INIT(32'h96696996)) lut_n10808 (.I0(x1959), .I1(x1960), .I2(x1961), .I3(n10804), .I4(n10805), .O(n10808));
  LUT5 #(.INIT(32'hFF969600)) lut_n10809 (.I0(x1965), .I1(x1966), .I2(x1967), .I3(n10807), .I4(n10808), .O(n10809));
  LUT3 #(.INIT(8'h96)) lut_n10810 (.I0(n10798), .I1(n10801), .I2(n10802), .O(n10810));
  LUT3 #(.INIT(8'hE8)) lut_n10811 (.I0(n10806), .I1(n10809), .I2(n10810), .O(n10811));
  LUT3 #(.INIT(8'h96)) lut_n10812 (.I0(n10781), .I1(n10789), .I2(n10790), .O(n10812));
  LUT3 #(.INIT(8'hE8)) lut_n10813 (.I0(n10803), .I1(n10811), .I2(n10812), .O(n10813));
  LUT3 #(.INIT(8'h96)) lut_n10814 (.I0(x1974), .I1(x1975), .I2(x1976), .O(n10814));
  LUT5 #(.INIT(32'h96696996)) lut_n10815 (.I0(x1965), .I1(x1966), .I2(x1967), .I3(n10807), .I4(n10808), .O(n10815));
  LUT5 #(.INIT(32'hFF969600)) lut_n10816 (.I0(x1971), .I1(x1972), .I2(x1973), .I3(n10814), .I4(n10815), .O(n10816));
  LUT3 #(.INIT(8'h96)) lut_n10817 (.I0(x1980), .I1(x1981), .I2(x1982), .O(n10817));
  LUT5 #(.INIT(32'h96696996)) lut_n10818 (.I0(x1971), .I1(x1972), .I2(x1973), .I3(n10814), .I4(n10815), .O(n10818));
  LUT5 #(.INIT(32'hFF969600)) lut_n10819 (.I0(x1977), .I1(x1978), .I2(x1979), .I3(n10817), .I4(n10818), .O(n10819));
  LUT3 #(.INIT(8'h96)) lut_n10820 (.I0(n10806), .I1(n10809), .I2(n10810), .O(n10820));
  LUT3 #(.INIT(8'hE8)) lut_n10821 (.I0(n10816), .I1(n10819), .I2(n10820), .O(n10821));
  LUT3 #(.INIT(8'h96)) lut_n10822 (.I0(x1986), .I1(x1987), .I2(x1988), .O(n10822));
  LUT5 #(.INIT(32'h96696996)) lut_n10823 (.I0(x1977), .I1(x1978), .I2(x1979), .I3(n10817), .I4(n10818), .O(n10823));
  LUT5 #(.INIT(32'hFF969600)) lut_n10824 (.I0(x1983), .I1(x1984), .I2(x1985), .I3(n10822), .I4(n10823), .O(n10824));
  LUT3 #(.INIT(8'h96)) lut_n10825 (.I0(x1992), .I1(x1993), .I2(x1994), .O(n10825));
  LUT5 #(.INIT(32'h96696996)) lut_n10826 (.I0(x1983), .I1(x1984), .I2(x1985), .I3(n10822), .I4(n10823), .O(n10826));
  LUT5 #(.INIT(32'hFF969600)) lut_n10827 (.I0(x1989), .I1(x1990), .I2(x1991), .I3(n10825), .I4(n10826), .O(n10827));
  LUT3 #(.INIT(8'h96)) lut_n10828 (.I0(n10816), .I1(n10819), .I2(n10820), .O(n10828));
  LUT3 #(.INIT(8'hE8)) lut_n10829 (.I0(n10824), .I1(n10827), .I2(n10828), .O(n10829));
  LUT3 #(.INIT(8'h96)) lut_n10830 (.I0(n10803), .I1(n10811), .I2(n10812), .O(n10830));
  LUT3 #(.INIT(8'hE8)) lut_n10831 (.I0(n10821), .I1(n10829), .I2(n10830), .O(n10831));
  LUT3 #(.INIT(8'h96)) lut_n10832 (.I0(n10773), .I1(n10791), .I2(n10792), .O(n10832));
  LUT3 #(.INIT(8'hE8)) lut_n10833 (.I0(n10813), .I1(n10831), .I2(n10832), .O(n10833));
  LUT3 #(.INIT(8'h96)) lut_n10834 (.I0(x1998), .I1(x1999), .I2(x2000), .O(n10834));
  LUT5 #(.INIT(32'h96696996)) lut_n10835 (.I0(x1989), .I1(x1990), .I2(x1991), .I3(n10825), .I4(n10826), .O(n10835));
  LUT5 #(.INIT(32'hFF969600)) lut_n10836 (.I0(x1995), .I1(x1996), .I2(x1997), .I3(n10834), .I4(n10835), .O(n10836));
  LUT3 #(.INIT(8'h96)) lut_n10837 (.I0(x2004), .I1(x2005), .I2(x2006), .O(n10837));
  LUT5 #(.INIT(32'h96696996)) lut_n10838 (.I0(x1995), .I1(x1996), .I2(x1997), .I3(n10834), .I4(n10835), .O(n10838));
  LUT5 #(.INIT(32'hFF969600)) lut_n10839 (.I0(x2001), .I1(x2002), .I2(x2003), .I3(n10837), .I4(n10838), .O(n10839));
  LUT3 #(.INIT(8'h96)) lut_n10840 (.I0(n10824), .I1(n10827), .I2(n10828), .O(n10840));
  LUT3 #(.INIT(8'hE8)) lut_n10841 (.I0(n10836), .I1(n10839), .I2(n10840), .O(n10841));
  LUT3 #(.INIT(8'h96)) lut_n10842 (.I0(x2010), .I1(x2011), .I2(x2012), .O(n10842));
  LUT5 #(.INIT(32'h96696996)) lut_n10843 (.I0(x2001), .I1(x2002), .I2(x2003), .I3(n10837), .I4(n10838), .O(n10843));
  LUT5 #(.INIT(32'hFF969600)) lut_n10844 (.I0(x2007), .I1(x2008), .I2(x2009), .I3(n10842), .I4(n10843), .O(n10844));
  LUT3 #(.INIT(8'h96)) lut_n10845 (.I0(x2016), .I1(x2017), .I2(x2018), .O(n10845));
  LUT5 #(.INIT(32'h96696996)) lut_n10846 (.I0(x2007), .I1(x2008), .I2(x2009), .I3(n10842), .I4(n10843), .O(n10846));
  LUT5 #(.INIT(32'hFF969600)) lut_n10847 (.I0(x2013), .I1(x2014), .I2(x2015), .I3(n10845), .I4(n10846), .O(n10847));
  LUT3 #(.INIT(8'h96)) lut_n10848 (.I0(n10836), .I1(n10839), .I2(n10840), .O(n10848));
  LUT3 #(.INIT(8'hE8)) lut_n10849 (.I0(n10844), .I1(n10847), .I2(n10848), .O(n10849));
  LUT3 #(.INIT(8'h96)) lut_n10850 (.I0(n10821), .I1(n10829), .I2(n10830), .O(n10850));
  LUT3 #(.INIT(8'hE8)) lut_n10851 (.I0(n10841), .I1(n10849), .I2(n10850), .O(n10851));
  LUT3 #(.INIT(8'h96)) lut_n10852 (.I0(x2022), .I1(x2023), .I2(x2024), .O(n10852));
  LUT5 #(.INIT(32'h96696996)) lut_n10853 (.I0(x2013), .I1(x2014), .I2(x2015), .I3(n10845), .I4(n10846), .O(n10853));
  LUT5 #(.INIT(32'hFF969600)) lut_n10854 (.I0(x2019), .I1(x2020), .I2(x2021), .I3(n10852), .I4(n10853), .O(n10854));
  LUT3 #(.INIT(8'h96)) lut_n10855 (.I0(x2028), .I1(x2029), .I2(x2030), .O(n10855));
  LUT5 #(.INIT(32'h96696996)) lut_n10856 (.I0(x2019), .I1(x2020), .I2(x2021), .I3(n10852), .I4(n10853), .O(n10856));
  LUT5 #(.INIT(32'hFF969600)) lut_n10857 (.I0(x2025), .I1(x2026), .I2(x2027), .I3(n10855), .I4(n10856), .O(n10857));
  LUT3 #(.INIT(8'h96)) lut_n10858 (.I0(n10844), .I1(n10847), .I2(n10848), .O(n10858));
  LUT3 #(.INIT(8'hE8)) lut_n10859 (.I0(n10854), .I1(n10857), .I2(n10858), .O(n10859));
  LUT3 #(.INIT(8'h96)) lut_n10860 (.I0(x2034), .I1(x2035), .I2(x2036), .O(n10860));
  LUT5 #(.INIT(32'h96696996)) lut_n10861 (.I0(x2025), .I1(x2026), .I2(x2027), .I3(n10855), .I4(n10856), .O(n10861));
  LUT5 #(.INIT(32'hFF969600)) lut_n10862 (.I0(x2031), .I1(x2032), .I2(x2033), .I3(n10860), .I4(n10861), .O(n10862));
  LUT3 #(.INIT(8'h96)) lut_n10863 (.I0(x2040), .I1(x2041), .I2(x2042), .O(n10863));
  LUT5 #(.INIT(32'h96696996)) lut_n10864 (.I0(x2031), .I1(x2032), .I2(x2033), .I3(n10860), .I4(n10861), .O(n10864));
  LUT5 #(.INIT(32'hFF969600)) lut_n10865 (.I0(x2037), .I1(x2038), .I2(x2039), .I3(n10863), .I4(n10864), .O(n10865));
  LUT3 #(.INIT(8'h96)) lut_n10866 (.I0(n10854), .I1(n10857), .I2(n10858), .O(n10866));
  LUT3 #(.INIT(8'hE8)) lut_n10867 (.I0(n10862), .I1(n10865), .I2(n10866), .O(n10867));
  LUT3 #(.INIT(8'h96)) lut_n10868 (.I0(n10841), .I1(n10849), .I2(n10850), .O(n10868));
  LUT3 #(.INIT(8'hE8)) lut_n10869 (.I0(n10859), .I1(n10867), .I2(n10868), .O(n10869));
  LUT3 #(.INIT(8'h96)) lut_n10870 (.I0(n10813), .I1(n10831), .I2(n10832), .O(n10870));
  LUT3 #(.INIT(8'hE8)) lut_n10871 (.I0(n10851), .I1(n10869), .I2(n10870), .O(n10871));
  LUT3 #(.INIT(8'h96)) lut_n10872 (.I0(n10755), .I1(n10793), .I2(n10794), .O(n10872));
  LUT3 #(.INIT(8'hE8)) lut_n10873 (.I0(n10833), .I1(n10871), .I2(n10872), .O(n10873));
  LUT3 #(.INIT(8'h96)) lut_n10874 (.I0(n10635), .I1(n10713), .I2(n10714), .O(n10874));
  LUT3 #(.INIT(8'hE8)) lut_n10875 (.I0(n10795), .I1(n10873), .I2(n10874), .O(n10875));
  LUT3 #(.INIT(8'h96)) lut_n10876 (.I0(x2046), .I1(x2047), .I2(x2048), .O(n10876));
  LUT5 #(.INIT(32'h96696996)) lut_n10877 (.I0(x2037), .I1(x2038), .I2(x2039), .I3(n10863), .I4(n10864), .O(n10877));
  LUT5 #(.INIT(32'hFF969600)) lut_n10878 (.I0(x2043), .I1(x2044), .I2(x2045), .I3(n10876), .I4(n10877), .O(n10878));
  LUT3 #(.INIT(8'h96)) lut_n10879 (.I0(x2052), .I1(x2053), .I2(x2054), .O(n10879));
  LUT5 #(.INIT(32'h96696996)) lut_n10880 (.I0(x2043), .I1(x2044), .I2(x2045), .I3(n10876), .I4(n10877), .O(n10880));
  LUT5 #(.INIT(32'hFF969600)) lut_n10881 (.I0(x2049), .I1(x2050), .I2(x2051), .I3(n10879), .I4(n10880), .O(n10881));
  LUT3 #(.INIT(8'h96)) lut_n10882 (.I0(n10862), .I1(n10865), .I2(n10866), .O(n10882));
  LUT3 #(.INIT(8'hE8)) lut_n10883 (.I0(n10878), .I1(n10881), .I2(n10882), .O(n10883));
  LUT3 #(.INIT(8'h96)) lut_n10884 (.I0(x2058), .I1(x2059), .I2(x2060), .O(n10884));
  LUT5 #(.INIT(32'h96696996)) lut_n10885 (.I0(x2049), .I1(x2050), .I2(x2051), .I3(n10879), .I4(n10880), .O(n10885));
  LUT5 #(.INIT(32'hFF969600)) lut_n10886 (.I0(x2055), .I1(x2056), .I2(x2057), .I3(n10884), .I4(n10885), .O(n10886));
  LUT3 #(.INIT(8'h96)) lut_n10887 (.I0(x2064), .I1(x2065), .I2(x2066), .O(n10887));
  LUT5 #(.INIT(32'h96696996)) lut_n10888 (.I0(x2055), .I1(x2056), .I2(x2057), .I3(n10884), .I4(n10885), .O(n10888));
  LUT5 #(.INIT(32'hFF969600)) lut_n10889 (.I0(x2061), .I1(x2062), .I2(x2063), .I3(n10887), .I4(n10888), .O(n10889));
  LUT3 #(.INIT(8'h96)) lut_n10890 (.I0(n10878), .I1(n10881), .I2(n10882), .O(n10890));
  LUT3 #(.INIT(8'hE8)) lut_n10891 (.I0(n10886), .I1(n10889), .I2(n10890), .O(n10891));
  LUT3 #(.INIT(8'h96)) lut_n10892 (.I0(n10859), .I1(n10867), .I2(n10868), .O(n10892));
  LUT3 #(.INIT(8'hE8)) lut_n10893 (.I0(n10883), .I1(n10891), .I2(n10892), .O(n10893));
  LUT3 #(.INIT(8'h96)) lut_n10894 (.I0(x2070), .I1(x2071), .I2(x2072), .O(n10894));
  LUT5 #(.INIT(32'h96696996)) lut_n10895 (.I0(x2061), .I1(x2062), .I2(x2063), .I3(n10887), .I4(n10888), .O(n10895));
  LUT5 #(.INIT(32'hFF969600)) lut_n10896 (.I0(x2067), .I1(x2068), .I2(x2069), .I3(n10894), .I4(n10895), .O(n10896));
  LUT3 #(.INIT(8'h96)) lut_n10897 (.I0(x2076), .I1(x2077), .I2(x2078), .O(n10897));
  LUT5 #(.INIT(32'h96696996)) lut_n10898 (.I0(x2067), .I1(x2068), .I2(x2069), .I3(n10894), .I4(n10895), .O(n10898));
  LUT5 #(.INIT(32'hFF969600)) lut_n10899 (.I0(x2073), .I1(x2074), .I2(x2075), .I3(n10897), .I4(n10898), .O(n10899));
  LUT3 #(.INIT(8'h96)) lut_n10900 (.I0(n10886), .I1(n10889), .I2(n10890), .O(n10900));
  LUT3 #(.INIT(8'hE8)) lut_n10901 (.I0(n10896), .I1(n10899), .I2(n10900), .O(n10901));
  LUT3 #(.INIT(8'h96)) lut_n10902 (.I0(x2082), .I1(x2083), .I2(x2084), .O(n10902));
  LUT5 #(.INIT(32'h96696996)) lut_n10903 (.I0(x2073), .I1(x2074), .I2(x2075), .I3(n10897), .I4(n10898), .O(n10903));
  LUT5 #(.INIT(32'hFF969600)) lut_n10904 (.I0(x2079), .I1(x2080), .I2(x2081), .I3(n10902), .I4(n10903), .O(n10904));
  LUT3 #(.INIT(8'h96)) lut_n10905 (.I0(x2088), .I1(x2089), .I2(x2090), .O(n10905));
  LUT5 #(.INIT(32'h96696996)) lut_n10906 (.I0(x2079), .I1(x2080), .I2(x2081), .I3(n10902), .I4(n10903), .O(n10906));
  LUT5 #(.INIT(32'hFF969600)) lut_n10907 (.I0(x2085), .I1(x2086), .I2(x2087), .I3(n10905), .I4(n10906), .O(n10907));
  LUT3 #(.INIT(8'h96)) lut_n10908 (.I0(n10896), .I1(n10899), .I2(n10900), .O(n10908));
  LUT3 #(.INIT(8'hE8)) lut_n10909 (.I0(n10904), .I1(n10907), .I2(n10908), .O(n10909));
  LUT3 #(.INIT(8'h96)) lut_n10910 (.I0(n10883), .I1(n10891), .I2(n10892), .O(n10910));
  LUT3 #(.INIT(8'hE8)) lut_n10911 (.I0(n10901), .I1(n10909), .I2(n10910), .O(n10911));
  LUT3 #(.INIT(8'h96)) lut_n10912 (.I0(n10851), .I1(n10869), .I2(n10870), .O(n10912));
  LUT3 #(.INIT(8'hE8)) lut_n10913 (.I0(n10893), .I1(n10911), .I2(n10912), .O(n10913));
  LUT3 #(.INIT(8'h96)) lut_n10914 (.I0(x2094), .I1(x2095), .I2(x2096), .O(n10914));
  LUT5 #(.INIT(32'h96696996)) lut_n10915 (.I0(x2085), .I1(x2086), .I2(x2087), .I3(n10905), .I4(n10906), .O(n10915));
  LUT5 #(.INIT(32'hFF969600)) lut_n10916 (.I0(x2091), .I1(x2092), .I2(x2093), .I3(n10914), .I4(n10915), .O(n10916));
  LUT3 #(.INIT(8'h96)) lut_n10917 (.I0(x2100), .I1(x2101), .I2(x2102), .O(n10917));
  LUT5 #(.INIT(32'h96696996)) lut_n10918 (.I0(x2091), .I1(x2092), .I2(x2093), .I3(n10914), .I4(n10915), .O(n10918));
  LUT5 #(.INIT(32'hFF969600)) lut_n10919 (.I0(x2097), .I1(x2098), .I2(x2099), .I3(n10917), .I4(n10918), .O(n10919));
  LUT3 #(.INIT(8'h96)) lut_n10920 (.I0(n10904), .I1(n10907), .I2(n10908), .O(n10920));
  LUT3 #(.INIT(8'hE8)) lut_n10921 (.I0(n10916), .I1(n10919), .I2(n10920), .O(n10921));
  LUT3 #(.INIT(8'h96)) lut_n10922 (.I0(x2106), .I1(x2107), .I2(x2108), .O(n10922));
  LUT5 #(.INIT(32'h96696996)) lut_n10923 (.I0(x2097), .I1(x2098), .I2(x2099), .I3(n10917), .I4(n10918), .O(n10923));
  LUT5 #(.INIT(32'hFF969600)) lut_n10924 (.I0(x2103), .I1(x2104), .I2(x2105), .I3(n10922), .I4(n10923), .O(n10924));
  LUT3 #(.INIT(8'h96)) lut_n10925 (.I0(x2112), .I1(x2113), .I2(x2114), .O(n10925));
  LUT5 #(.INIT(32'h96696996)) lut_n10926 (.I0(x2103), .I1(x2104), .I2(x2105), .I3(n10922), .I4(n10923), .O(n10926));
  LUT5 #(.INIT(32'hFF969600)) lut_n10927 (.I0(x2109), .I1(x2110), .I2(x2111), .I3(n10925), .I4(n10926), .O(n10927));
  LUT3 #(.INIT(8'h96)) lut_n10928 (.I0(n10916), .I1(n10919), .I2(n10920), .O(n10928));
  LUT3 #(.INIT(8'hE8)) lut_n10929 (.I0(n10924), .I1(n10927), .I2(n10928), .O(n10929));
  LUT3 #(.INIT(8'h96)) lut_n10930 (.I0(n10901), .I1(n10909), .I2(n10910), .O(n10930));
  LUT3 #(.INIT(8'hE8)) lut_n10931 (.I0(n10921), .I1(n10929), .I2(n10930), .O(n10931));
  LUT3 #(.INIT(8'h96)) lut_n10932 (.I0(x2118), .I1(x2119), .I2(x2120), .O(n10932));
  LUT5 #(.INIT(32'h96696996)) lut_n10933 (.I0(x2109), .I1(x2110), .I2(x2111), .I3(n10925), .I4(n10926), .O(n10933));
  LUT5 #(.INIT(32'hFF969600)) lut_n10934 (.I0(x2115), .I1(x2116), .I2(x2117), .I3(n10932), .I4(n10933), .O(n10934));
  LUT3 #(.INIT(8'h96)) lut_n10935 (.I0(x2124), .I1(x2125), .I2(x2126), .O(n10935));
  LUT5 #(.INIT(32'h96696996)) lut_n10936 (.I0(x2115), .I1(x2116), .I2(x2117), .I3(n10932), .I4(n10933), .O(n10936));
  LUT5 #(.INIT(32'hFF969600)) lut_n10937 (.I0(x2121), .I1(x2122), .I2(x2123), .I3(n10935), .I4(n10936), .O(n10937));
  LUT3 #(.INIT(8'h96)) lut_n10938 (.I0(n10924), .I1(n10927), .I2(n10928), .O(n10938));
  LUT3 #(.INIT(8'hE8)) lut_n10939 (.I0(n10934), .I1(n10937), .I2(n10938), .O(n10939));
  LUT3 #(.INIT(8'h96)) lut_n10940 (.I0(x2130), .I1(x2131), .I2(x2132), .O(n10940));
  LUT5 #(.INIT(32'h96696996)) lut_n10941 (.I0(x2121), .I1(x2122), .I2(x2123), .I3(n10935), .I4(n10936), .O(n10941));
  LUT5 #(.INIT(32'hFF969600)) lut_n10942 (.I0(x2127), .I1(x2128), .I2(x2129), .I3(n10940), .I4(n10941), .O(n10942));
  LUT3 #(.INIT(8'h96)) lut_n10943 (.I0(x2136), .I1(x2137), .I2(x2138), .O(n10943));
  LUT5 #(.INIT(32'h96696996)) lut_n10944 (.I0(x2127), .I1(x2128), .I2(x2129), .I3(n10940), .I4(n10941), .O(n10944));
  LUT5 #(.INIT(32'hFF969600)) lut_n10945 (.I0(x2133), .I1(x2134), .I2(x2135), .I3(n10943), .I4(n10944), .O(n10945));
  LUT3 #(.INIT(8'h96)) lut_n10946 (.I0(n10934), .I1(n10937), .I2(n10938), .O(n10946));
  LUT3 #(.INIT(8'hE8)) lut_n10947 (.I0(n10942), .I1(n10945), .I2(n10946), .O(n10947));
  LUT3 #(.INIT(8'h96)) lut_n10948 (.I0(n10921), .I1(n10929), .I2(n10930), .O(n10948));
  LUT3 #(.INIT(8'hE8)) lut_n10949 (.I0(n10939), .I1(n10947), .I2(n10948), .O(n10949));
  LUT3 #(.INIT(8'h96)) lut_n10950 (.I0(n10893), .I1(n10911), .I2(n10912), .O(n10950));
  LUT3 #(.INIT(8'hE8)) lut_n10951 (.I0(n10931), .I1(n10949), .I2(n10950), .O(n10951));
  LUT3 #(.INIT(8'h96)) lut_n10952 (.I0(n10833), .I1(n10871), .I2(n10872), .O(n10952));
  LUT3 #(.INIT(8'hE8)) lut_n10953 (.I0(n10913), .I1(n10951), .I2(n10952), .O(n10953));
  LUT3 #(.INIT(8'h96)) lut_n10954 (.I0(x2142), .I1(x2143), .I2(x2144), .O(n10954));
  LUT5 #(.INIT(32'h96696996)) lut_n10955 (.I0(x2133), .I1(x2134), .I2(x2135), .I3(n10943), .I4(n10944), .O(n10955));
  LUT5 #(.INIT(32'hFF969600)) lut_n10956 (.I0(x2139), .I1(x2140), .I2(x2141), .I3(n10954), .I4(n10955), .O(n10956));
  LUT3 #(.INIT(8'h96)) lut_n10957 (.I0(x2148), .I1(x2149), .I2(x2150), .O(n10957));
  LUT5 #(.INIT(32'h96696996)) lut_n10958 (.I0(x2139), .I1(x2140), .I2(x2141), .I3(n10954), .I4(n10955), .O(n10958));
  LUT5 #(.INIT(32'hFF969600)) lut_n10959 (.I0(x2145), .I1(x2146), .I2(x2147), .I3(n10957), .I4(n10958), .O(n10959));
  LUT3 #(.INIT(8'h96)) lut_n10960 (.I0(n10942), .I1(n10945), .I2(n10946), .O(n10960));
  LUT3 #(.INIT(8'hE8)) lut_n10961 (.I0(n10956), .I1(n10959), .I2(n10960), .O(n10961));
  LUT3 #(.INIT(8'h96)) lut_n10962 (.I0(x2154), .I1(x2155), .I2(x2156), .O(n10962));
  LUT5 #(.INIT(32'h96696996)) lut_n10963 (.I0(x2145), .I1(x2146), .I2(x2147), .I3(n10957), .I4(n10958), .O(n10963));
  LUT5 #(.INIT(32'hFF969600)) lut_n10964 (.I0(x2151), .I1(x2152), .I2(x2153), .I3(n10962), .I4(n10963), .O(n10964));
  LUT3 #(.INIT(8'h96)) lut_n10965 (.I0(x2160), .I1(x2161), .I2(x2162), .O(n10965));
  LUT5 #(.INIT(32'h96696996)) lut_n10966 (.I0(x2151), .I1(x2152), .I2(x2153), .I3(n10962), .I4(n10963), .O(n10966));
  LUT5 #(.INIT(32'hFF969600)) lut_n10967 (.I0(x2157), .I1(x2158), .I2(x2159), .I3(n10965), .I4(n10966), .O(n10967));
  LUT3 #(.INIT(8'h96)) lut_n10968 (.I0(n10956), .I1(n10959), .I2(n10960), .O(n10968));
  LUT3 #(.INIT(8'hE8)) lut_n10969 (.I0(n10964), .I1(n10967), .I2(n10968), .O(n10969));
  LUT3 #(.INIT(8'h96)) lut_n10970 (.I0(n10939), .I1(n10947), .I2(n10948), .O(n10970));
  LUT3 #(.INIT(8'hE8)) lut_n10971 (.I0(n10961), .I1(n10969), .I2(n10970), .O(n10971));
  LUT3 #(.INIT(8'h96)) lut_n10972 (.I0(x2166), .I1(x2167), .I2(x2168), .O(n10972));
  LUT5 #(.INIT(32'h96696996)) lut_n10973 (.I0(x2157), .I1(x2158), .I2(x2159), .I3(n10965), .I4(n10966), .O(n10973));
  LUT5 #(.INIT(32'hFF969600)) lut_n10974 (.I0(x2163), .I1(x2164), .I2(x2165), .I3(n10972), .I4(n10973), .O(n10974));
  LUT3 #(.INIT(8'h96)) lut_n10975 (.I0(x2172), .I1(x2173), .I2(x2174), .O(n10975));
  LUT5 #(.INIT(32'h96696996)) lut_n10976 (.I0(x2163), .I1(x2164), .I2(x2165), .I3(n10972), .I4(n10973), .O(n10976));
  LUT5 #(.INIT(32'hFF969600)) lut_n10977 (.I0(x2169), .I1(x2170), .I2(x2171), .I3(n10975), .I4(n10976), .O(n10977));
  LUT3 #(.INIT(8'h96)) lut_n10978 (.I0(n10964), .I1(n10967), .I2(n10968), .O(n10978));
  LUT3 #(.INIT(8'hE8)) lut_n10979 (.I0(n10974), .I1(n10977), .I2(n10978), .O(n10979));
  LUT3 #(.INIT(8'h96)) lut_n10980 (.I0(x2178), .I1(x2179), .I2(x2180), .O(n10980));
  LUT5 #(.INIT(32'h96696996)) lut_n10981 (.I0(x2169), .I1(x2170), .I2(x2171), .I3(n10975), .I4(n10976), .O(n10981));
  LUT5 #(.INIT(32'hFF969600)) lut_n10982 (.I0(x2175), .I1(x2176), .I2(x2177), .I3(n10980), .I4(n10981), .O(n10982));
  LUT3 #(.INIT(8'h96)) lut_n10983 (.I0(x2184), .I1(x2185), .I2(x2186), .O(n10983));
  LUT5 #(.INIT(32'h96696996)) lut_n10984 (.I0(x2175), .I1(x2176), .I2(x2177), .I3(n10980), .I4(n10981), .O(n10984));
  LUT5 #(.INIT(32'hFF969600)) lut_n10985 (.I0(x2181), .I1(x2182), .I2(x2183), .I3(n10983), .I4(n10984), .O(n10985));
  LUT3 #(.INIT(8'h96)) lut_n10986 (.I0(n10974), .I1(n10977), .I2(n10978), .O(n10986));
  LUT3 #(.INIT(8'hE8)) lut_n10987 (.I0(n10982), .I1(n10985), .I2(n10986), .O(n10987));
  LUT3 #(.INIT(8'h96)) lut_n10988 (.I0(n10961), .I1(n10969), .I2(n10970), .O(n10988));
  LUT3 #(.INIT(8'hE8)) lut_n10989 (.I0(n10979), .I1(n10987), .I2(n10988), .O(n10989));
  LUT3 #(.INIT(8'h96)) lut_n10990 (.I0(n10931), .I1(n10949), .I2(n10950), .O(n10990));
  LUT3 #(.INIT(8'hE8)) lut_n10991 (.I0(n10971), .I1(n10989), .I2(n10990), .O(n10991));
  LUT3 #(.INIT(8'h96)) lut_n10992 (.I0(x2190), .I1(x2191), .I2(x2192), .O(n10992));
  LUT5 #(.INIT(32'h96696996)) lut_n10993 (.I0(x2181), .I1(x2182), .I2(x2183), .I3(n10983), .I4(n10984), .O(n10993));
  LUT5 #(.INIT(32'hFF969600)) lut_n10994 (.I0(x2187), .I1(x2188), .I2(x2189), .I3(n10992), .I4(n10993), .O(n10994));
  LUT3 #(.INIT(8'h96)) lut_n10995 (.I0(x2196), .I1(x2197), .I2(x2198), .O(n10995));
  LUT5 #(.INIT(32'h96696996)) lut_n10996 (.I0(x2187), .I1(x2188), .I2(x2189), .I3(n10992), .I4(n10993), .O(n10996));
  LUT5 #(.INIT(32'hFF969600)) lut_n10997 (.I0(x2193), .I1(x2194), .I2(x2195), .I3(n10995), .I4(n10996), .O(n10997));
  LUT3 #(.INIT(8'h96)) lut_n10998 (.I0(n10982), .I1(n10985), .I2(n10986), .O(n10998));
  LUT3 #(.INIT(8'hE8)) lut_n10999 (.I0(n10994), .I1(n10997), .I2(n10998), .O(n10999));
  LUT3 #(.INIT(8'h96)) lut_n11000 (.I0(x2202), .I1(x2203), .I2(x2204), .O(n11000));
  LUT5 #(.INIT(32'h96696996)) lut_n11001 (.I0(x2193), .I1(x2194), .I2(x2195), .I3(n10995), .I4(n10996), .O(n11001));
  LUT5 #(.INIT(32'hFF969600)) lut_n11002 (.I0(x2199), .I1(x2200), .I2(x2201), .I3(n11000), .I4(n11001), .O(n11002));
  LUT3 #(.INIT(8'h96)) lut_n11003 (.I0(x2208), .I1(x2209), .I2(x2210), .O(n11003));
  LUT5 #(.INIT(32'h96696996)) lut_n11004 (.I0(x2199), .I1(x2200), .I2(x2201), .I3(n11000), .I4(n11001), .O(n11004));
  LUT5 #(.INIT(32'hFF969600)) lut_n11005 (.I0(x2205), .I1(x2206), .I2(x2207), .I3(n11003), .I4(n11004), .O(n11005));
  LUT3 #(.INIT(8'h96)) lut_n11006 (.I0(n10994), .I1(n10997), .I2(n10998), .O(n11006));
  LUT3 #(.INIT(8'hE8)) lut_n11007 (.I0(n11002), .I1(n11005), .I2(n11006), .O(n11007));
  LUT3 #(.INIT(8'h96)) lut_n11008 (.I0(n10979), .I1(n10987), .I2(n10988), .O(n11008));
  LUT3 #(.INIT(8'hE8)) lut_n11009 (.I0(n10999), .I1(n11007), .I2(n11008), .O(n11009));
  LUT3 #(.INIT(8'h96)) lut_n11010 (.I0(x2214), .I1(x2215), .I2(x2216), .O(n11010));
  LUT5 #(.INIT(32'h96696996)) lut_n11011 (.I0(x2205), .I1(x2206), .I2(x2207), .I3(n11003), .I4(n11004), .O(n11011));
  LUT5 #(.INIT(32'hFF969600)) lut_n11012 (.I0(x2211), .I1(x2212), .I2(x2213), .I3(n11010), .I4(n11011), .O(n11012));
  LUT3 #(.INIT(8'h96)) lut_n11013 (.I0(x2220), .I1(x2221), .I2(x2222), .O(n11013));
  LUT5 #(.INIT(32'h96696996)) lut_n11014 (.I0(x2211), .I1(x2212), .I2(x2213), .I3(n11010), .I4(n11011), .O(n11014));
  LUT5 #(.INIT(32'hFF969600)) lut_n11015 (.I0(x2217), .I1(x2218), .I2(x2219), .I3(n11013), .I4(n11014), .O(n11015));
  LUT3 #(.INIT(8'h96)) lut_n11016 (.I0(n11002), .I1(n11005), .I2(n11006), .O(n11016));
  LUT3 #(.INIT(8'hE8)) lut_n11017 (.I0(n11012), .I1(n11015), .I2(n11016), .O(n11017));
  LUT3 #(.INIT(8'h96)) lut_n11018 (.I0(x2226), .I1(x2227), .I2(x2228), .O(n11018));
  LUT5 #(.INIT(32'h96696996)) lut_n11019 (.I0(x2217), .I1(x2218), .I2(x2219), .I3(n11013), .I4(n11014), .O(n11019));
  LUT5 #(.INIT(32'hFF969600)) lut_n11020 (.I0(x2223), .I1(x2224), .I2(x2225), .I3(n11018), .I4(n11019), .O(n11020));
  LUT3 #(.INIT(8'h96)) lut_n11021 (.I0(x2232), .I1(x2233), .I2(x2234), .O(n11021));
  LUT5 #(.INIT(32'h96696996)) lut_n11022 (.I0(x2223), .I1(x2224), .I2(x2225), .I3(n11018), .I4(n11019), .O(n11022));
  LUT5 #(.INIT(32'hFF969600)) lut_n11023 (.I0(x2229), .I1(x2230), .I2(x2231), .I3(n11021), .I4(n11022), .O(n11023));
  LUT3 #(.INIT(8'h96)) lut_n11024 (.I0(n11012), .I1(n11015), .I2(n11016), .O(n11024));
  LUT3 #(.INIT(8'hE8)) lut_n11025 (.I0(n11020), .I1(n11023), .I2(n11024), .O(n11025));
  LUT3 #(.INIT(8'h96)) lut_n11026 (.I0(n10999), .I1(n11007), .I2(n11008), .O(n11026));
  LUT3 #(.INIT(8'hE8)) lut_n11027 (.I0(n11017), .I1(n11025), .I2(n11026), .O(n11027));
  LUT3 #(.INIT(8'h96)) lut_n11028 (.I0(n10971), .I1(n10989), .I2(n10990), .O(n11028));
  LUT3 #(.INIT(8'hE8)) lut_n11029 (.I0(n11009), .I1(n11027), .I2(n11028), .O(n11029));
  LUT3 #(.INIT(8'h96)) lut_n11030 (.I0(n10913), .I1(n10951), .I2(n10952), .O(n11030));
  LUT3 #(.INIT(8'hE8)) lut_n11031 (.I0(n10991), .I1(n11029), .I2(n11030), .O(n11031));
  LUT3 #(.INIT(8'h96)) lut_n11032 (.I0(n10795), .I1(n10873), .I2(n10874), .O(n11032));
  LUT3 #(.INIT(8'hE8)) lut_n11033 (.I0(n10953), .I1(n11031), .I2(n11032), .O(n11033));
  LUT3 #(.INIT(8'h96)) lut_n11034 (.I0(n10557), .I1(n10715), .I2(n10716), .O(n11034));
  LUT3 #(.INIT(8'hE8)) lut_n11035 (.I0(n10875), .I1(n11033), .I2(n11034), .O(n11035));
  LUT3 #(.INIT(8'h96)) lut_n11036 (.I0(n10079), .I1(n10397), .I2(n10398), .O(n11036));
  LUT3 #(.INIT(8'hE8)) lut_n11037 (.I0(n10717), .I1(n11035), .I2(n11036), .O(n11037));
  LUT3 #(.INIT(8'h96)) lut_n11038 (.I0(n9151), .I1(n9759), .I2(n9760), .O(n11038));
  LUT3 #(.INIT(8'hE8)) lut_n11039 (.I0(n10399), .I1(n11037), .I2(n11038), .O(n11039));
  LUT3 #(.INIT(8'h96)) lut_n11040 (.I0(n8193), .I1(n8831), .I2(n8832), .O(n11040));
  LUT3 #(.INIT(8'hE8)) lut_n11041 (.I0(n9761), .I1(n11039), .I2(n11040), .O(n11041));
  LUT3 #(.INIT(8'hE8)) lut_n11042 (.I0(n7555), .I1(n8833), .I2(n11041), .O(n11042));
  LUT3 #(.INIT(8'h96)) lut_n11043 (.I0(x2238), .I1(x2239), .I2(x2240), .O(n11043));
  LUT5 #(.INIT(32'h96696996)) lut_n11044 (.I0(x2229), .I1(x2230), .I2(x2231), .I3(n11021), .I4(n11022), .O(n11044));
  LUT5 #(.INIT(32'hFF969600)) lut_n11045 (.I0(x2235), .I1(x2236), .I2(x2237), .I3(n11043), .I4(n11044), .O(n11045));
  LUT3 #(.INIT(8'h96)) lut_n11046 (.I0(x2244), .I1(x2245), .I2(x2246), .O(n11046));
  LUT5 #(.INIT(32'h96696996)) lut_n11047 (.I0(x2235), .I1(x2236), .I2(x2237), .I3(n11043), .I4(n11044), .O(n11047));
  LUT5 #(.INIT(32'hFF969600)) lut_n11048 (.I0(x2241), .I1(x2242), .I2(x2243), .I3(n11046), .I4(n11047), .O(n11048));
  LUT3 #(.INIT(8'h96)) lut_n11049 (.I0(n11020), .I1(n11023), .I2(n11024), .O(n11049));
  LUT3 #(.INIT(8'hE8)) lut_n11050 (.I0(n11045), .I1(n11048), .I2(n11049), .O(n11050));
  LUT3 #(.INIT(8'h96)) lut_n11051 (.I0(x2250), .I1(x2251), .I2(x2252), .O(n11051));
  LUT5 #(.INIT(32'h96696996)) lut_n11052 (.I0(x2241), .I1(x2242), .I2(x2243), .I3(n11046), .I4(n11047), .O(n11052));
  LUT5 #(.INIT(32'hFF969600)) lut_n11053 (.I0(x2247), .I1(x2248), .I2(x2249), .I3(n11051), .I4(n11052), .O(n11053));
  LUT3 #(.INIT(8'h96)) lut_n11054 (.I0(x2256), .I1(x2257), .I2(x2258), .O(n11054));
  LUT5 #(.INIT(32'h96696996)) lut_n11055 (.I0(x2247), .I1(x2248), .I2(x2249), .I3(n11051), .I4(n11052), .O(n11055));
  LUT5 #(.INIT(32'hFF969600)) lut_n11056 (.I0(x2253), .I1(x2254), .I2(x2255), .I3(n11054), .I4(n11055), .O(n11056));
  LUT3 #(.INIT(8'h96)) lut_n11057 (.I0(n11045), .I1(n11048), .I2(n11049), .O(n11057));
  LUT3 #(.INIT(8'hE8)) lut_n11058 (.I0(n11053), .I1(n11056), .I2(n11057), .O(n11058));
  LUT3 #(.INIT(8'h96)) lut_n11059 (.I0(n11017), .I1(n11025), .I2(n11026), .O(n11059));
  LUT3 #(.INIT(8'hE8)) lut_n11060 (.I0(n11050), .I1(n11058), .I2(n11059), .O(n11060));
  LUT3 #(.INIT(8'h96)) lut_n11061 (.I0(x2262), .I1(x2263), .I2(x2264), .O(n11061));
  LUT5 #(.INIT(32'h96696996)) lut_n11062 (.I0(x2253), .I1(x2254), .I2(x2255), .I3(n11054), .I4(n11055), .O(n11062));
  LUT5 #(.INIT(32'hFF969600)) lut_n11063 (.I0(x2259), .I1(x2260), .I2(x2261), .I3(n11061), .I4(n11062), .O(n11063));
  LUT3 #(.INIT(8'h96)) lut_n11064 (.I0(x2268), .I1(x2269), .I2(x2270), .O(n11064));
  LUT5 #(.INIT(32'h96696996)) lut_n11065 (.I0(x2259), .I1(x2260), .I2(x2261), .I3(n11061), .I4(n11062), .O(n11065));
  LUT5 #(.INIT(32'hFF969600)) lut_n11066 (.I0(x2265), .I1(x2266), .I2(x2267), .I3(n11064), .I4(n11065), .O(n11066));
  LUT3 #(.INIT(8'h96)) lut_n11067 (.I0(n11053), .I1(n11056), .I2(n11057), .O(n11067));
  LUT3 #(.INIT(8'hE8)) lut_n11068 (.I0(n11063), .I1(n11066), .I2(n11067), .O(n11068));
  LUT3 #(.INIT(8'h96)) lut_n11069 (.I0(x2274), .I1(x2275), .I2(x2276), .O(n11069));
  LUT5 #(.INIT(32'h96696996)) lut_n11070 (.I0(x2265), .I1(x2266), .I2(x2267), .I3(n11064), .I4(n11065), .O(n11070));
  LUT5 #(.INIT(32'hFF969600)) lut_n11071 (.I0(x2271), .I1(x2272), .I2(x2273), .I3(n11069), .I4(n11070), .O(n11071));
  LUT3 #(.INIT(8'h96)) lut_n11072 (.I0(x2280), .I1(x2281), .I2(x2282), .O(n11072));
  LUT5 #(.INIT(32'h96696996)) lut_n11073 (.I0(x2271), .I1(x2272), .I2(x2273), .I3(n11069), .I4(n11070), .O(n11073));
  LUT5 #(.INIT(32'hFF969600)) lut_n11074 (.I0(x2277), .I1(x2278), .I2(x2279), .I3(n11072), .I4(n11073), .O(n11074));
  LUT3 #(.INIT(8'h96)) lut_n11075 (.I0(n11063), .I1(n11066), .I2(n11067), .O(n11075));
  LUT3 #(.INIT(8'hE8)) lut_n11076 (.I0(n11071), .I1(n11074), .I2(n11075), .O(n11076));
  LUT3 #(.INIT(8'h96)) lut_n11077 (.I0(n11050), .I1(n11058), .I2(n11059), .O(n11077));
  LUT3 #(.INIT(8'hE8)) lut_n11078 (.I0(n11068), .I1(n11076), .I2(n11077), .O(n11078));
  LUT3 #(.INIT(8'h96)) lut_n11079 (.I0(n11009), .I1(n11027), .I2(n11028), .O(n11079));
  LUT3 #(.INIT(8'hE8)) lut_n11080 (.I0(n11060), .I1(n11078), .I2(n11079), .O(n11080));
  LUT3 #(.INIT(8'h96)) lut_n11081 (.I0(x2286), .I1(x2287), .I2(x2288), .O(n11081));
  LUT5 #(.INIT(32'h96696996)) lut_n11082 (.I0(x2277), .I1(x2278), .I2(x2279), .I3(n11072), .I4(n11073), .O(n11082));
  LUT5 #(.INIT(32'hFF969600)) lut_n11083 (.I0(x2283), .I1(x2284), .I2(x2285), .I3(n11081), .I4(n11082), .O(n11083));
  LUT3 #(.INIT(8'h96)) lut_n11084 (.I0(x2292), .I1(x2293), .I2(x2294), .O(n11084));
  LUT5 #(.INIT(32'h96696996)) lut_n11085 (.I0(x2283), .I1(x2284), .I2(x2285), .I3(n11081), .I4(n11082), .O(n11085));
  LUT5 #(.INIT(32'hFF969600)) lut_n11086 (.I0(x2289), .I1(x2290), .I2(x2291), .I3(n11084), .I4(n11085), .O(n11086));
  LUT3 #(.INIT(8'h96)) lut_n11087 (.I0(n11071), .I1(n11074), .I2(n11075), .O(n11087));
  LUT3 #(.INIT(8'hE8)) lut_n11088 (.I0(n11083), .I1(n11086), .I2(n11087), .O(n11088));
  LUT3 #(.INIT(8'h96)) lut_n11089 (.I0(x2298), .I1(x2299), .I2(x2300), .O(n11089));
  LUT5 #(.INIT(32'h96696996)) lut_n11090 (.I0(x2289), .I1(x2290), .I2(x2291), .I3(n11084), .I4(n11085), .O(n11090));
  LUT5 #(.INIT(32'hFF969600)) lut_n11091 (.I0(x2295), .I1(x2296), .I2(x2297), .I3(n11089), .I4(n11090), .O(n11091));
  LUT3 #(.INIT(8'h96)) lut_n11092 (.I0(x2304), .I1(x2305), .I2(x2306), .O(n11092));
  LUT5 #(.INIT(32'h96696996)) lut_n11093 (.I0(x2295), .I1(x2296), .I2(x2297), .I3(n11089), .I4(n11090), .O(n11093));
  LUT5 #(.INIT(32'hFF969600)) lut_n11094 (.I0(x2301), .I1(x2302), .I2(x2303), .I3(n11092), .I4(n11093), .O(n11094));
  LUT3 #(.INIT(8'h96)) lut_n11095 (.I0(n11083), .I1(n11086), .I2(n11087), .O(n11095));
  LUT3 #(.INIT(8'hE8)) lut_n11096 (.I0(n11091), .I1(n11094), .I2(n11095), .O(n11096));
  LUT3 #(.INIT(8'h96)) lut_n11097 (.I0(n11068), .I1(n11076), .I2(n11077), .O(n11097));
  LUT3 #(.INIT(8'hE8)) lut_n11098 (.I0(n11088), .I1(n11096), .I2(n11097), .O(n11098));
  LUT3 #(.INIT(8'h96)) lut_n11099 (.I0(x2310), .I1(x2311), .I2(x2312), .O(n11099));
  LUT5 #(.INIT(32'h96696996)) lut_n11100 (.I0(x2301), .I1(x2302), .I2(x2303), .I3(n11092), .I4(n11093), .O(n11100));
  LUT5 #(.INIT(32'hFF969600)) lut_n11101 (.I0(x2307), .I1(x2308), .I2(x2309), .I3(n11099), .I4(n11100), .O(n11101));
  LUT3 #(.INIT(8'h96)) lut_n11102 (.I0(x2316), .I1(x2317), .I2(x2318), .O(n11102));
  LUT5 #(.INIT(32'h96696996)) lut_n11103 (.I0(x2307), .I1(x2308), .I2(x2309), .I3(n11099), .I4(n11100), .O(n11103));
  LUT5 #(.INIT(32'hFF969600)) lut_n11104 (.I0(x2313), .I1(x2314), .I2(x2315), .I3(n11102), .I4(n11103), .O(n11104));
  LUT3 #(.INIT(8'h96)) lut_n11105 (.I0(n11091), .I1(n11094), .I2(n11095), .O(n11105));
  LUT3 #(.INIT(8'hE8)) lut_n11106 (.I0(n11101), .I1(n11104), .I2(n11105), .O(n11106));
  LUT3 #(.INIT(8'h96)) lut_n11107 (.I0(x2322), .I1(x2323), .I2(x2324), .O(n11107));
  LUT5 #(.INIT(32'h96696996)) lut_n11108 (.I0(x2313), .I1(x2314), .I2(x2315), .I3(n11102), .I4(n11103), .O(n11108));
  LUT5 #(.INIT(32'hFF969600)) lut_n11109 (.I0(x2319), .I1(x2320), .I2(x2321), .I3(n11107), .I4(n11108), .O(n11109));
  LUT3 #(.INIT(8'h96)) lut_n11110 (.I0(x2328), .I1(x2329), .I2(x2330), .O(n11110));
  LUT5 #(.INIT(32'h96696996)) lut_n11111 (.I0(x2319), .I1(x2320), .I2(x2321), .I3(n11107), .I4(n11108), .O(n11111));
  LUT5 #(.INIT(32'hFF969600)) lut_n11112 (.I0(x2325), .I1(x2326), .I2(x2327), .I3(n11110), .I4(n11111), .O(n11112));
  LUT3 #(.INIT(8'h96)) lut_n11113 (.I0(n11101), .I1(n11104), .I2(n11105), .O(n11113));
  LUT3 #(.INIT(8'hE8)) lut_n11114 (.I0(n11109), .I1(n11112), .I2(n11113), .O(n11114));
  LUT3 #(.INIT(8'h96)) lut_n11115 (.I0(n11088), .I1(n11096), .I2(n11097), .O(n11115));
  LUT3 #(.INIT(8'hE8)) lut_n11116 (.I0(n11106), .I1(n11114), .I2(n11115), .O(n11116));
  LUT3 #(.INIT(8'h96)) lut_n11117 (.I0(n11060), .I1(n11078), .I2(n11079), .O(n11117));
  LUT3 #(.INIT(8'hE8)) lut_n11118 (.I0(n11098), .I1(n11116), .I2(n11117), .O(n11118));
  LUT3 #(.INIT(8'h96)) lut_n11119 (.I0(n10991), .I1(n11029), .I2(n11030), .O(n11119));
  LUT3 #(.INIT(8'hE8)) lut_n11120 (.I0(n11080), .I1(n11118), .I2(n11119), .O(n11120));
  LUT3 #(.INIT(8'h96)) lut_n11121 (.I0(x2334), .I1(x2335), .I2(x2336), .O(n11121));
  LUT5 #(.INIT(32'h96696996)) lut_n11122 (.I0(x2325), .I1(x2326), .I2(x2327), .I3(n11110), .I4(n11111), .O(n11122));
  LUT5 #(.INIT(32'hFF969600)) lut_n11123 (.I0(x2331), .I1(x2332), .I2(x2333), .I3(n11121), .I4(n11122), .O(n11123));
  LUT3 #(.INIT(8'h96)) lut_n11124 (.I0(x2340), .I1(x2341), .I2(x2342), .O(n11124));
  LUT5 #(.INIT(32'h96696996)) lut_n11125 (.I0(x2331), .I1(x2332), .I2(x2333), .I3(n11121), .I4(n11122), .O(n11125));
  LUT5 #(.INIT(32'hFF969600)) lut_n11126 (.I0(x2337), .I1(x2338), .I2(x2339), .I3(n11124), .I4(n11125), .O(n11126));
  LUT3 #(.INIT(8'h96)) lut_n11127 (.I0(n11109), .I1(n11112), .I2(n11113), .O(n11127));
  LUT3 #(.INIT(8'hE8)) lut_n11128 (.I0(n11123), .I1(n11126), .I2(n11127), .O(n11128));
  LUT3 #(.INIT(8'h96)) lut_n11129 (.I0(x2346), .I1(x2347), .I2(x2348), .O(n11129));
  LUT5 #(.INIT(32'h96696996)) lut_n11130 (.I0(x2337), .I1(x2338), .I2(x2339), .I3(n11124), .I4(n11125), .O(n11130));
  LUT5 #(.INIT(32'hFF969600)) lut_n11131 (.I0(x2343), .I1(x2344), .I2(x2345), .I3(n11129), .I4(n11130), .O(n11131));
  LUT3 #(.INIT(8'h96)) lut_n11132 (.I0(x2352), .I1(x2353), .I2(x2354), .O(n11132));
  LUT5 #(.INIT(32'h96696996)) lut_n11133 (.I0(x2343), .I1(x2344), .I2(x2345), .I3(n11129), .I4(n11130), .O(n11133));
  LUT5 #(.INIT(32'hFF969600)) lut_n11134 (.I0(x2349), .I1(x2350), .I2(x2351), .I3(n11132), .I4(n11133), .O(n11134));
  LUT3 #(.INIT(8'h96)) lut_n11135 (.I0(n11123), .I1(n11126), .I2(n11127), .O(n11135));
  LUT3 #(.INIT(8'hE8)) lut_n11136 (.I0(n11131), .I1(n11134), .I2(n11135), .O(n11136));
  LUT3 #(.INIT(8'h96)) lut_n11137 (.I0(n11106), .I1(n11114), .I2(n11115), .O(n11137));
  LUT3 #(.INIT(8'hE8)) lut_n11138 (.I0(n11128), .I1(n11136), .I2(n11137), .O(n11138));
  LUT3 #(.INIT(8'h96)) lut_n11139 (.I0(x2358), .I1(x2359), .I2(x2360), .O(n11139));
  LUT5 #(.INIT(32'h96696996)) lut_n11140 (.I0(x2349), .I1(x2350), .I2(x2351), .I3(n11132), .I4(n11133), .O(n11140));
  LUT5 #(.INIT(32'hFF969600)) lut_n11141 (.I0(x2355), .I1(x2356), .I2(x2357), .I3(n11139), .I4(n11140), .O(n11141));
  LUT3 #(.INIT(8'h96)) lut_n11142 (.I0(x2364), .I1(x2365), .I2(x2366), .O(n11142));
  LUT5 #(.INIT(32'h96696996)) lut_n11143 (.I0(x2355), .I1(x2356), .I2(x2357), .I3(n11139), .I4(n11140), .O(n11143));
  LUT5 #(.INIT(32'hFF969600)) lut_n11144 (.I0(x2361), .I1(x2362), .I2(x2363), .I3(n11142), .I4(n11143), .O(n11144));
  LUT3 #(.INIT(8'h96)) lut_n11145 (.I0(n11131), .I1(n11134), .I2(n11135), .O(n11145));
  LUT3 #(.INIT(8'hE8)) lut_n11146 (.I0(n11141), .I1(n11144), .I2(n11145), .O(n11146));
  LUT3 #(.INIT(8'h96)) lut_n11147 (.I0(x2370), .I1(x2371), .I2(x2372), .O(n11147));
  LUT5 #(.INIT(32'h96696996)) lut_n11148 (.I0(x2361), .I1(x2362), .I2(x2363), .I3(n11142), .I4(n11143), .O(n11148));
  LUT5 #(.INIT(32'hFF969600)) lut_n11149 (.I0(x2367), .I1(x2368), .I2(x2369), .I3(n11147), .I4(n11148), .O(n11149));
  LUT3 #(.INIT(8'h96)) lut_n11150 (.I0(x2376), .I1(x2377), .I2(x2378), .O(n11150));
  LUT5 #(.INIT(32'h96696996)) lut_n11151 (.I0(x2367), .I1(x2368), .I2(x2369), .I3(n11147), .I4(n11148), .O(n11151));
  LUT5 #(.INIT(32'hFF969600)) lut_n11152 (.I0(x2373), .I1(x2374), .I2(x2375), .I3(n11150), .I4(n11151), .O(n11152));
  LUT3 #(.INIT(8'h96)) lut_n11153 (.I0(n11141), .I1(n11144), .I2(n11145), .O(n11153));
  LUT3 #(.INIT(8'hE8)) lut_n11154 (.I0(n11149), .I1(n11152), .I2(n11153), .O(n11154));
  LUT3 #(.INIT(8'h96)) lut_n11155 (.I0(n11128), .I1(n11136), .I2(n11137), .O(n11155));
  LUT3 #(.INIT(8'hE8)) lut_n11156 (.I0(n11146), .I1(n11154), .I2(n11155), .O(n11156));
  LUT3 #(.INIT(8'h96)) lut_n11157 (.I0(n11098), .I1(n11116), .I2(n11117), .O(n11157));
  LUT3 #(.INIT(8'hE8)) lut_n11158 (.I0(n11138), .I1(n11156), .I2(n11157), .O(n11158));
  LUT3 #(.INIT(8'h96)) lut_n11159 (.I0(x2382), .I1(x2383), .I2(x2384), .O(n11159));
  LUT5 #(.INIT(32'h96696996)) lut_n11160 (.I0(x2373), .I1(x2374), .I2(x2375), .I3(n11150), .I4(n11151), .O(n11160));
  LUT5 #(.INIT(32'hFF969600)) lut_n11161 (.I0(x2379), .I1(x2380), .I2(x2381), .I3(n11159), .I4(n11160), .O(n11161));
  LUT3 #(.INIT(8'h96)) lut_n11162 (.I0(x2388), .I1(x2389), .I2(x2390), .O(n11162));
  LUT5 #(.INIT(32'h96696996)) lut_n11163 (.I0(x2379), .I1(x2380), .I2(x2381), .I3(n11159), .I4(n11160), .O(n11163));
  LUT5 #(.INIT(32'hFF969600)) lut_n11164 (.I0(x2385), .I1(x2386), .I2(x2387), .I3(n11162), .I4(n11163), .O(n11164));
  LUT3 #(.INIT(8'h96)) lut_n11165 (.I0(n11149), .I1(n11152), .I2(n11153), .O(n11165));
  LUT3 #(.INIT(8'hE8)) lut_n11166 (.I0(n11161), .I1(n11164), .I2(n11165), .O(n11166));
  LUT3 #(.INIT(8'h96)) lut_n11167 (.I0(x2394), .I1(x2395), .I2(x2396), .O(n11167));
  LUT5 #(.INIT(32'h96696996)) lut_n11168 (.I0(x2385), .I1(x2386), .I2(x2387), .I3(n11162), .I4(n11163), .O(n11168));
  LUT5 #(.INIT(32'hFF969600)) lut_n11169 (.I0(x2391), .I1(x2392), .I2(x2393), .I3(n11167), .I4(n11168), .O(n11169));
  LUT3 #(.INIT(8'h96)) lut_n11170 (.I0(x2400), .I1(x2401), .I2(x2402), .O(n11170));
  LUT5 #(.INIT(32'h96696996)) lut_n11171 (.I0(x2391), .I1(x2392), .I2(x2393), .I3(n11167), .I4(n11168), .O(n11171));
  LUT5 #(.INIT(32'hFF969600)) lut_n11172 (.I0(x2397), .I1(x2398), .I2(x2399), .I3(n11170), .I4(n11171), .O(n11172));
  LUT3 #(.INIT(8'h96)) lut_n11173 (.I0(n11161), .I1(n11164), .I2(n11165), .O(n11173));
  LUT3 #(.INIT(8'hE8)) lut_n11174 (.I0(n11169), .I1(n11172), .I2(n11173), .O(n11174));
  LUT3 #(.INIT(8'h96)) lut_n11175 (.I0(n11146), .I1(n11154), .I2(n11155), .O(n11175));
  LUT3 #(.INIT(8'hE8)) lut_n11176 (.I0(n11166), .I1(n11174), .I2(n11175), .O(n11176));
  LUT3 #(.INIT(8'h96)) lut_n11177 (.I0(x2406), .I1(x2407), .I2(x2408), .O(n11177));
  LUT5 #(.INIT(32'h96696996)) lut_n11178 (.I0(x2397), .I1(x2398), .I2(x2399), .I3(n11170), .I4(n11171), .O(n11178));
  LUT5 #(.INIT(32'hFF969600)) lut_n11179 (.I0(x2403), .I1(x2404), .I2(x2405), .I3(n11177), .I4(n11178), .O(n11179));
  LUT3 #(.INIT(8'h96)) lut_n11180 (.I0(x2412), .I1(x2413), .I2(x2414), .O(n11180));
  LUT5 #(.INIT(32'h96696996)) lut_n11181 (.I0(x2403), .I1(x2404), .I2(x2405), .I3(n11177), .I4(n11178), .O(n11181));
  LUT5 #(.INIT(32'hFF969600)) lut_n11182 (.I0(x2409), .I1(x2410), .I2(x2411), .I3(n11180), .I4(n11181), .O(n11182));
  LUT3 #(.INIT(8'h96)) lut_n11183 (.I0(n11169), .I1(n11172), .I2(n11173), .O(n11183));
  LUT3 #(.INIT(8'hE8)) lut_n11184 (.I0(n11179), .I1(n11182), .I2(n11183), .O(n11184));
  LUT3 #(.INIT(8'h96)) lut_n11185 (.I0(x2418), .I1(x2419), .I2(x2420), .O(n11185));
  LUT5 #(.INIT(32'h96696996)) lut_n11186 (.I0(x2409), .I1(x2410), .I2(x2411), .I3(n11180), .I4(n11181), .O(n11186));
  LUT5 #(.INIT(32'hFF969600)) lut_n11187 (.I0(x2415), .I1(x2416), .I2(x2417), .I3(n11185), .I4(n11186), .O(n11187));
  LUT3 #(.INIT(8'h96)) lut_n11188 (.I0(x2424), .I1(x2425), .I2(x2426), .O(n11188));
  LUT5 #(.INIT(32'h96696996)) lut_n11189 (.I0(x2415), .I1(x2416), .I2(x2417), .I3(n11185), .I4(n11186), .O(n11189));
  LUT5 #(.INIT(32'hFF969600)) lut_n11190 (.I0(x2421), .I1(x2422), .I2(x2423), .I3(n11188), .I4(n11189), .O(n11190));
  LUT3 #(.INIT(8'h96)) lut_n11191 (.I0(n11179), .I1(n11182), .I2(n11183), .O(n11191));
  LUT3 #(.INIT(8'hE8)) lut_n11192 (.I0(n11187), .I1(n11190), .I2(n11191), .O(n11192));
  LUT3 #(.INIT(8'h96)) lut_n11193 (.I0(n11166), .I1(n11174), .I2(n11175), .O(n11193));
  LUT3 #(.INIT(8'hE8)) lut_n11194 (.I0(n11184), .I1(n11192), .I2(n11193), .O(n11194));
  LUT3 #(.INIT(8'h96)) lut_n11195 (.I0(n11138), .I1(n11156), .I2(n11157), .O(n11195));
  LUT3 #(.INIT(8'hE8)) lut_n11196 (.I0(n11176), .I1(n11194), .I2(n11195), .O(n11196));
  LUT3 #(.INIT(8'h96)) lut_n11197 (.I0(n11080), .I1(n11118), .I2(n11119), .O(n11197));
  LUT3 #(.INIT(8'hE8)) lut_n11198 (.I0(n11158), .I1(n11196), .I2(n11197), .O(n11198));
  LUT3 #(.INIT(8'h96)) lut_n11199 (.I0(n10953), .I1(n11031), .I2(n11032), .O(n11199));
  LUT3 #(.INIT(8'hE8)) lut_n11200 (.I0(n11120), .I1(n11198), .I2(n11199), .O(n11200));
  LUT3 #(.INIT(8'h96)) lut_n11201 (.I0(x2430), .I1(x2431), .I2(x2432), .O(n11201));
  LUT5 #(.INIT(32'h96696996)) lut_n11202 (.I0(x2421), .I1(x2422), .I2(x2423), .I3(n11188), .I4(n11189), .O(n11202));
  LUT5 #(.INIT(32'hFF969600)) lut_n11203 (.I0(x2427), .I1(x2428), .I2(x2429), .I3(n11201), .I4(n11202), .O(n11203));
  LUT3 #(.INIT(8'h96)) lut_n11204 (.I0(x2436), .I1(x2437), .I2(x2438), .O(n11204));
  LUT5 #(.INIT(32'h96696996)) lut_n11205 (.I0(x2427), .I1(x2428), .I2(x2429), .I3(n11201), .I4(n11202), .O(n11205));
  LUT5 #(.INIT(32'hFF969600)) lut_n11206 (.I0(x2433), .I1(x2434), .I2(x2435), .I3(n11204), .I4(n11205), .O(n11206));
  LUT3 #(.INIT(8'h96)) lut_n11207 (.I0(n11187), .I1(n11190), .I2(n11191), .O(n11207));
  LUT3 #(.INIT(8'hE8)) lut_n11208 (.I0(n11203), .I1(n11206), .I2(n11207), .O(n11208));
  LUT3 #(.INIT(8'h96)) lut_n11209 (.I0(x2442), .I1(x2443), .I2(x2444), .O(n11209));
  LUT5 #(.INIT(32'h96696996)) lut_n11210 (.I0(x2433), .I1(x2434), .I2(x2435), .I3(n11204), .I4(n11205), .O(n11210));
  LUT5 #(.INIT(32'hFF969600)) lut_n11211 (.I0(x2439), .I1(x2440), .I2(x2441), .I3(n11209), .I4(n11210), .O(n11211));
  LUT3 #(.INIT(8'h96)) lut_n11212 (.I0(x2448), .I1(x2449), .I2(x2450), .O(n11212));
  LUT5 #(.INIT(32'h96696996)) lut_n11213 (.I0(x2439), .I1(x2440), .I2(x2441), .I3(n11209), .I4(n11210), .O(n11213));
  LUT5 #(.INIT(32'hFF969600)) lut_n11214 (.I0(x2445), .I1(x2446), .I2(x2447), .I3(n11212), .I4(n11213), .O(n11214));
  LUT3 #(.INIT(8'h96)) lut_n11215 (.I0(n11203), .I1(n11206), .I2(n11207), .O(n11215));
  LUT3 #(.INIT(8'hE8)) lut_n11216 (.I0(n11211), .I1(n11214), .I2(n11215), .O(n11216));
  LUT3 #(.INIT(8'h96)) lut_n11217 (.I0(n11184), .I1(n11192), .I2(n11193), .O(n11217));
  LUT3 #(.INIT(8'hE8)) lut_n11218 (.I0(n11208), .I1(n11216), .I2(n11217), .O(n11218));
  LUT3 #(.INIT(8'h96)) lut_n11219 (.I0(x2454), .I1(x2455), .I2(x2456), .O(n11219));
  LUT5 #(.INIT(32'h96696996)) lut_n11220 (.I0(x2445), .I1(x2446), .I2(x2447), .I3(n11212), .I4(n11213), .O(n11220));
  LUT5 #(.INIT(32'hFF969600)) lut_n11221 (.I0(x2451), .I1(x2452), .I2(x2453), .I3(n11219), .I4(n11220), .O(n11221));
  LUT3 #(.INIT(8'h96)) lut_n11222 (.I0(x2460), .I1(x2461), .I2(x2462), .O(n11222));
  LUT5 #(.INIT(32'h96696996)) lut_n11223 (.I0(x2451), .I1(x2452), .I2(x2453), .I3(n11219), .I4(n11220), .O(n11223));
  LUT5 #(.INIT(32'hFF969600)) lut_n11224 (.I0(x2457), .I1(x2458), .I2(x2459), .I3(n11222), .I4(n11223), .O(n11224));
  LUT3 #(.INIT(8'h96)) lut_n11225 (.I0(n11211), .I1(n11214), .I2(n11215), .O(n11225));
  LUT3 #(.INIT(8'hE8)) lut_n11226 (.I0(n11221), .I1(n11224), .I2(n11225), .O(n11226));
  LUT3 #(.INIT(8'h96)) lut_n11227 (.I0(x2466), .I1(x2467), .I2(x2468), .O(n11227));
  LUT5 #(.INIT(32'h96696996)) lut_n11228 (.I0(x2457), .I1(x2458), .I2(x2459), .I3(n11222), .I4(n11223), .O(n11228));
  LUT5 #(.INIT(32'hFF969600)) lut_n11229 (.I0(x2463), .I1(x2464), .I2(x2465), .I3(n11227), .I4(n11228), .O(n11229));
  LUT3 #(.INIT(8'h96)) lut_n11230 (.I0(x2472), .I1(x2473), .I2(x2474), .O(n11230));
  LUT5 #(.INIT(32'h96696996)) lut_n11231 (.I0(x2463), .I1(x2464), .I2(x2465), .I3(n11227), .I4(n11228), .O(n11231));
  LUT5 #(.INIT(32'hFF969600)) lut_n11232 (.I0(x2469), .I1(x2470), .I2(x2471), .I3(n11230), .I4(n11231), .O(n11232));
  LUT3 #(.INIT(8'h96)) lut_n11233 (.I0(n11221), .I1(n11224), .I2(n11225), .O(n11233));
  LUT3 #(.INIT(8'hE8)) lut_n11234 (.I0(n11229), .I1(n11232), .I2(n11233), .O(n11234));
  LUT3 #(.INIT(8'h96)) lut_n11235 (.I0(n11208), .I1(n11216), .I2(n11217), .O(n11235));
  LUT3 #(.INIT(8'hE8)) lut_n11236 (.I0(n11226), .I1(n11234), .I2(n11235), .O(n11236));
  LUT3 #(.INIT(8'h96)) lut_n11237 (.I0(n11176), .I1(n11194), .I2(n11195), .O(n11237));
  LUT3 #(.INIT(8'hE8)) lut_n11238 (.I0(n11218), .I1(n11236), .I2(n11237), .O(n11238));
  LUT3 #(.INIT(8'h96)) lut_n11239 (.I0(x2478), .I1(x2479), .I2(x2480), .O(n11239));
  LUT5 #(.INIT(32'h96696996)) lut_n11240 (.I0(x2469), .I1(x2470), .I2(x2471), .I3(n11230), .I4(n11231), .O(n11240));
  LUT5 #(.INIT(32'hFF969600)) lut_n11241 (.I0(x2475), .I1(x2476), .I2(x2477), .I3(n11239), .I4(n11240), .O(n11241));
  LUT3 #(.INIT(8'h96)) lut_n11242 (.I0(x2484), .I1(x2485), .I2(x2486), .O(n11242));
  LUT5 #(.INIT(32'h96696996)) lut_n11243 (.I0(x2475), .I1(x2476), .I2(x2477), .I3(n11239), .I4(n11240), .O(n11243));
  LUT5 #(.INIT(32'hFF969600)) lut_n11244 (.I0(x2481), .I1(x2482), .I2(x2483), .I3(n11242), .I4(n11243), .O(n11244));
  LUT3 #(.INIT(8'h96)) lut_n11245 (.I0(n11229), .I1(n11232), .I2(n11233), .O(n11245));
  LUT3 #(.INIT(8'hE8)) lut_n11246 (.I0(n11241), .I1(n11244), .I2(n11245), .O(n11246));
  LUT3 #(.INIT(8'h96)) lut_n11247 (.I0(x2490), .I1(x2491), .I2(x2492), .O(n11247));
  LUT5 #(.INIT(32'h96696996)) lut_n11248 (.I0(x2481), .I1(x2482), .I2(x2483), .I3(n11242), .I4(n11243), .O(n11248));
  LUT5 #(.INIT(32'hFF969600)) lut_n11249 (.I0(x2487), .I1(x2488), .I2(x2489), .I3(n11247), .I4(n11248), .O(n11249));
  LUT3 #(.INIT(8'h96)) lut_n11250 (.I0(x2496), .I1(x2497), .I2(x2498), .O(n11250));
  LUT5 #(.INIT(32'h96696996)) lut_n11251 (.I0(x2487), .I1(x2488), .I2(x2489), .I3(n11247), .I4(n11248), .O(n11251));
  LUT5 #(.INIT(32'hFF969600)) lut_n11252 (.I0(x2493), .I1(x2494), .I2(x2495), .I3(n11250), .I4(n11251), .O(n11252));
  LUT3 #(.INIT(8'h96)) lut_n11253 (.I0(n11241), .I1(n11244), .I2(n11245), .O(n11253));
  LUT3 #(.INIT(8'hE8)) lut_n11254 (.I0(n11249), .I1(n11252), .I2(n11253), .O(n11254));
  LUT3 #(.INIT(8'h96)) lut_n11255 (.I0(n11226), .I1(n11234), .I2(n11235), .O(n11255));
  LUT3 #(.INIT(8'hE8)) lut_n11256 (.I0(n11246), .I1(n11254), .I2(n11255), .O(n11256));
  LUT3 #(.INIT(8'h96)) lut_n11257 (.I0(x2502), .I1(x2503), .I2(x2504), .O(n11257));
  LUT5 #(.INIT(32'h96696996)) lut_n11258 (.I0(x2493), .I1(x2494), .I2(x2495), .I3(n11250), .I4(n11251), .O(n11258));
  LUT5 #(.INIT(32'hFF969600)) lut_n11259 (.I0(x2499), .I1(x2500), .I2(x2501), .I3(n11257), .I4(n11258), .O(n11259));
  LUT3 #(.INIT(8'h96)) lut_n11260 (.I0(x2508), .I1(x2509), .I2(x2510), .O(n11260));
  LUT5 #(.INIT(32'h96696996)) lut_n11261 (.I0(x2499), .I1(x2500), .I2(x2501), .I3(n11257), .I4(n11258), .O(n11261));
  LUT5 #(.INIT(32'hFF969600)) lut_n11262 (.I0(x2505), .I1(x2506), .I2(x2507), .I3(n11260), .I4(n11261), .O(n11262));
  LUT3 #(.INIT(8'h96)) lut_n11263 (.I0(n11249), .I1(n11252), .I2(n11253), .O(n11263));
  LUT3 #(.INIT(8'hE8)) lut_n11264 (.I0(n11259), .I1(n11262), .I2(n11263), .O(n11264));
  LUT3 #(.INIT(8'h96)) lut_n11265 (.I0(x2514), .I1(x2515), .I2(x2516), .O(n11265));
  LUT5 #(.INIT(32'h96696996)) lut_n11266 (.I0(x2505), .I1(x2506), .I2(x2507), .I3(n11260), .I4(n11261), .O(n11266));
  LUT5 #(.INIT(32'hFF969600)) lut_n11267 (.I0(x2511), .I1(x2512), .I2(x2513), .I3(n11265), .I4(n11266), .O(n11267));
  LUT3 #(.INIT(8'h96)) lut_n11268 (.I0(x2520), .I1(x2521), .I2(x2522), .O(n11268));
  LUT5 #(.INIT(32'h96696996)) lut_n11269 (.I0(x2511), .I1(x2512), .I2(x2513), .I3(n11265), .I4(n11266), .O(n11269));
  LUT5 #(.INIT(32'hFF969600)) lut_n11270 (.I0(x2517), .I1(x2518), .I2(x2519), .I3(n11268), .I4(n11269), .O(n11270));
  LUT3 #(.INIT(8'h96)) lut_n11271 (.I0(n11259), .I1(n11262), .I2(n11263), .O(n11271));
  LUT3 #(.INIT(8'hE8)) lut_n11272 (.I0(n11267), .I1(n11270), .I2(n11271), .O(n11272));
  LUT3 #(.INIT(8'h96)) lut_n11273 (.I0(n11246), .I1(n11254), .I2(n11255), .O(n11273));
  LUT3 #(.INIT(8'hE8)) lut_n11274 (.I0(n11264), .I1(n11272), .I2(n11273), .O(n11274));
  LUT3 #(.INIT(8'h96)) lut_n11275 (.I0(n11218), .I1(n11236), .I2(n11237), .O(n11275));
  LUT3 #(.INIT(8'hE8)) lut_n11276 (.I0(n11256), .I1(n11274), .I2(n11275), .O(n11276));
  LUT3 #(.INIT(8'h96)) lut_n11277 (.I0(n11158), .I1(n11196), .I2(n11197), .O(n11277));
  LUT3 #(.INIT(8'hE8)) lut_n11278 (.I0(n11238), .I1(n11276), .I2(n11277), .O(n11278));
  LUT3 #(.INIT(8'h96)) lut_n11279 (.I0(x2526), .I1(x2527), .I2(x2528), .O(n11279));
  LUT5 #(.INIT(32'h96696996)) lut_n11280 (.I0(x2517), .I1(x2518), .I2(x2519), .I3(n11268), .I4(n11269), .O(n11280));
  LUT5 #(.INIT(32'hFF969600)) lut_n11281 (.I0(x2523), .I1(x2524), .I2(x2525), .I3(n11279), .I4(n11280), .O(n11281));
  LUT3 #(.INIT(8'h96)) lut_n11282 (.I0(x2532), .I1(x2533), .I2(x2534), .O(n11282));
  LUT5 #(.INIT(32'h96696996)) lut_n11283 (.I0(x2523), .I1(x2524), .I2(x2525), .I3(n11279), .I4(n11280), .O(n11283));
  LUT5 #(.INIT(32'hFF969600)) lut_n11284 (.I0(x2529), .I1(x2530), .I2(x2531), .I3(n11282), .I4(n11283), .O(n11284));
  LUT3 #(.INIT(8'h96)) lut_n11285 (.I0(n11267), .I1(n11270), .I2(n11271), .O(n11285));
  LUT3 #(.INIT(8'hE8)) lut_n11286 (.I0(n11281), .I1(n11284), .I2(n11285), .O(n11286));
  LUT3 #(.INIT(8'h96)) lut_n11287 (.I0(x2538), .I1(x2539), .I2(x2540), .O(n11287));
  LUT5 #(.INIT(32'h96696996)) lut_n11288 (.I0(x2529), .I1(x2530), .I2(x2531), .I3(n11282), .I4(n11283), .O(n11288));
  LUT5 #(.INIT(32'hFF969600)) lut_n11289 (.I0(x2535), .I1(x2536), .I2(x2537), .I3(n11287), .I4(n11288), .O(n11289));
  LUT3 #(.INIT(8'h96)) lut_n11290 (.I0(x2544), .I1(x2545), .I2(x2546), .O(n11290));
  LUT5 #(.INIT(32'h96696996)) lut_n11291 (.I0(x2535), .I1(x2536), .I2(x2537), .I3(n11287), .I4(n11288), .O(n11291));
  LUT5 #(.INIT(32'hFF969600)) lut_n11292 (.I0(x2541), .I1(x2542), .I2(x2543), .I3(n11290), .I4(n11291), .O(n11292));
  LUT3 #(.INIT(8'h96)) lut_n11293 (.I0(n11281), .I1(n11284), .I2(n11285), .O(n11293));
  LUT3 #(.INIT(8'hE8)) lut_n11294 (.I0(n11289), .I1(n11292), .I2(n11293), .O(n11294));
  LUT3 #(.INIT(8'h96)) lut_n11295 (.I0(n11264), .I1(n11272), .I2(n11273), .O(n11295));
  LUT3 #(.INIT(8'hE8)) lut_n11296 (.I0(n11286), .I1(n11294), .I2(n11295), .O(n11296));
  LUT3 #(.INIT(8'h96)) lut_n11297 (.I0(x2550), .I1(x2551), .I2(x2552), .O(n11297));
  LUT5 #(.INIT(32'h96696996)) lut_n11298 (.I0(x2541), .I1(x2542), .I2(x2543), .I3(n11290), .I4(n11291), .O(n11298));
  LUT5 #(.INIT(32'hFF969600)) lut_n11299 (.I0(x2547), .I1(x2548), .I2(x2549), .I3(n11297), .I4(n11298), .O(n11299));
  LUT3 #(.INIT(8'h96)) lut_n11300 (.I0(x2556), .I1(x2557), .I2(x2558), .O(n11300));
  LUT5 #(.INIT(32'h96696996)) lut_n11301 (.I0(x2547), .I1(x2548), .I2(x2549), .I3(n11297), .I4(n11298), .O(n11301));
  LUT5 #(.INIT(32'hFF969600)) lut_n11302 (.I0(x2553), .I1(x2554), .I2(x2555), .I3(n11300), .I4(n11301), .O(n11302));
  LUT3 #(.INIT(8'h96)) lut_n11303 (.I0(n11289), .I1(n11292), .I2(n11293), .O(n11303));
  LUT3 #(.INIT(8'hE8)) lut_n11304 (.I0(n11299), .I1(n11302), .I2(n11303), .O(n11304));
  LUT3 #(.INIT(8'h96)) lut_n11305 (.I0(x2562), .I1(x2563), .I2(x2564), .O(n11305));
  LUT5 #(.INIT(32'h96696996)) lut_n11306 (.I0(x2553), .I1(x2554), .I2(x2555), .I3(n11300), .I4(n11301), .O(n11306));
  LUT5 #(.INIT(32'hFF969600)) lut_n11307 (.I0(x2559), .I1(x2560), .I2(x2561), .I3(n11305), .I4(n11306), .O(n11307));
  LUT3 #(.INIT(8'h96)) lut_n11308 (.I0(x2568), .I1(x2569), .I2(x2570), .O(n11308));
  LUT5 #(.INIT(32'h96696996)) lut_n11309 (.I0(x2559), .I1(x2560), .I2(x2561), .I3(n11305), .I4(n11306), .O(n11309));
  LUT5 #(.INIT(32'hFF969600)) lut_n11310 (.I0(x2565), .I1(x2566), .I2(x2567), .I3(n11308), .I4(n11309), .O(n11310));
  LUT3 #(.INIT(8'h96)) lut_n11311 (.I0(n11299), .I1(n11302), .I2(n11303), .O(n11311));
  LUT3 #(.INIT(8'hE8)) lut_n11312 (.I0(n11307), .I1(n11310), .I2(n11311), .O(n11312));
  LUT3 #(.INIT(8'h96)) lut_n11313 (.I0(n11286), .I1(n11294), .I2(n11295), .O(n11313));
  LUT3 #(.INIT(8'hE8)) lut_n11314 (.I0(n11304), .I1(n11312), .I2(n11313), .O(n11314));
  LUT3 #(.INIT(8'h96)) lut_n11315 (.I0(n11256), .I1(n11274), .I2(n11275), .O(n11315));
  LUT3 #(.INIT(8'hE8)) lut_n11316 (.I0(n11296), .I1(n11314), .I2(n11315), .O(n11316));
  LUT3 #(.INIT(8'h96)) lut_n11317 (.I0(x2574), .I1(x2575), .I2(x2576), .O(n11317));
  LUT5 #(.INIT(32'h96696996)) lut_n11318 (.I0(x2565), .I1(x2566), .I2(x2567), .I3(n11308), .I4(n11309), .O(n11318));
  LUT5 #(.INIT(32'hFF969600)) lut_n11319 (.I0(x2571), .I1(x2572), .I2(x2573), .I3(n11317), .I4(n11318), .O(n11319));
  LUT3 #(.INIT(8'h96)) lut_n11320 (.I0(x2580), .I1(x2581), .I2(x2582), .O(n11320));
  LUT5 #(.INIT(32'h96696996)) lut_n11321 (.I0(x2571), .I1(x2572), .I2(x2573), .I3(n11317), .I4(n11318), .O(n11321));
  LUT5 #(.INIT(32'hFF969600)) lut_n11322 (.I0(x2577), .I1(x2578), .I2(x2579), .I3(n11320), .I4(n11321), .O(n11322));
  LUT3 #(.INIT(8'h96)) lut_n11323 (.I0(n11307), .I1(n11310), .I2(n11311), .O(n11323));
  LUT3 #(.INIT(8'hE8)) lut_n11324 (.I0(n11319), .I1(n11322), .I2(n11323), .O(n11324));
  LUT3 #(.INIT(8'h96)) lut_n11325 (.I0(x2586), .I1(x2587), .I2(x2588), .O(n11325));
  LUT5 #(.INIT(32'h96696996)) lut_n11326 (.I0(x2577), .I1(x2578), .I2(x2579), .I3(n11320), .I4(n11321), .O(n11326));
  LUT5 #(.INIT(32'hFF969600)) lut_n11327 (.I0(x2583), .I1(x2584), .I2(x2585), .I3(n11325), .I4(n11326), .O(n11327));
  LUT3 #(.INIT(8'h96)) lut_n11328 (.I0(x2592), .I1(x2593), .I2(x2594), .O(n11328));
  LUT5 #(.INIT(32'h96696996)) lut_n11329 (.I0(x2583), .I1(x2584), .I2(x2585), .I3(n11325), .I4(n11326), .O(n11329));
  LUT5 #(.INIT(32'hFF969600)) lut_n11330 (.I0(x2589), .I1(x2590), .I2(x2591), .I3(n11328), .I4(n11329), .O(n11330));
  LUT3 #(.INIT(8'h96)) lut_n11331 (.I0(n11319), .I1(n11322), .I2(n11323), .O(n11331));
  LUT3 #(.INIT(8'hE8)) lut_n11332 (.I0(n11327), .I1(n11330), .I2(n11331), .O(n11332));
  LUT3 #(.INIT(8'h96)) lut_n11333 (.I0(n11304), .I1(n11312), .I2(n11313), .O(n11333));
  LUT3 #(.INIT(8'hE8)) lut_n11334 (.I0(n11324), .I1(n11332), .I2(n11333), .O(n11334));
  LUT3 #(.INIT(8'h96)) lut_n11335 (.I0(x2598), .I1(x2599), .I2(x2600), .O(n11335));
  LUT5 #(.INIT(32'h96696996)) lut_n11336 (.I0(x2589), .I1(x2590), .I2(x2591), .I3(n11328), .I4(n11329), .O(n11336));
  LUT5 #(.INIT(32'hFF969600)) lut_n11337 (.I0(x2595), .I1(x2596), .I2(x2597), .I3(n11335), .I4(n11336), .O(n11337));
  LUT3 #(.INIT(8'h96)) lut_n11338 (.I0(x2604), .I1(x2605), .I2(x2606), .O(n11338));
  LUT5 #(.INIT(32'h96696996)) lut_n11339 (.I0(x2595), .I1(x2596), .I2(x2597), .I3(n11335), .I4(n11336), .O(n11339));
  LUT5 #(.INIT(32'hFF969600)) lut_n11340 (.I0(x2601), .I1(x2602), .I2(x2603), .I3(n11338), .I4(n11339), .O(n11340));
  LUT3 #(.INIT(8'h96)) lut_n11341 (.I0(n11327), .I1(n11330), .I2(n11331), .O(n11341));
  LUT3 #(.INIT(8'hE8)) lut_n11342 (.I0(n11337), .I1(n11340), .I2(n11341), .O(n11342));
  LUT3 #(.INIT(8'h96)) lut_n11343 (.I0(x2610), .I1(x2611), .I2(x2612), .O(n11343));
  LUT5 #(.INIT(32'h96696996)) lut_n11344 (.I0(x2601), .I1(x2602), .I2(x2603), .I3(n11338), .I4(n11339), .O(n11344));
  LUT5 #(.INIT(32'hFF969600)) lut_n11345 (.I0(x2607), .I1(x2608), .I2(x2609), .I3(n11343), .I4(n11344), .O(n11345));
  LUT3 #(.INIT(8'h96)) lut_n11346 (.I0(x2616), .I1(x2617), .I2(x2618), .O(n11346));
  LUT5 #(.INIT(32'h96696996)) lut_n11347 (.I0(x2607), .I1(x2608), .I2(x2609), .I3(n11343), .I4(n11344), .O(n11347));
  LUT5 #(.INIT(32'hFF969600)) lut_n11348 (.I0(x2613), .I1(x2614), .I2(x2615), .I3(n11346), .I4(n11347), .O(n11348));
  LUT3 #(.INIT(8'h96)) lut_n11349 (.I0(n11337), .I1(n11340), .I2(n11341), .O(n11349));
  LUT3 #(.INIT(8'hE8)) lut_n11350 (.I0(n11345), .I1(n11348), .I2(n11349), .O(n11350));
  LUT3 #(.INIT(8'h96)) lut_n11351 (.I0(n11324), .I1(n11332), .I2(n11333), .O(n11351));
  LUT3 #(.INIT(8'hE8)) lut_n11352 (.I0(n11342), .I1(n11350), .I2(n11351), .O(n11352));
  LUT3 #(.INIT(8'h96)) lut_n11353 (.I0(n11296), .I1(n11314), .I2(n11315), .O(n11353));
  LUT3 #(.INIT(8'hE8)) lut_n11354 (.I0(n11334), .I1(n11352), .I2(n11353), .O(n11354));
  LUT3 #(.INIT(8'h96)) lut_n11355 (.I0(n11238), .I1(n11276), .I2(n11277), .O(n11355));
  LUT3 #(.INIT(8'hE8)) lut_n11356 (.I0(n11316), .I1(n11354), .I2(n11355), .O(n11356));
  LUT3 #(.INIT(8'h96)) lut_n11357 (.I0(n11120), .I1(n11198), .I2(n11199), .O(n11357));
  LUT3 #(.INIT(8'hE8)) lut_n11358 (.I0(n11278), .I1(n11356), .I2(n11357), .O(n11358));
  LUT3 #(.INIT(8'h96)) lut_n11359 (.I0(n10875), .I1(n11033), .I2(n11034), .O(n11359));
  LUT3 #(.INIT(8'hE8)) lut_n11360 (.I0(n11200), .I1(n11358), .I2(n11359), .O(n11360));
  LUT3 #(.INIT(8'h96)) lut_n11361 (.I0(x2622), .I1(x2623), .I2(x2624), .O(n11361));
  LUT5 #(.INIT(32'h96696996)) lut_n11362 (.I0(x2613), .I1(x2614), .I2(x2615), .I3(n11346), .I4(n11347), .O(n11362));
  LUT5 #(.INIT(32'hFF969600)) lut_n11363 (.I0(x2619), .I1(x2620), .I2(x2621), .I3(n11361), .I4(n11362), .O(n11363));
  LUT3 #(.INIT(8'h96)) lut_n11364 (.I0(x2628), .I1(x2629), .I2(x2630), .O(n11364));
  LUT5 #(.INIT(32'h96696996)) lut_n11365 (.I0(x2619), .I1(x2620), .I2(x2621), .I3(n11361), .I4(n11362), .O(n11365));
  LUT5 #(.INIT(32'hFF969600)) lut_n11366 (.I0(x2625), .I1(x2626), .I2(x2627), .I3(n11364), .I4(n11365), .O(n11366));
  LUT3 #(.INIT(8'h96)) lut_n11367 (.I0(n11345), .I1(n11348), .I2(n11349), .O(n11367));
  LUT3 #(.INIT(8'hE8)) lut_n11368 (.I0(n11363), .I1(n11366), .I2(n11367), .O(n11368));
  LUT3 #(.INIT(8'h96)) lut_n11369 (.I0(x2634), .I1(x2635), .I2(x2636), .O(n11369));
  LUT5 #(.INIT(32'h96696996)) lut_n11370 (.I0(x2625), .I1(x2626), .I2(x2627), .I3(n11364), .I4(n11365), .O(n11370));
  LUT5 #(.INIT(32'hFF969600)) lut_n11371 (.I0(x2631), .I1(x2632), .I2(x2633), .I3(n11369), .I4(n11370), .O(n11371));
  LUT3 #(.INIT(8'h96)) lut_n11372 (.I0(x2640), .I1(x2641), .I2(x2642), .O(n11372));
  LUT5 #(.INIT(32'h96696996)) lut_n11373 (.I0(x2631), .I1(x2632), .I2(x2633), .I3(n11369), .I4(n11370), .O(n11373));
  LUT5 #(.INIT(32'hFF969600)) lut_n11374 (.I0(x2637), .I1(x2638), .I2(x2639), .I3(n11372), .I4(n11373), .O(n11374));
  LUT3 #(.INIT(8'h96)) lut_n11375 (.I0(n11363), .I1(n11366), .I2(n11367), .O(n11375));
  LUT3 #(.INIT(8'hE8)) lut_n11376 (.I0(n11371), .I1(n11374), .I2(n11375), .O(n11376));
  LUT3 #(.INIT(8'h96)) lut_n11377 (.I0(n11342), .I1(n11350), .I2(n11351), .O(n11377));
  LUT3 #(.INIT(8'hE8)) lut_n11378 (.I0(n11368), .I1(n11376), .I2(n11377), .O(n11378));
  LUT3 #(.INIT(8'h96)) lut_n11379 (.I0(x2646), .I1(x2647), .I2(x2648), .O(n11379));
  LUT5 #(.INIT(32'h96696996)) lut_n11380 (.I0(x2637), .I1(x2638), .I2(x2639), .I3(n11372), .I4(n11373), .O(n11380));
  LUT5 #(.INIT(32'hFF969600)) lut_n11381 (.I0(x2643), .I1(x2644), .I2(x2645), .I3(n11379), .I4(n11380), .O(n11381));
  LUT3 #(.INIT(8'h96)) lut_n11382 (.I0(x2652), .I1(x2653), .I2(x2654), .O(n11382));
  LUT5 #(.INIT(32'h96696996)) lut_n11383 (.I0(x2643), .I1(x2644), .I2(x2645), .I3(n11379), .I4(n11380), .O(n11383));
  LUT5 #(.INIT(32'hFF969600)) lut_n11384 (.I0(x2649), .I1(x2650), .I2(x2651), .I3(n11382), .I4(n11383), .O(n11384));
  LUT3 #(.INIT(8'h96)) lut_n11385 (.I0(n11371), .I1(n11374), .I2(n11375), .O(n11385));
  LUT3 #(.INIT(8'hE8)) lut_n11386 (.I0(n11381), .I1(n11384), .I2(n11385), .O(n11386));
  LUT3 #(.INIT(8'h96)) lut_n11387 (.I0(x2658), .I1(x2659), .I2(x2660), .O(n11387));
  LUT5 #(.INIT(32'h96696996)) lut_n11388 (.I0(x2649), .I1(x2650), .I2(x2651), .I3(n11382), .I4(n11383), .O(n11388));
  LUT5 #(.INIT(32'hFF969600)) lut_n11389 (.I0(x2655), .I1(x2656), .I2(x2657), .I3(n11387), .I4(n11388), .O(n11389));
  LUT3 #(.INIT(8'h96)) lut_n11390 (.I0(x2664), .I1(x2665), .I2(x2666), .O(n11390));
  LUT5 #(.INIT(32'h96696996)) lut_n11391 (.I0(x2655), .I1(x2656), .I2(x2657), .I3(n11387), .I4(n11388), .O(n11391));
  LUT5 #(.INIT(32'hFF969600)) lut_n11392 (.I0(x2661), .I1(x2662), .I2(x2663), .I3(n11390), .I4(n11391), .O(n11392));
  LUT3 #(.INIT(8'h96)) lut_n11393 (.I0(n11381), .I1(n11384), .I2(n11385), .O(n11393));
  LUT3 #(.INIT(8'hE8)) lut_n11394 (.I0(n11389), .I1(n11392), .I2(n11393), .O(n11394));
  LUT3 #(.INIT(8'h96)) lut_n11395 (.I0(n11368), .I1(n11376), .I2(n11377), .O(n11395));
  LUT3 #(.INIT(8'hE8)) lut_n11396 (.I0(n11386), .I1(n11394), .I2(n11395), .O(n11396));
  LUT3 #(.INIT(8'h96)) lut_n11397 (.I0(n11334), .I1(n11352), .I2(n11353), .O(n11397));
  LUT3 #(.INIT(8'hE8)) lut_n11398 (.I0(n11378), .I1(n11396), .I2(n11397), .O(n11398));
  LUT3 #(.INIT(8'h96)) lut_n11399 (.I0(x2670), .I1(x2671), .I2(x2672), .O(n11399));
  LUT5 #(.INIT(32'h96696996)) lut_n11400 (.I0(x2661), .I1(x2662), .I2(x2663), .I3(n11390), .I4(n11391), .O(n11400));
  LUT5 #(.INIT(32'hFF969600)) lut_n11401 (.I0(x2667), .I1(x2668), .I2(x2669), .I3(n11399), .I4(n11400), .O(n11401));
  LUT3 #(.INIT(8'h96)) lut_n11402 (.I0(x2676), .I1(x2677), .I2(x2678), .O(n11402));
  LUT5 #(.INIT(32'h96696996)) lut_n11403 (.I0(x2667), .I1(x2668), .I2(x2669), .I3(n11399), .I4(n11400), .O(n11403));
  LUT5 #(.INIT(32'hFF969600)) lut_n11404 (.I0(x2673), .I1(x2674), .I2(x2675), .I3(n11402), .I4(n11403), .O(n11404));
  LUT3 #(.INIT(8'h96)) lut_n11405 (.I0(n11389), .I1(n11392), .I2(n11393), .O(n11405));
  LUT3 #(.INIT(8'hE8)) lut_n11406 (.I0(n11401), .I1(n11404), .I2(n11405), .O(n11406));
  LUT3 #(.INIT(8'h96)) lut_n11407 (.I0(x2682), .I1(x2683), .I2(x2684), .O(n11407));
  LUT5 #(.INIT(32'h96696996)) lut_n11408 (.I0(x2673), .I1(x2674), .I2(x2675), .I3(n11402), .I4(n11403), .O(n11408));
  LUT5 #(.INIT(32'hFF969600)) lut_n11409 (.I0(x2679), .I1(x2680), .I2(x2681), .I3(n11407), .I4(n11408), .O(n11409));
  LUT3 #(.INIT(8'h96)) lut_n11410 (.I0(x2688), .I1(x2689), .I2(x2690), .O(n11410));
  LUT5 #(.INIT(32'h96696996)) lut_n11411 (.I0(x2679), .I1(x2680), .I2(x2681), .I3(n11407), .I4(n11408), .O(n11411));
  LUT5 #(.INIT(32'hFF969600)) lut_n11412 (.I0(x2685), .I1(x2686), .I2(x2687), .I3(n11410), .I4(n11411), .O(n11412));
  LUT3 #(.INIT(8'h96)) lut_n11413 (.I0(n11401), .I1(n11404), .I2(n11405), .O(n11413));
  LUT3 #(.INIT(8'hE8)) lut_n11414 (.I0(n11409), .I1(n11412), .I2(n11413), .O(n11414));
  LUT3 #(.INIT(8'h96)) lut_n11415 (.I0(n11386), .I1(n11394), .I2(n11395), .O(n11415));
  LUT3 #(.INIT(8'hE8)) lut_n11416 (.I0(n11406), .I1(n11414), .I2(n11415), .O(n11416));
  LUT3 #(.INIT(8'h96)) lut_n11417 (.I0(x2694), .I1(x2695), .I2(x2696), .O(n11417));
  LUT5 #(.INIT(32'h96696996)) lut_n11418 (.I0(x2685), .I1(x2686), .I2(x2687), .I3(n11410), .I4(n11411), .O(n11418));
  LUT5 #(.INIT(32'hFF969600)) lut_n11419 (.I0(x2691), .I1(x2692), .I2(x2693), .I3(n11417), .I4(n11418), .O(n11419));
  LUT3 #(.INIT(8'h96)) lut_n11420 (.I0(x2700), .I1(x2701), .I2(x2702), .O(n11420));
  LUT5 #(.INIT(32'h96696996)) lut_n11421 (.I0(x2691), .I1(x2692), .I2(x2693), .I3(n11417), .I4(n11418), .O(n11421));
  LUT5 #(.INIT(32'hFF969600)) lut_n11422 (.I0(x2697), .I1(x2698), .I2(x2699), .I3(n11420), .I4(n11421), .O(n11422));
  LUT3 #(.INIT(8'h96)) lut_n11423 (.I0(n11409), .I1(n11412), .I2(n11413), .O(n11423));
  LUT3 #(.INIT(8'hE8)) lut_n11424 (.I0(n11419), .I1(n11422), .I2(n11423), .O(n11424));
  LUT3 #(.INIT(8'h96)) lut_n11425 (.I0(x2706), .I1(x2707), .I2(x2708), .O(n11425));
  LUT5 #(.INIT(32'h96696996)) lut_n11426 (.I0(x2697), .I1(x2698), .I2(x2699), .I3(n11420), .I4(n11421), .O(n11426));
  LUT5 #(.INIT(32'hFF969600)) lut_n11427 (.I0(x2703), .I1(x2704), .I2(x2705), .I3(n11425), .I4(n11426), .O(n11427));
  LUT3 #(.INIT(8'h96)) lut_n11428 (.I0(x2712), .I1(x2713), .I2(x2714), .O(n11428));
  LUT5 #(.INIT(32'h96696996)) lut_n11429 (.I0(x2703), .I1(x2704), .I2(x2705), .I3(n11425), .I4(n11426), .O(n11429));
  LUT5 #(.INIT(32'hFF969600)) lut_n11430 (.I0(x2709), .I1(x2710), .I2(x2711), .I3(n11428), .I4(n11429), .O(n11430));
  LUT3 #(.INIT(8'h96)) lut_n11431 (.I0(n11419), .I1(n11422), .I2(n11423), .O(n11431));
  LUT3 #(.INIT(8'hE8)) lut_n11432 (.I0(n11427), .I1(n11430), .I2(n11431), .O(n11432));
  LUT3 #(.INIT(8'h96)) lut_n11433 (.I0(n11406), .I1(n11414), .I2(n11415), .O(n11433));
  LUT3 #(.INIT(8'hE8)) lut_n11434 (.I0(n11424), .I1(n11432), .I2(n11433), .O(n11434));
  LUT3 #(.INIT(8'h96)) lut_n11435 (.I0(n11378), .I1(n11396), .I2(n11397), .O(n11435));
  LUT3 #(.INIT(8'hE8)) lut_n11436 (.I0(n11416), .I1(n11434), .I2(n11435), .O(n11436));
  LUT3 #(.INIT(8'h96)) lut_n11437 (.I0(n11316), .I1(n11354), .I2(n11355), .O(n11437));
  LUT3 #(.INIT(8'hE8)) lut_n11438 (.I0(n11398), .I1(n11436), .I2(n11437), .O(n11438));
  LUT3 #(.INIT(8'h96)) lut_n11439 (.I0(x2718), .I1(x2719), .I2(x2720), .O(n11439));
  LUT5 #(.INIT(32'h96696996)) lut_n11440 (.I0(x2709), .I1(x2710), .I2(x2711), .I3(n11428), .I4(n11429), .O(n11440));
  LUT5 #(.INIT(32'hFF969600)) lut_n11441 (.I0(x2715), .I1(x2716), .I2(x2717), .I3(n11439), .I4(n11440), .O(n11441));
  LUT3 #(.INIT(8'h96)) lut_n11442 (.I0(x2724), .I1(x2725), .I2(x2726), .O(n11442));
  LUT5 #(.INIT(32'h96696996)) lut_n11443 (.I0(x2715), .I1(x2716), .I2(x2717), .I3(n11439), .I4(n11440), .O(n11443));
  LUT5 #(.INIT(32'hFF969600)) lut_n11444 (.I0(x2721), .I1(x2722), .I2(x2723), .I3(n11442), .I4(n11443), .O(n11444));
  LUT3 #(.INIT(8'h96)) lut_n11445 (.I0(n11427), .I1(n11430), .I2(n11431), .O(n11445));
  LUT3 #(.INIT(8'hE8)) lut_n11446 (.I0(n11441), .I1(n11444), .I2(n11445), .O(n11446));
  LUT3 #(.INIT(8'h96)) lut_n11447 (.I0(x2730), .I1(x2731), .I2(x2732), .O(n11447));
  LUT5 #(.INIT(32'h96696996)) lut_n11448 (.I0(x2721), .I1(x2722), .I2(x2723), .I3(n11442), .I4(n11443), .O(n11448));
  LUT5 #(.INIT(32'hFF969600)) lut_n11449 (.I0(x2727), .I1(x2728), .I2(x2729), .I3(n11447), .I4(n11448), .O(n11449));
  LUT3 #(.INIT(8'h96)) lut_n11450 (.I0(x2736), .I1(x2737), .I2(x2738), .O(n11450));
  LUT5 #(.INIT(32'h96696996)) lut_n11451 (.I0(x2727), .I1(x2728), .I2(x2729), .I3(n11447), .I4(n11448), .O(n11451));
  LUT5 #(.INIT(32'hFF969600)) lut_n11452 (.I0(x2733), .I1(x2734), .I2(x2735), .I3(n11450), .I4(n11451), .O(n11452));
  LUT3 #(.INIT(8'h96)) lut_n11453 (.I0(n11441), .I1(n11444), .I2(n11445), .O(n11453));
  LUT3 #(.INIT(8'hE8)) lut_n11454 (.I0(n11449), .I1(n11452), .I2(n11453), .O(n11454));
  LUT3 #(.INIT(8'h96)) lut_n11455 (.I0(n11424), .I1(n11432), .I2(n11433), .O(n11455));
  LUT3 #(.INIT(8'hE8)) lut_n11456 (.I0(n11446), .I1(n11454), .I2(n11455), .O(n11456));
  LUT3 #(.INIT(8'h96)) lut_n11457 (.I0(x2742), .I1(x2743), .I2(x2744), .O(n11457));
  LUT5 #(.INIT(32'h96696996)) lut_n11458 (.I0(x2733), .I1(x2734), .I2(x2735), .I3(n11450), .I4(n11451), .O(n11458));
  LUT5 #(.INIT(32'hFF969600)) lut_n11459 (.I0(x2739), .I1(x2740), .I2(x2741), .I3(n11457), .I4(n11458), .O(n11459));
  LUT3 #(.INIT(8'h96)) lut_n11460 (.I0(x2748), .I1(x2749), .I2(x2750), .O(n11460));
  LUT5 #(.INIT(32'h96696996)) lut_n11461 (.I0(x2739), .I1(x2740), .I2(x2741), .I3(n11457), .I4(n11458), .O(n11461));
  LUT5 #(.INIT(32'hFF969600)) lut_n11462 (.I0(x2745), .I1(x2746), .I2(x2747), .I3(n11460), .I4(n11461), .O(n11462));
  LUT3 #(.INIT(8'h96)) lut_n11463 (.I0(n11449), .I1(n11452), .I2(n11453), .O(n11463));
  LUT3 #(.INIT(8'hE8)) lut_n11464 (.I0(n11459), .I1(n11462), .I2(n11463), .O(n11464));
  LUT3 #(.INIT(8'h96)) lut_n11465 (.I0(x2754), .I1(x2755), .I2(x2756), .O(n11465));
  LUT5 #(.INIT(32'h96696996)) lut_n11466 (.I0(x2745), .I1(x2746), .I2(x2747), .I3(n11460), .I4(n11461), .O(n11466));
  LUT5 #(.INIT(32'hFF969600)) lut_n11467 (.I0(x2751), .I1(x2752), .I2(x2753), .I3(n11465), .I4(n11466), .O(n11467));
  LUT3 #(.INIT(8'h96)) lut_n11468 (.I0(x2760), .I1(x2761), .I2(x2762), .O(n11468));
  LUT5 #(.INIT(32'h96696996)) lut_n11469 (.I0(x2751), .I1(x2752), .I2(x2753), .I3(n11465), .I4(n11466), .O(n11469));
  LUT5 #(.INIT(32'hFF969600)) lut_n11470 (.I0(x2757), .I1(x2758), .I2(x2759), .I3(n11468), .I4(n11469), .O(n11470));
  LUT3 #(.INIT(8'h96)) lut_n11471 (.I0(n11459), .I1(n11462), .I2(n11463), .O(n11471));
  LUT3 #(.INIT(8'hE8)) lut_n11472 (.I0(n11467), .I1(n11470), .I2(n11471), .O(n11472));
  LUT3 #(.INIT(8'h96)) lut_n11473 (.I0(n11446), .I1(n11454), .I2(n11455), .O(n11473));
  LUT3 #(.INIT(8'hE8)) lut_n11474 (.I0(n11464), .I1(n11472), .I2(n11473), .O(n11474));
  LUT3 #(.INIT(8'h96)) lut_n11475 (.I0(n11416), .I1(n11434), .I2(n11435), .O(n11475));
  LUT3 #(.INIT(8'hE8)) lut_n11476 (.I0(n11456), .I1(n11474), .I2(n11475), .O(n11476));
  LUT3 #(.INIT(8'h96)) lut_n11477 (.I0(x2766), .I1(x2767), .I2(x2768), .O(n11477));
  LUT5 #(.INIT(32'h96696996)) lut_n11478 (.I0(x2757), .I1(x2758), .I2(x2759), .I3(n11468), .I4(n11469), .O(n11478));
  LUT5 #(.INIT(32'hFF969600)) lut_n11479 (.I0(x2763), .I1(x2764), .I2(x2765), .I3(n11477), .I4(n11478), .O(n11479));
  LUT3 #(.INIT(8'h96)) lut_n11480 (.I0(x2772), .I1(x2773), .I2(x2774), .O(n11480));
  LUT5 #(.INIT(32'h96696996)) lut_n11481 (.I0(x2763), .I1(x2764), .I2(x2765), .I3(n11477), .I4(n11478), .O(n11481));
  LUT5 #(.INIT(32'hFF969600)) lut_n11482 (.I0(x2769), .I1(x2770), .I2(x2771), .I3(n11480), .I4(n11481), .O(n11482));
  LUT3 #(.INIT(8'h96)) lut_n11483 (.I0(n11467), .I1(n11470), .I2(n11471), .O(n11483));
  LUT3 #(.INIT(8'hE8)) lut_n11484 (.I0(n11479), .I1(n11482), .I2(n11483), .O(n11484));
  LUT3 #(.INIT(8'h96)) lut_n11485 (.I0(x2778), .I1(x2779), .I2(x2780), .O(n11485));
  LUT5 #(.INIT(32'h96696996)) lut_n11486 (.I0(x2769), .I1(x2770), .I2(x2771), .I3(n11480), .I4(n11481), .O(n11486));
  LUT5 #(.INIT(32'hFF969600)) lut_n11487 (.I0(x2775), .I1(x2776), .I2(x2777), .I3(n11485), .I4(n11486), .O(n11487));
  LUT3 #(.INIT(8'h96)) lut_n11488 (.I0(x2784), .I1(x2785), .I2(x2786), .O(n11488));
  LUT5 #(.INIT(32'h96696996)) lut_n11489 (.I0(x2775), .I1(x2776), .I2(x2777), .I3(n11485), .I4(n11486), .O(n11489));
  LUT5 #(.INIT(32'hFF969600)) lut_n11490 (.I0(x2781), .I1(x2782), .I2(x2783), .I3(n11488), .I4(n11489), .O(n11490));
  LUT3 #(.INIT(8'h96)) lut_n11491 (.I0(n11479), .I1(n11482), .I2(n11483), .O(n11491));
  LUT3 #(.INIT(8'hE8)) lut_n11492 (.I0(n11487), .I1(n11490), .I2(n11491), .O(n11492));
  LUT3 #(.INIT(8'h96)) lut_n11493 (.I0(n11464), .I1(n11472), .I2(n11473), .O(n11493));
  LUT3 #(.INIT(8'hE8)) lut_n11494 (.I0(n11484), .I1(n11492), .I2(n11493), .O(n11494));
  LUT3 #(.INIT(8'h96)) lut_n11495 (.I0(x2790), .I1(x2791), .I2(x2792), .O(n11495));
  LUT5 #(.INIT(32'h96696996)) lut_n11496 (.I0(x2781), .I1(x2782), .I2(x2783), .I3(n11488), .I4(n11489), .O(n11496));
  LUT5 #(.INIT(32'hFF969600)) lut_n11497 (.I0(x2787), .I1(x2788), .I2(x2789), .I3(n11495), .I4(n11496), .O(n11497));
  LUT3 #(.INIT(8'h96)) lut_n11498 (.I0(x2796), .I1(x2797), .I2(x2798), .O(n11498));
  LUT5 #(.INIT(32'h96696996)) lut_n11499 (.I0(x2787), .I1(x2788), .I2(x2789), .I3(n11495), .I4(n11496), .O(n11499));
  LUT5 #(.INIT(32'hFF969600)) lut_n11500 (.I0(x2793), .I1(x2794), .I2(x2795), .I3(n11498), .I4(n11499), .O(n11500));
  LUT3 #(.INIT(8'h96)) lut_n11501 (.I0(n11487), .I1(n11490), .I2(n11491), .O(n11501));
  LUT3 #(.INIT(8'hE8)) lut_n11502 (.I0(n11497), .I1(n11500), .I2(n11501), .O(n11502));
  LUT3 #(.INIT(8'h96)) lut_n11503 (.I0(x2802), .I1(x2803), .I2(x2804), .O(n11503));
  LUT5 #(.INIT(32'h96696996)) lut_n11504 (.I0(x2793), .I1(x2794), .I2(x2795), .I3(n11498), .I4(n11499), .O(n11504));
  LUT5 #(.INIT(32'hFF969600)) lut_n11505 (.I0(x2799), .I1(x2800), .I2(x2801), .I3(n11503), .I4(n11504), .O(n11505));
  LUT3 #(.INIT(8'h96)) lut_n11506 (.I0(x2808), .I1(x2809), .I2(x2810), .O(n11506));
  LUT5 #(.INIT(32'h96696996)) lut_n11507 (.I0(x2799), .I1(x2800), .I2(x2801), .I3(n11503), .I4(n11504), .O(n11507));
  LUT5 #(.INIT(32'hFF969600)) lut_n11508 (.I0(x2805), .I1(x2806), .I2(x2807), .I3(n11506), .I4(n11507), .O(n11508));
  LUT3 #(.INIT(8'h96)) lut_n11509 (.I0(n11497), .I1(n11500), .I2(n11501), .O(n11509));
  LUT3 #(.INIT(8'hE8)) lut_n11510 (.I0(n11505), .I1(n11508), .I2(n11509), .O(n11510));
  LUT3 #(.INIT(8'h96)) lut_n11511 (.I0(n11484), .I1(n11492), .I2(n11493), .O(n11511));
  LUT3 #(.INIT(8'hE8)) lut_n11512 (.I0(n11502), .I1(n11510), .I2(n11511), .O(n11512));
  LUT3 #(.INIT(8'h96)) lut_n11513 (.I0(n11456), .I1(n11474), .I2(n11475), .O(n11513));
  LUT3 #(.INIT(8'hE8)) lut_n11514 (.I0(n11494), .I1(n11512), .I2(n11513), .O(n11514));
  LUT3 #(.INIT(8'h96)) lut_n11515 (.I0(n11398), .I1(n11436), .I2(n11437), .O(n11515));
  LUT3 #(.INIT(8'hE8)) lut_n11516 (.I0(n11476), .I1(n11514), .I2(n11515), .O(n11516));
  LUT3 #(.INIT(8'h96)) lut_n11517 (.I0(n11278), .I1(n11356), .I2(n11357), .O(n11517));
  LUT3 #(.INIT(8'hE8)) lut_n11518 (.I0(n11438), .I1(n11516), .I2(n11517), .O(n11518));
  LUT3 #(.INIT(8'h96)) lut_n11519 (.I0(x2814), .I1(x2815), .I2(x2816), .O(n11519));
  LUT5 #(.INIT(32'h96696996)) lut_n11520 (.I0(x2805), .I1(x2806), .I2(x2807), .I3(n11506), .I4(n11507), .O(n11520));
  LUT5 #(.INIT(32'hFF969600)) lut_n11521 (.I0(x2811), .I1(x2812), .I2(x2813), .I3(n11519), .I4(n11520), .O(n11521));
  LUT3 #(.INIT(8'h96)) lut_n11522 (.I0(x2820), .I1(x2821), .I2(x2822), .O(n11522));
  LUT5 #(.INIT(32'h96696996)) lut_n11523 (.I0(x2811), .I1(x2812), .I2(x2813), .I3(n11519), .I4(n11520), .O(n11523));
  LUT5 #(.INIT(32'hFF969600)) lut_n11524 (.I0(x2817), .I1(x2818), .I2(x2819), .I3(n11522), .I4(n11523), .O(n11524));
  LUT3 #(.INIT(8'h96)) lut_n11525 (.I0(n11505), .I1(n11508), .I2(n11509), .O(n11525));
  LUT3 #(.INIT(8'hE8)) lut_n11526 (.I0(n11521), .I1(n11524), .I2(n11525), .O(n11526));
  LUT3 #(.INIT(8'h96)) lut_n11527 (.I0(x2826), .I1(x2827), .I2(x2828), .O(n11527));
  LUT5 #(.INIT(32'h96696996)) lut_n11528 (.I0(x2817), .I1(x2818), .I2(x2819), .I3(n11522), .I4(n11523), .O(n11528));
  LUT5 #(.INIT(32'hFF969600)) lut_n11529 (.I0(x2823), .I1(x2824), .I2(x2825), .I3(n11527), .I4(n11528), .O(n11529));
  LUT3 #(.INIT(8'h96)) lut_n11530 (.I0(x2832), .I1(x2833), .I2(x2834), .O(n11530));
  LUT5 #(.INIT(32'h96696996)) lut_n11531 (.I0(x2823), .I1(x2824), .I2(x2825), .I3(n11527), .I4(n11528), .O(n11531));
  LUT5 #(.INIT(32'hFF969600)) lut_n11532 (.I0(x2829), .I1(x2830), .I2(x2831), .I3(n11530), .I4(n11531), .O(n11532));
  LUT3 #(.INIT(8'h96)) lut_n11533 (.I0(n11521), .I1(n11524), .I2(n11525), .O(n11533));
  LUT3 #(.INIT(8'hE8)) lut_n11534 (.I0(n11529), .I1(n11532), .I2(n11533), .O(n11534));
  LUT3 #(.INIT(8'h96)) lut_n11535 (.I0(n11502), .I1(n11510), .I2(n11511), .O(n11535));
  LUT3 #(.INIT(8'hE8)) lut_n11536 (.I0(n11526), .I1(n11534), .I2(n11535), .O(n11536));
  LUT3 #(.INIT(8'h96)) lut_n11537 (.I0(x2838), .I1(x2839), .I2(x2840), .O(n11537));
  LUT5 #(.INIT(32'h96696996)) lut_n11538 (.I0(x2829), .I1(x2830), .I2(x2831), .I3(n11530), .I4(n11531), .O(n11538));
  LUT5 #(.INIT(32'hFF969600)) lut_n11539 (.I0(x2835), .I1(x2836), .I2(x2837), .I3(n11537), .I4(n11538), .O(n11539));
  LUT3 #(.INIT(8'h96)) lut_n11540 (.I0(x2844), .I1(x2845), .I2(x2846), .O(n11540));
  LUT5 #(.INIT(32'h96696996)) lut_n11541 (.I0(x2835), .I1(x2836), .I2(x2837), .I3(n11537), .I4(n11538), .O(n11541));
  LUT5 #(.INIT(32'hFF969600)) lut_n11542 (.I0(x2841), .I1(x2842), .I2(x2843), .I3(n11540), .I4(n11541), .O(n11542));
  LUT3 #(.INIT(8'h96)) lut_n11543 (.I0(n11529), .I1(n11532), .I2(n11533), .O(n11543));
  LUT3 #(.INIT(8'hE8)) lut_n11544 (.I0(n11539), .I1(n11542), .I2(n11543), .O(n11544));
  LUT3 #(.INIT(8'h96)) lut_n11545 (.I0(x2850), .I1(x2851), .I2(x2852), .O(n11545));
  LUT5 #(.INIT(32'h96696996)) lut_n11546 (.I0(x2841), .I1(x2842), .I2(x2843), .I3(n11540), .I4(n11541), .O(n11546));
  LUT5 #(.INIT(32'hFF969600)) lut_n11547 (.I0(x2847), .I1(x2848), .I2(x2849), .I3(n11545), .I4(n11546), .O(n11547));
  LUT3 #(.INIT(8'h96)) lut_n11548 (.I0(x2856), .I1(x2857), .I2(x2858), .O(n11548));
  LUT5 #(.INIT(32'h96696996)) lut_n11549 (.I0(x2847), .I1(x2848), .I2(x2849), .I3(n11545), .I4(n11546), .O(n11549));
  LUT5 #(.INIT(32'hFF969600)) lut_n11550 (.I0(x2853), .I1(x2854), .I2(x2855), .I3(n11548), .I4(n11549), .O(n11550));
  LUT3 #(.INIT(8'h96)) lut_n11551 (.I0(n11539), .I1(n11542), .I2(n11543), .O(n11551));
  LUT3 #(.INIT(8'hE8)) lut_n11552 (.I0(n11547), .I1(n11550), .I2(n11551), .O(n11552));
  LUT3 #(.INIT(8'h96)) lut_n11553 (.I0(n11526), .I1(n11534), .I2(n11535), .O(n11553));
  LUT3 #(.INIT(8'hE8)) lut_n11554 (.I0(n11544), .I1(n11552), .I2(n11553), .O(n11554));
  LUT3 #(.INIT(8'h96)) lut_n11555 (.I0(n11494), .I1(n11512), .I2(n11513), .O(n11555));
  LUT3 #(.INIT(8'hE8)) lut_n11556 (.I0(n11536), .I1(n11554), .I2(n11555), .O(n11556));
  LUT3 #(.INIT(8'h96)) lut_n11557 (.I0(x2862), .I1(x2863), .I2(x2864), .O(n11557));
  LUT5 #(.INIT(32'h96696996)) lut_n11558 (.I0(x2853), .I1(x2854), .I2(x2855), .I3(n11548), .I4(n11549), .O(n11558));
  LUT5 #(.INIT(32'hFF969600)) lut_n11559 (.I0(x2859), .I1(x2860), .I2(x2861), .I3(n11557), .I4(n11558), .O(n11559));
  LUT3 #(.INIT(8'h96)) lut_n11560 (.I0(x2868), .I1(x2869), .I2(x2870), .O(n11560));
  LUT5 #(.INIT(32'h96696996)) lut_n11561 (.I0(x2859), .I1(x2860), .I2(x2861), .I3(n11557), .I4(n11558), .O(n11561));
  LUT5 #(.INIT(32'hFF969600)) lut_n11562 (.I0(x2865), .I1(x2866), .I2(x2867), .I3(n11560), .I4(n11561), .O(n11562));
  LUT3 #(.INIT(8'h96)) lut_n11563 (.I0(n11547), .I1(n11550), .I2(n11551), .O(n11563));
  LUT3 #(.INIT(8'hE8)) lut_n11564 (.I0(n11559), .I1(n11562), .I2(n11563), .O(n11564));
  LUT3 #(.INIT(8'h96)) lut_n11565 (.I0(x2874), .I1(x2875), .I2(x2876), .O(n11565));
  LUT5 #(.INIT(32'h96696996)) lut_n11566 (.I0(x2865), .I1(x2866), .I2(x2867), .I3(n11560), .I4(n11561), .O(n11566));
  LUT5 #(.INIT(32'hFF969600)) lut_n11567 (.I0(x2871), .I1(x2872), .I2(x2873), .I3(n11565), .I4(n11566), .O(n11567));
  LUT3 #(.INIT(8'h96)) lut_n11568 (.I0(x2880), .I1(x2881), .I2(x2882), .O(n11568));
  LUT5 #(.INIT(32'h96696996)) lut_n11569 (.I0(x2871), .I1(x2872), .I2(x2873), .I3(n11565), .I4(n11566), .O(n11569));
  LUT5 #(.INIT(32'hFF969600)) lut_n11570 (.I0(x2877), .I1(x2878), .I2(x2879), .I3(n11568), .I4(n11569), .O(n11570));
  LUT3 #(.INIT(8'h96)) lut_n11571 (.I0(n11559), .I1(n11562), .I2(n11563), .O(n11571));
  LUT3 #(.INIT(8'hE8)) lut_n11572 (.I0(n11567), .I1(n11570), .I2(n11571), .O(n11572));
  LUT3 #(.INIT(8'h96)) lut_n11573 (.I0(n11544), .I1(n11552), .I2(n11553), .O(n11573));
  LUT3 #(.INIT(8'hE8)) lut_n11574 (.I0(n11564), .I1(n11572), .I2(n11573), .O(n11574));
  LUT3 #(.INIT(8'h96)) lut_n11575 (.I0(x2886), .I1(x2887), .I2(x2888), .O(n11575));
  LUT5 #(.INIT(32'h96696996)) lut_n11576 (.I0(x2877), .I1(x2878), .I2(x2879), .I3(n11568), .I4(n11569), .O(n11576));
  LUT5 #(.INIT(32'hFF969600)) lut_n11577 (.I0(x2883), .I1(x2884), .I2(x2885), .I3(n11575), .I4(n11576), .O(n11577));
  LUT3 #(.INIT(8'h96)) lut_n11578 (.I0(x2892), .I1(x2893), .I2(x2894), .O(n11578));
  LUT5 #(.INIT(32'h96696996)) lut_n11579 (.I0(x2883), .I1(x2884), .I2(x2885), .I3(n11575), .I4(n11576), .O(n11579));
  LUT5 #(.INIT(32'hFF969600)) lut_n11580 (.I0(x2889), .I1(x2890), .I2(x2891), .I3(n11578), .I4(n11579), .O(n11580));
  LUT3 #(.INIT(8'h96)) lut_n11581 (.I0(n11567), .I1(n11570), .I2(n11571), .O(n11581));
  LUT3 #(.INIT(8'hE8)) lut_n11582 (.I0(n11577), .I1(n11580), .I2(n11581), .O(n11582));
  LUT3 #(.INIT(8'h96)) lut_n11583 (.I0(x2898), .I1(x2899), .I2(x2900), .O(n11583));
  LUT5 #(.INIT(32'h96696996)) lut_n11584 (.I0(x2889), .I1(x2890), .I2(x2891), .I3(n11578), .I4(n11579), .O(n11584));
  LUT5 #(.INIT(32'hFF969600)) lut_n11585 (.I0(x2895), .I1(x2896), .I2(x2897), .I3(n11583), .I4(n11584), .O(n11585));
  LUT3 #(.INIT(8'h96)) lut_n11586 (.I0(x2904), .I1(x2905), .I2(x2906), .O(n11586));
  LUT5 #(.INIT(32'h96696996)) lut_n11587 (.I0(x2895), .I1(x2896), .I2(x2897), .I3(n11583), .I4(n11584), .O(n11587));
  LUT5 #(.INIT(32'hFF969600)) lut_n11588 (.I0(x2901), .I1(x2902), .I2(x2903), .I3(n11586), .I4(n11587), .O(n11588));
  LUT3 #(.INIT(8'h96)) lut_n11589 (.I0(n11577), .I1(n11580), .I2(n11581), .O(n11589));
  LUT3 #(.INIT(8'hE8)) lut_n11590 (.I0(n11585), .I1(n11588), .I2(n11589), .O(n11590));
  LUT3 #(.INIT(8'h96)) lut_n11591 (.I0(n11564), .I1(n11572), .I2(n11573), .O(n11591));
  LUT3 #(.INIT(8'hE8)) lut_n11592 (.I0(n11582), .I1(n11590), .I2(n11591), .O(n11592));
  LUT3 #(.INIT(8'h96)) lut_n11593 (.I0(n11536), .I1(n11554), .I2(n11555), .O(n11593));
  LUT3 #(.INIT(8'hE8)) lut_n11594 (.I0(n11574), .I1(n11592), .I2(n11593), .O(n11594));
  LUT3 #(.INIT(8'h96)) lut_n11595 (.I0(n11476), .I1(n11514), .I2(n11515), .O(n11595));
  LUT3 #(.INIT(8'hE8)) lut_n11596 (.I0(n11556), .I1(n11594), .I2(n11595), .O(n11596));
  LUT3 #(.INIT(8'h96)) lut_n11597 (.I0(x2910), .I1(x2911), .I2(x2912), .O(n11597));
  LUT5 #(.INIT(32'h96696996)) lut_n11598 (.I0(x2901), .I1(x2902), .I2(x2903), .I3(n11586), .I4(n11587), .O(n11598));
  LUT5 #(.INIT(32'hFF969600)) lut_n11599 (.I0(x2907), .I1(x2908), .I2(x2909), .I3(n11597), .I4(n11598), .O(n11599));
  LUT3 #(.INIT(8'h96)) lut_n11600 (.I0(x2916), .I1(x2917), .I2(x2918), .O(n11600));
  LUT5 #(.INIT(32'h96696996)) lut_n11601 (.I0(x2907), .I1(x2908), .I2(x2909), .I3(n11597), .I4(n11598), .O(n11601));
  LUT5 #(.INIT(32'hFF969600)) lut_n11602 (.I0(x2913), .I1(x2914), .I2(x2915), .I3(n11600), .I4(n11601), .O(n11602));
  LUT3 #(.INIT(8'h96)) lut_n11603 (.I0(n11585), .I1(n11588), .I2(n11589), .O(n11603));
  LUT3 #(.INIT(8'hE8)) lut_n11604 (.I0(n11599), .I1(n11602), .I2(n11603), .O(n11604));
  LUT3 #(.INIT(8'h96)) lut_n11605 (.I0(x2922), .I1(x2923), .I2(x2924), .O(n11605));
  LUT5 #(.INIT(32'h96696996)) lut_n11606 (.I0(x2913), .I1(x2914), .I2(x2915), .I3(n11600), .I4(n11601), .O(n11606));
  LUT5 #(.INIT(32'hFF969600)) lut_n11607 (.I0(x2919), .I1(x2920), .I2(x2921), .I3(n11605), .I4(n11606), .O(n11607));
  LUT3 #(.INIT(8'h96)) lut_n11608 (.I0(x2928), .I1(x2929), .I2(x2930), .O(n11608));
  LUT5 #(.INIT(32'h96696996)) lut_n11609 (.I0(x2919), .I1(x2920), .I2(x2921), .I3(n11605), .I4(n11606), .O(n11609));
  LUT5 #(.INIT(32'hFF969600)) lut_n11610 (.I0(x2925), .I1(x2926), .I2(x2927), .I3(n11608), .I4(n11609), .O(n11610));
  LUT3 #(.INIT(8'h96)) lut_n11611 (.I0(n11599), .I1(n11602), .I2(n11603), .O(n11611));
  LUT3 #(.INIT(8'hE8)) lut_n11612 (.I0(n11607), .I1(n11610), .I2(n11611), .O(n11612));
  LUT3 #(.INIT(8'h96)) lut_n11613 (.I0(n11582), .I1(n11590), .I2(n11591), .O(n11613));
  LUT3 #(.INIT(8'hE8)) lut_n11614 (.I0(n11604), .I1(n11612), .I2(n11613), .O(n11614));
  LUT3 #(.INIT(8'h96)) lut_n11615 (.I0(x2934), .I1(x2935), .I2(x2936), .O(n11615));
  LUT5 #(.INIT(32'h96696996)) lut_n11616 (.I0(x2925), .I1(x2926), .I2(x2927), .I3(n11608), .I4(n11609), .O(n11616));
  LUT5 #(.INIT(32'hFF969600)) lut_n11617 (.I0(x2931), .I1(x2932), .I2(x2933), .I3(n11615), .I4(n11616), .O(n11617));
  LUT3 #(.INIT(8'h96)) lut_n11618 (.I0(x2940), .I1(x2941), .I2(x2942), .O(n11618));
  LUT5 #(.INIT(32'h96696996)) lut_n11619 (.I0(x2931), .I1(x2932), .I2(x2933), .I3(n11615), .I4(n11616), .O(n11619));
  LUT5 #(.INIT(32'hFF969600)) lut_n11620 (.I0(x2937), .I1(x2938), .I2(x2939), .I3(n11618), .I4(n11619), .O(n11620));
  LUT3 #(.INIT(8'h96)) lut_n11621 (.I0(n11607), .I1(n11610), .I2(n11611), .O(n11621));
  LUT3 #(.INIT(8'hE8)) lut_n11622 (.I0(n11617), .I1(n11620), .I2(n11621), .O(n11622));
  LUT3 #(.INIT(8'h96)) lut_n11623 (.I0(x2946), .I1(x2947), .I2(x2948), .O(n11623));
  LUT5 #(.INIT(32'h96696996)) lut_n11624 (.I0(x2937), .I1(x2938), .I2(x2939), .I3(n11618), .I4(n11619), .O(n11624));
  LUT5 #(.INIT(32'hFF969600)) lut_n11625 (.I0(x2943), .I1(x2944), .I2(x2945), .I3(n11623), .I4(n11624), .O(n11625));
  LUT3 #(.INIT(8'h96)) lut_n11626 (.I0(x2952), .I1(x2953), .I2(x2954), .O(n11626));
  LUT5 #(.INIT(32'h96696996)) lut_n11627 (.I0(x2943), .I1(x2944), .I2(x2945), .I3(n11623), .I4(n11624), .O(n11627));
  LUT5 #(.INIT(32'hFF969600)) lut_n11628 (.I0(x2949), .I1(x2950), .I2(x2951), .I3(n11626), .I4(n11627), .O(n11628));
  LUT3 #(.INIT(8'h96)) lut_n11629 (.I0(n11617), .I1(n11620), .I2(n11621), .O(n11629));
  LUT3 #(.INIT(8'hE8)) lut_n11630 (.I0(n11625), .I1(n11628), .I2(n11629), .O(n11630));
  LUT3 #(.INIT(8'h96)) lut_n11631 (.I0(n11604), .I1(n11612), .I2(n11613), .O(n11631));
  LUT3 #(.INIT(8'hE8)) lut_n11632 (.I0(n11622), .I1(n11630), .I2(n11631), .O(n11632));
  LUT3 #(.INIT(8'h96)) lut_n11633 (.I0(n11574), .I1(n11592), .I2(n11593), .O(n11633));
  LUT3 #(.INIT(8'hE8)) lut_n11634 (.I0(n11614), .I1(n11632), .I2(n11633), .O(n11634));
  LUT3 #(.INIT(8'h96)) lut_n11635 (.I0(x2958), .I1(x2959), .I2(x2960), .O(n11635));
  LUT5 #(.INIT(32'h96696996)) lut_n11636 (.I0(x2949), .I1(x2950), .I2(x2951), .I3(n11626), .I4(n11627), .O(n11636));
  LUT5 #(.INIT(32'hFF969600)) lut_n11637 (.I0(x2955), .I1(x2956), .I2(x2957), .I3(n11635), .I4(n11636), .O(n11637));
  LUT3 #(.INIT(8'h96)) lut_n11638 (.I0(x2964), .I1(x2965), .I2(x2966), .O(n11638));
  LUT5 #(.INIT(32'h96696996)) lut_n11639 (.I0(x2955), .I1(x2956), .I2(x2957), .I3(n11635), .I4(n11636), .O(n11639));
  LUT5 #(.INIT(32'hFF969600)) lut_n11640 (.I0(x2961), .I1(x2962), .I2(x2963), .I3(n11638), .I4(n11639), .O(n11640));
  LUT3 #(.INIT(8'h96)) lut_n11641 (.I0(n11625), .I1(n11628), .I2(n11629), .O(n11641));
  LUT3 #(.INIT(8'hE8)) lut_n11642 (.I0(n11637), .I1(n11640), .I2(n11641), .O(n11642));
  LUT3 #(.INIT(8'h96)) lut_n11643 (.I0(x2970), .I1(x2971), .I2(x2972), .O(n11643));
  LUT5 #(.INIT(32'h96696996)) lut_n11644 (.I0(x2961), .I1(x2962), .I2(x2963), .I3(n11638), .I4(n11639), .O(n11644));
  LUT5 #(.INIT(32'hFF969600)) lut_n11645 (.I0(x2967), .I1(x2968), .I2(x2969), .I3(n11643), .I4(n11644), .O(n11645));
  LUT3 #(.INIT(8'h96)) lut_n11646 (.I0(x2976), .I1(x2977), .I2(x2978), .O(n11646));
  LUT5 #(.INIT(32'h96696996)) lut_n11647 (.I0(x2967), .I1(x2968), .I2(x2969), .I3(n11643), .I4(n11644), .O(n11647));
  LUT5 #(.INIT(32'hFF969600)) lut_n11648 (.I0(x2973), .I1(x2974), .I2(x2975), .I3(n11646), .I4(n11647), .O(n11648));
  LUT3 #(.INIT(8'h96)) lut_n11649 (.I0(n11637), .I1(n11640), .I2(n11641), .O(n11649));
  LUT3 #(.INIT(8'hE8)) lut_n11650 (.I0(n11645), .I1(n11648), .I2(n11649), .O(n11650));
  LUT3 #(.INIT(8'h96)) lut_n11651 (.I0(n11622), .I1(n11630), .I2(n11631), .O(n11651));
  LUT3 #(.INIT(8'hE8)) lut_n11652 (.I0(n11642), .I1(n11650), .I2(n11651), .O(n11652));
  LUT3 #(.INIT(8'h96)) lut_n11653 (.I0(x2982), .I1(x2983), .I2(x2984), .O(n11653));
  LUT5 #(.INIT(32'h96696996)) lut_n11654 (.I0(x2973), .I1(x2974), .I2(x2975), .I3(n11646), .I4(n11647), .O(n11654));
  LUT5 #(.INIT(32'hFF969600)) lut_n11655 (.I0(x2979), .I1(x2980), .I2(x2981), .I3(n11653), .I4(n11654), .O(n11655));
  LUT3 #(.INIT(8'h96)) lut_n11656 (.I0(x2988), .I1(x2989), .I2(x2990), .O(n11656));
  LUT5 #(.INIT(32'h96696996)) lut_n11657 (.I0(x2979), .I1(x2980), .I2(x2981), .I3(n11653), .I4(n11654), .O(n11657));
  LUT5 #(.INIT(32'hFF969600)) lut_n11658 (.I0(x2985), .I1(x2986), .I2(x2987), .I3(n11656), .I4(n11657), .O(n11658));
  LUT3 #(.INIT(8'h96)) lut_n11659 (.I0(n11645), .I1(n11648), .I2(n11649), .O(n11659));
  LUT3 #(.INIT(8'hE8)) lut_n11660 (.I0(n11655), .I1(n11658), .I2(n11659), .O(n11660));
  LUT3 #(.INIT(8'h96)) lut_n11661 (.I0(x2994), .I1(x2995), .I2(x2996), .O(n11661));
  LUT5 #(.INIT(32'h96696996)) lut_n11662 (.I0(x2985), .I1(x2986), .I2(x2987), .I3(n11656), .I4(n11657), .O(n11662));
  LUT5 #(.INIT(32'hFF969600)) lut_n11663 (.I0(x2991), .I1(x2992), .I2(x2993), .I3(n11661), .I4(n11662), .O(n11663));
  LUT3 #(.INIT(8'h96)) lut_n11664 (.I0(x2997), .I1(x2998), .I2(x2999), .O(n11664));
  LUT5 #(.INIT(32'h96696996)) lut_n11665 (.I0(x2991), .I1(x2992), .I2(x2993), .I3(n11661), .I4(n11662), .O(n11665));
  LUT5 #(.INIT(32'hFF969600)) lut_n11666 (.I0(x3000), .I1(x3001), .I2(x3002), .I3(n11664), .I4(n11665), .O(n11666));
  LUT3 #(.INIT(8'h96)) lut_n11667 (.I0(n11655), .I1(n11658), .I2(n11659), .O(n11667));
  LUT3 #(.INIT(8'hE8)) lut_n11668 (.I0(n11663), .I1(n11666), .I2(n11667), .O(n11668));
  LUT3 #(.INIT(8'h96)) lut_n11669 (.I0(n11642), .I1(n11650), .I2(n11651), .O(n11669));
  LUT3 #(.INIT(8'hE8)) lut_n11670 (.I0(n11660), .I1(n11668), .I2(n11669), .O(n11670));
  LUT3 #(.INIT(8'h96)) lut_n11671 (.I0(n11614), .I1(n11632), .I2(n11633), .O(n11671));
  LUT3 #(.INIT(8'hE8)) lut_n11672 (.I0(n11652), .I1(n11670), .I2(n11671), .O(n11672));
  LUT3 #(.INIT(8'h96)) lut_n11673 (.I0(n11556), .I1(n11594), .I2(n11595), .O(n11673));
  LUT3 #(.INIT(8'hE8)) lut_n11674 (.I0(n11634), .I1(n11672), .I2(n11673), .O(n11674));
  LUT3 #(.INIT(8'h96)) lut_n11675 (.I0(n11438), .I1(n11516), .I2(n11517), .O(n11675));
  LUT3 #(.INIT(8'hE8)) lut_n11676 (.I0(n11596), .I1(n11674), .I2(n11675), .O(n11676));
  LUT3 #(.INIT(8'h96)) lut_n11677 (.I0(n11200), .I1(n11358), .I2(n11359), .O(n11677));
  LUT3 #(.INIT(8'hE8)) lut_n11678 (.I0(n11518), .I1(n11676), .I2(n11677), .O(n11678));
  LUT3 #(.INIT(8'h96)) lut_n11679 (.I0(n10717), .I1(n11035), .I2(n11036), .O(n11679));
  LUT3 #(.INIT(8'hE8)) lut_n11680 (.I0(n11360), .I1(n11678), .I2(n11679), .O(n11680));
  LUT3 #(.INIT(8'h96)) lut_n11681 (.I0(x3006), .I1(x3007), .I2(x3008), .O(n11681));
  LUT5 #(.INIT(32'h96696996)) lut_n11682 (.I0(x3000), .I1(x3001), .I2(x3002), .I3(n11664), .I4(n11665), .O(n11682));
  LUT5 #(.INIT(32'hFF969600)) lut_n11683 (.I0(x3003), .I1(x3004), .I2(x3005), .I3(n11681), .I4(n11682), .O(n11683));
  LUT3 #(.INIT(8'h96)) lut_n11684 (.I0(x3012), .I1(x3013), .I2(x3014), .O(n11684));
  LUT5 #(.INIT(32'h96696996)) lut_n11685 (.I0(x3003), .I1(x3004), .I2(x3005), .I3(n11681), .I4(n11682), .O(n11685));
  LUT5 #(.INIT(32'hFF969600)) lut_n11686 (.I0(x3009), .I1(x3010), .I2(x3011), .I3(n11684), .I4(n11685), .O(n11686));
  LUT3 #(.INIT(8'h96)) lut_n11687 (.I0(n11663), .I1(n11666), .I2(n11667), .O(n11687));
  LUT3 #(.INIT(8'hE8)) lut_n11688 (.I0(n11683), .I1(n11686), .I2(n11687), .O(n11688));
  LUT3 #(.INIT(8'h96)) lut_n11689 (.I0(x3018), .I1(x3019), .I2(x3020), .O(n11689));
  LUT5 #(.INIT(32'h96696996)) lut_n11690 (.I0(x3009), .I1(x3010), .I2(x3011), .I3(n11684), .I4(n11685), .O(n11690));
  LUT5 #(.INIT(32'hFF969600)) lut_n11691 (.I0(x3015), .I1(x3016), .I2(x3017), .I3(n11689), .I4(n11690), .O(n11691));
  LUT3 #(.INIT(8'h96)) lut_n11692 (.I0(x3024), .I1(x3025), .I2(x3026), .O(n11692));
  LUT5 #(.INIT(32'h96696996)) lut_n11693 (.I0(x3015), .I1(x3016), .I2(x3017), .I3(n11689), .I4(n11690), .O(n11693));
  LUT5 #(.INIT(32'hFF969600)) lut_n11694 (.I0(x3021), .I1(x3022), .I2(x3023), .I3(n11692), .I4(n11693), .O(n11694));
  LUT3 #(.INIT(8'h96)) lut_n11695 (.I0(n11683), .I1(n11686), .I2(n11687), .O(n11695));
  LUT3 #(.INIT(8'hE8)) lut_n11696 (.I0(n11691), .I1(n11694), .I2(n11695), .O(n11696));
  LUT3 #(.INIT(8'h96)) lut_n11697 (.I0(n11660), .I1(n11668), .I2(n11669), .O(n11697));
  LUT3 #(.INIT(8'hE8)) lut_n11698 (.I0(n11688), .I1(n11696), .I2(n11697), .O(n11698));
  LUT3 #(.INIT(8'h96)) lut_n11699 (.I0(x3030), .I1(x3031), .I2(x3032), .O(n11699));
  LUT5 #(.INIT(32'h96696996)) lut_n11700 (.I0(x3021), .I1(x3022), .I2(x3023), .I3(n11692), .I4(n11693), .O(n11700));
  LUT5 #(.INIT(32'hFF969600)) lut_n11701 (.I0(x3027), .I1(x3028), .I2(x3029), .I3(n11699), .I4(n11700), .O(n11701));
  LUT3 #(.INIT(8'h96)) lut_n11702 (.I0(x3036), .I1(x3037), .I2(x3038), .O(n11702));
  LUT5 #(.INIT(32'h96696996)) lut_n11703 (.I0(x3027), .I1(x3028), .I2(x3029), .I3(n11699), .I4(n11700), .O(n11703));
  LUT5 #(.INIT(32'hFF969600)) lut_n11704 (.I0(x3033), .I1(x3034), .I2(x3035), .I3(n11702), .I4(n11703), .O(n11704));
  LUT3 #(.INIT(8'h96)) lut_n11705 (.I0(n11691), .I1(n11694), .I2(n11695), .O(n11705));
  LUT3 #(.INIT(8'hE8)) lut_n11706 (.I0(n11701), .I1(n11704), .I2(n11705), .O(n11706));
  LUT3 #(.INIT(8'h96)) lut_n11707 (.I0(x3042), .I1(x3043), .I2(x3044), .O(n11707));
  LUT5 #(.INIT(32'h96696996)) lut_n11708 (.I0(x3033), .I1(x3034), .I2(x3035), .I3(n11702), .I4(n11703), .O(n11708));
  LUT5 #(.INIT(32'hFF969600)) lut_n11709 (.I0(x3039), .I1(x3040), .I2(x3041), .I3(n11707), .I4(n11708), .O(n11709));
  LUT3 #(.INIT(8'h96)) lut_n11710 (.I0(x3048), .I1(x3049), .I2(x3050), .O(n11710));
  LUT5 #(.INIT(32'h96696996)) lut_n11711 (.I0(x3039), .I1(x3040), .I2(x3041), .I3(n11707), .I4(n11708), .O(n11711));
  LUT5 #(.INIT(32'hFF969600)) lut_n11712 (.I0(x3045), .I1(x3046), .I2(x3047), .I3(n11710), .I4(n11711), .O(n11712));
  LUT3 #(.INIT(8'h96)) lut_n11713 (.I0(n11701), .I1(n11704), .I2(n11705), .O(n11713));
  LUT3 #(.INIT(8'hE8)) lut_n11714 (.I0(n11709), .I1(n11712), .I2(n11713), .O(n11714));
  LUT3 #(.INIT(8'h96)) lut_n11715 (.I0(n11688), .I1(n11696), .I2(n11697), .O(n11715));
  LUT3 #(.INIT(8'hE8)) lut_n11716 (.I0(n11706), .I1(n11714), .I2(n11715), .O(n11716));
  LUT3 #(.INIT(8'h96)) lut_n11717 (.I0(n11652), .I1(n11670), .I2(n11671), .O(n11717));
  LUT3 #(.INIT(8'hE8)) lut_n11718 (.I0(n11698), .I1(n11716), .I2(n11717), .O(n11718));
  LUT3 #(.INIT(8'h96)) lut_n11719 (.I0(x3054), .I1(x3055), .I2(x3056), .O(n11719));
  LUT5 #(.INIT(32'h96696996)) lut_n11720 (.I0(x3045), .I1(x3046), .I2(x3047), .I3(n11710), .I4(n11711), .O(n11720));
  LUT5 #(.INIT(32'hFF969600)) lut_n11721 (.I0(x3051), .I1(x3052), .I2(x3053), .I3(n11719), .I4(n11720), .O(n11721));
  LUT3 #(.INIT(8'h96)) lut_n11722 (.I0(x3060), .I1(x3061), .I2(x3062), .O(n11722));
  LUT5 #(.INIT(32'h96696996)) lut_n11723 (.I0(x3051), .I1(x3052), .I2(x3053), .I3(n11719), .I4(n11720), .O(n11723));
  LUT5 #(.INIT(32'hFF969600)) lut_n11724 (.I0(x3057), .I1(x3058), .I2(x3059), .I3(n11722), .I4(n11723), .O(n11724));
  LUT3 #(.INIT(8'h96)) lut_n11725 (.I0(n11709), .I1(n11712), .I2(n11713), .O(n11725));
  LUT3 #(.INIT(8'hE8)) lut_n11726 (.I0(n11721), .I1(n11724), .I2(n11725), .O(n11726));
  LUT3 #(.INIT(8'h96)) lut_n11727 (.I0(x3066), .I1(x3067), .I2(x3068), .O(n11727));
  LUT5 #(.INIT(32'h96696996)) lut_n11728 (.I0(x3057), .I1(x3058), .I2(x3059), .I3(n11722), .I4(n11723), .O(n11728));
  LUT5 #(.INIT(32'hFF969600)) lut_n11729 (.I0(x3063), .I1(x3064), .I2(x3065), .I3(n11727), .I4(n11728), .O(n11729));
  LUT3 #(.INIT(8'h96)) lut_n11730 (.I0(x3072), .I1(x3073), .I2(x3074), .O(n11730));
  LUT5 #(.INIT(32'h96696996)) lut_n11731 (.I0(x3063), .I1(x3064), .I2(x3065), .I3(n11727), .I4(n11728), .O(n11731));
  LUT5 #(.INIT(32'hFF969600)) lut_n11732 (.I0(x3069), .I1(x3070), .I2(x3071), .I3(n11730), .I4(n11731), .O(n11732));
  LUT3 #(.INIT(8'h96)) lut_n11733 (.I0(n11721), .I1(n11724), .I2(n11725), .O(n11733));
  LUT3 #(.INIT(8'hE8)) lut_n11734 (.I0(n11729), .I1(n11732), .I2(n11733), .O(n11734));
  LUT3 #(.INIT(8'h96)) lut_n11735 (.I0(n11706), .I1(n11714), .I2(n11715), .O(n11735));
  LUT3 #(.INIT(8'hE8)) lut_n11736 (.I0(n11726), .I1(n11734), .I2(n11735), .O(n11736));
  LUT3 #(.INIT(8'h96)) lut_n11737 (.I0(x3078), .I1(x3079), .I2(x3080), .O(n11737));
  LUT5 #(.INIT(32'h96696996)) lut_n11738 (.I0(x3069), .I1(x3070), .I2(x3071), .I3(n11730), .I4(n11731), .O(n11738));
  LUT5 #(.INIT(32'hFF969600)) lut_n11739 (.I0(x3075), .I1(x3076), .I2(x3077), .I3(n11737), .I4(n11738), .O(n11739));
  LUT3 #(.INIT(8'h96)) lut_n11740 (.I0(x3084), .I1(x3085), .I2(x3086), .O(n11740));
  LUT5 #(.INIT(32'h96696996)) lut_n11741 (.I0(x3075), .I1(x3076), .I2(x3077), .I3(n11737), .I4(n11738), .O(n11741));
  LUT5 #(.INIT(32'hFF969600)) lut_n11742 (.I0(x3081), .I1(x3082), .I2(x3083), .I3(n11740), .I4(n11741), .O(n11742));
  LUT3 #(.INIT(8'h96)) lut_n11743 (.I0(n11729), .I1(n11732), .I2(n11733), .O(n11743));
  LUT3 #(.INIT(8'hE8)) lut_n11744 (.I0(n11739), .I1(n11742), .I2(n11743), .O(n11744));
  LUT3 #(.INIT(8'h96)) lut_n11745 (.I0(x3090), .I1(x3091), .I2(x3092), .O(n11745));
  LUT5 #(.INIT(32'h96696996)) lut_n11746 (.I0(x3081), .I1(x3082), .I2(x3083), .I3(n11740), .I4(n11741), .O(n11746));
  LUT5 #(.INIT(32'hFF969600)) lut_n11747 (.I0(x3087), .I1(x3088), .I2(x3089), .I3(n11745), .I4(n11746), .O(n11747));
  LUT3 #(.INIT(8'h96)) lut_n11748 (.I0(x3096), .I1(x3097), .I2(x3098), .O(n11748));
  LUT5 #(.INIT(32'h96696996)) lut_n11749 (.I0(x3087), .I1(x3088), .I2(x3089), .I3(n11745), .I4(n11746), .O(n11749));
  LUT5 #(.INIT(32'hFF969600)) lut_n11750 (.I0(x3093), .I1(x3094), .I2(x3095), .I3(n11748), .I4(n11749), .O(n11750));
  LUT3 #(.INIT(8'h96)) lut_n11751 (.I0(n11739), .I1(n11742), .I2(n11743), .O(n11751));
  LUT3 #(.INIT(8'hE8)) lut_n11752 (.I0(n11747), .I1(n11750), .I2(n11751), .O(n11752));
  LUT3 #(.INIT(8'h96)) lut_n11753 (.I0(n11726), .I1(n11734), .I2(n11735), .O(n11753));
  LUT3 #(.INIT(8'hE8)) lut_n11754 (.I0(n11744), .I1(n11752), .I2(n11753), .O(n11754));
  LUT3 #(.INIT(8'h96)) lut_n11755 (.I0(n11698), .I1(n11716), .I2(n11717), .O(n11755));
  LUT3 #(.INIT(8'hE8)) lut_n11756 (.I0(n11736), .I1(n11754), .I2(n11755), .O(n11756));
  LUT3 #(.INIT(8'h96)) lut_n11757 (.I0(n11634), .I1(n11672), .I2(n11673), .O(n11757));
  LUT3 #(.INIT(8'hE8)) lut_n11758 (.I0(n11718), .I1(n11756), .I2(n11757), .O(n11758));
  LUT3 #(.INIT(8'h96)) lut_n11759 (.I0(x3102), .I1(x3103), .I2(x3104), .O(n11759));
  LUT5 #(.INIT(32'h96696996)) lut_n11760 (.I0(x3093), .I1(x3094), .I2(x3095), .I3(n11748), .I4(n11749), .O(n11760));
  LUT5 #(.INIT(32'hFF969600)) lut_n11761 (.I0(x3099), .I1(x3100), .I2(x3101), .I3(n11759), .I4(n11760), .O(n11761));
  LUT3 #(.INIT(8'h96)) lut_n11762 (.I0(x3108), .I1(x3109), .I2(x3110), .O(n11762));
  LUT5 #(.INIT(32'h96696996)) lut_n11763 (.I0(x3099), .I1(x3100), .I2(x3101), .I3(n11759), .I4(n11760), .O(n11763));
  LUT5 #(.INIT(32'hFF969600)) lut_n11764 (.I0(x3105), .I1(x3106), .I2(x3107), .I3(n11762), .I4(n11763), .O(n11764));
  LUT3 #(.INIT(8'h96)) lut_n11765 (.I0(n11747), .I1(n11750), .I2(n11751), .O(n11765));
  LUT3 #(.INIT(8'hE8)) lut_n11766 (.I0(n11761), .I1(n11764), .I2(n11765), .O(n11766));
  LUT3 #(.INIT(8'h96)) lut_n11767 (.I0(x3114), .I1(x3115), .I2(x3116), .O(n11767));
  LUT5 #(.INIT(32'h96696996)) lut_n11768 (.I0(x3105), .I1(x3106), .I2(x3107), .I3(n11762), .I4(n11763), .O(n11768));
  LUT5 #(.INIT(32'hFF969600)) lut_n11769 (.I0(x3111), .I1(x3112), .I2(x3113), .I3(n11767), .I4(n11768), .O(n11769));
  LUT3 #(.INIT(8'h96)) lut_n11770 (.I0(x3120), .I1(x3121), .I2(x3122), .O(n11770));
  LUT5 #(.INIT(32'h96696996)) lut_n11771 (.I0(x3111), .I1(x3112), .I2(x3113), .I3(n11767), .I4(n11768), .O(n11771));
  LUT5 #(.INIT(32'hFF969600)) lut_n11772 (.I0(x3117), .I1(x3118), .I2(x3119), .I3(n11770), .I4(n11771), .O(n11772));
  LUT3 #(.INIT(8'h96)) lut_n11773 (.I0(n11761), .I1(n11764), .I2(n11765), .O(n11773));
  LUT3 #(.INIT(8'hE8)) lut_n11774 (.I0(n11769), .I1(n11772), .I2(n11773), .O(n11774));
  LUT3 #(.INIT(8'h96)) lut_n11775 (.I0(n11744), .I1(n11752), .I2(n11753), .O(n11775));
  LUT3 #(.INIT(8'hE8)) lut_n11776 (.I0(n11766), .I1(n11774), .I2(n11775), .O(n11776));
  LUT3 #(.INIT(8'h96)) lut_n11777 (.I0(x3126), .I1(x3127), .I2(x3128), .O(n11777));
  LUT5 #(.INIT(32'h96696996)) lut_n11778 (.I0(x3117), .I1(x3118), .I2(x3119), .I3(n11770), .I4(n11771), .O(n11778));
  LUT5 #(.INIT(32'hFF969600)) lut_n11779 (.I0(x3123), .I1(x3124), .I2(x3125), .I3(n11777), .I4(n11778), .O(n11779));
  LUT3 #(.INIT(8'h96)) lut_n11780 (.I0(x3132), .I1(x3133), .I2(x3134), .O(n11780));
  LUT5 #(.INIT(32'h96696996)) lut_n11781 (.I0(x3123), .I1(x3124), .I2(x3125), .I3(n11777), .I4(n11778), .O(n11781));
  LUT5 #(.INIT(32'hFF969600)) lut_n11782 (.I0(x3129), .I1(x3130), .I2(x3131), .I3(n11780), .I4(n11781), .O(n11782));
  LUT3 #(.INIT(8'h96)) lut_n11783 (.I0(n11769), .I1(n11772), .I2(n11773), .O(n11783));
  LUT3 #(.INIT(8'hE8)) lut_n11784 (.I0(n11779), .I1(n11782), .I2(n11783), .O(n11784));
  LUT3 #(.INIT(8'h96)) lut_n11785 (.I0(x3138), .I1(x3139), .I2(x3140), .O(n11785));
  LUT5 #(.INIT(32'h96696996)) lut_n11786 (.I0(x3129), .I1(x3130), .I2(x3131), .I3(n11780), .I4(n11781), .O(n11786));
  LUT5 #(.INIT(32'hFF969600)) lut_n11787 (.I0(x3135), .I1(x3136), .I2(x3137), .I3(n11785), .I4(n11786), .O(n11787));
  LUT3 #(.INIT(8'h96)) lut_n11788 (.I0(x3144), .I1(x3145), .I2(x3146), .O(n11788));
  LUT5 #(.INIT(32'h96696996)) lut_n11789 (.I0(x3135), .I1(x3136), .I2(x3137), .I3(n11785), .I4(n11786), .O(n11789));
  LUT5 #(.INIT(32'hFF969600)) lut_n11790 (.I0(x3141), .I1(x3142), .I2(x3143), .I3(n11788), .I4(n11789), .O(n11790));
  LUT3 #(.INIT(8'h96)) lut_n11791 (.I0(n11779), .I1(n11782), .I2(n11783), .O(n11791));
  LUT3 #(.INIT(8'hE8)) lut_n11792 (.I0(n11787), .I1(n11790), .I2(n11791), .O(n11792));
  LUT3 #(.INIT(8'h96)) lut_n11793 (.I0(n11766), .I1(n11774), .I2(n11775), .O(n11793));
  LUT3 #(.INIT(8'hE8)) lut_n11794 (.I0(n11784), .I1(n11792), .I2(n11793), .O(n11794));
  LUT3 #(.INIT(8'h96)) lut_n11795 (.I0(n11736), .I1(n11754), .I2(n11755), .O(n11795));
  LUT3 #(.INIT(8'hE8)) lut_n11796 (.I0(n11776), .I1(n11794), .I2(n11795), .O(n11796));
  LUT3 #(.INIT(8'h96)) lut_n11797 (.I0(x3150), .I1(x3151), .I2(x3152), .O(n11797));
  LUT5 #(.INIT(32'h96696996)) lut_n11798 (.I0(x3141), .I1(x3142), .I2(x3143), .I3(n11788), .I4(n11789), .O(n11798));
  LUT5 #(.INIT(32'hFF969600)) lut_n11799 (.I0(x3147), .I1(x3148), .I2(x3149), .I3(n11797), .I4(n11798), .O(n11799));
  LUT3 #(.INIT(8'h96)) lut_n11800 (.I0(x3156), .I1(x3157), .I2(x3158), .O(n11800));
  LUT5 #(.INIT(32'h96696996)) lut_n11801 (.I0(x3147), .I1(x3148), .I2(x3149), .I3(n11797), .I4(n11798), .O(n11801));
  LUT5 #(.INIT(32'hFF969600)) lut_n11802 (.I0(x3153), .I1(x3154), .I2(x3155), .I3(n11800), .I4(n11801), .O(n11802));
  LUT3 #(.INIT(8'h96)) lut_n11803 (.I0(n11787), .I1(n11790), .I2(n11791), .O(n11803));
  LUT3 #(.INIT(8'hE8)) lut_n11804 (.I0(n11799), .I1(n11802), .I2(n11803), .O(n11804));
  LUT3 #(.INIT(8'h96)) lut_n11805 (.I0(x3162), .I1(x3163), .I2(x3164), .O(n11805));
  LUT5 #(.INIT(32'h96696996)) lut_n11806 (.I0(x3153), .I1(x3154), .I2(x3155), .I3(n11800), .I4(n11801), .O(n11806));
  LUT5 #(.INIT(32'hFF969600)) lut_n11807 (.I0(x3159), .I1(x3160), .I2(x3161), .I3(n11805), .I4(n11806), .O(n11807));
  LUT3 #(.INIT(8'h96)) lut_n11808 (.I0(x3168), .I1(x3169), .I2(x3170), .O(n11808));
  LUT5 #(.INIT(32'h96696996)) lut_n11809 (.I0(x3159), .I1(x3160), .I2(x3161), .I3(n11805), .I4(n11806), .O(n11809));
  LUT5 #(.INIT(32'hFF969600)) lut_n11810 (.I0(x3165), .I1(x3166), .I2(x3167), .I3(n11808), .I4(n11809), .O(n11810));
  LUT3 #(.INIT(8'h96)) lut_n11811 (.I0(n11799), .I1(n11802), .I2(n11803), .O(n11811));
  LUT3 #(.INIT(8'hE8)) lut_n11812 (.I0(n11807), .I1(n11810), .I2(n11811), .O(n11812));
  LUT3 #(.INIT(8'h96)) lut_n11813 (.I0(n11784), .I1(n11792), .I2(n11793), .O(n11813));
  LUT3 #(.INIT(8'hE8)) lut_n11814 (.I0(n11804), .I1(n11812), .I2(n11813), .O(n11814));
  LUT3 #(.INIT(8'h96)) lut_n11815 (.I0(x3174), .I1(x3175), .I2(x3176), .O(n11815));
  LUT5 #(.INIT(32'h96696996)) lut_n11816 (.I0(x3165), .I1(x3166), .I2(x3167), .I3(n11808), .I4(n11809), .O(n11816));
  LUT5 #(.INIT(32'hFF969600)) lut_n11817 (.I0(x3171), .I1(x3172), .I2(x3173), .I3(n11815), .I4(n11816), .O(n11817));
  LUT3 #(.INIT(8'h96)) lut_n11818 (.I0(x3180), .I1(x3181), .I2(x3182), .O(n11818));
  LUT5 #(.INIT(32'h96696996)) lut_n11819 (.I0(x3171), .I1(x3172), .I2(x3173), .I3(n11815), .I4(n11816), .O(n11819));
  LUT5 #(.INIT(32'hFF969600)) lut_n11820 (.I0(x3177), .I1(x3178), .I2(x3179), .I3(n11818), .I4(n11819), .O(n11820));
  LUT3 #(.INIT(8'h96)) lut_n11821 (.I0(n11807), .I1(n11810), .I2(n11811), .O(n11821));
  LUT3 #(.INIT(8'hE8)) lut_n11822 (.I0(n11817), .I1(n11820), .I2(n11821), .O(n11822));
  LUT3 #(.INIT(8'h96)) lut_n11823 (.I0(x3186), .I1(x3187), .I2(x3188), .O(n11823));
  LUT5 #(.INIT(32'h96696996)) lut_n11824 (.I0(x3177), .I1(x3178), .I2(x3179), .I3(n11818), .I4(n11819), .O(n11824));
  LUT5 #(.INIT(32'hFF969600)) lut_n11825 (.I0(x3183), .I1(x3184), .I2(x3185), .I3(n11823), .I4(n11824), .O(n11825));
  LUT3 #(.INIT(8'h96)) lut_n11826 (.I0(x3192), .I1(x3193), .I2(x3194), .O(n11826));
  LUT5 #(.INIT(32'h96696996)) lut_n11827 (.I0(x3183), .I1(x3184), .I2(x3185), .I3(n11823), .I4(n11824), .O(n11827));
  LUT5 #(.INIT(32'hFF969600)) lut_n11828 (.I0(x3189), .I1(x3190), .I2(x3191), .I3(n11826), .I4(n11827), .O(n11828));
  LUT3 #(.INIT(8'h96)) lut_n11829 (.I0(n11817), .I1(n11820), .I2(n11821), .O(n11829));
  LUT3 #(.INIT(8'hE8)) lut_n11830 (.I0(n11825), .I1(n11828), .I2(n11829), .O(n11830));
  LUT3 #(.INIT(8'h96)) lut_n11831 (.I0(n11804), .I1(n11812), .I2(n11813), .O(n11831));
  LUT3 #(.INIT(8'hE8)) lut_n11832 (.I0(n11822), .I1(n11830), .I2(n11831), .O(n11832));
  LUT3 #(.INIT(8'h96)) lut_n11833 (.I0(n11776), .I1(n11794), .I2(n11795), .O(n11833));
  LUT3 #(.INIT(8'hE8)) lut_n11834 (.I0(n11814), .I1(n11832), .I2(n11833), .O(n11834));
  LUT3 #(.INIT(8'h96)) lut_n11835 (.I0(n11718), .I1(n11756), .I2(n11757), .O(n11835));
  LUT3 #(.INIT(8'hE8)) lut_n11836 (.I0(n11796), .I1(n11834), .I2(n11835), .O(n11836));
  LUT3 #(.INIT(8'h96)) lut_n11837 (.I0(n11596), .I1(n11674), .I2(n11675), .O(n11837));
  LUT3 #(.INIT(8'hE8)) lut_n11838 (.I0(n11758), .I1(n11836), .I2(n11837), .O(n11838));
  LUT3 #(.INIT(8'h96)) lut_n11839 (.I0(x3198), .I1(x3199), .I2(x3200), .O(n11839));
  LUT5 #(.INIT(32'h96696996)) lut_n11840 (.I0(x3189), .I1(x3190), .I2(x3191), .I3(n11826), .I4(n11827), .O(n11840));
  LUT5 #(.INIT(32'hFF969600)) lut_n11841 (.I0(x3195), .I1(x3196), .I2(x3197), .I3(n11839), .I4(n11840), .O(n11841));
  LUT3 #(.INIT(8'h96)) lut_n11842 (.I0(x3204), .I1(x3205), .I2(x3206), .O(n11842));
  LUT5 #(.INIT(32'h96696996)) lut_n11843 (.I0(x3195), .I1(x3196), .I2(x3197), .I3(n11839), .I4(n11840), .O(n11843));
  LUT5 #(.INIT(32'hFF969600)) lut_n11844 (.I0(x3201), .I1(x3202), .I2(x3203), .I3(n11842), .I4(n11843), .O(n11844));
  LUT3 #(.INIT(8'h96)) lut_n11845 (.I0(n11825), .I1(n11828), .I2(n11829), .O(n11845));
  LUT3 #(.INIT(8'hE8)) lut_n11846 (.I0(n11841), .I1(n11844), .I2(n11845), .O(n11846));
  LUT3 #(.INIT(8'h96)) lut_n11847 (.I0(x3210), .I1(x3211), .I2(x3212), .O(n11847));
  LUT5 #(.INIT(32'h96696996)) lut_n11848 (.I0(x3201), .I1(x3202), .I2(x3203), .I3(n11842), .I4(n11843), .O(n11848));
  LUT5 #(.INIT(32'hFF969600)) lut_n11849 (.I0(x3207), .I1(x3208), .I2(x3209), .I3(n11847), .I4(n11848), .O(n11849));
  LUT3 #(.INIT(8'h96)) lut_n11850 (.I0(x3216), .I1(x3217), .I2(x3218), .O(n11850));
  LUT5 #(.INIT(32'h96696996)) lut_n11851 (.I0(x3207), .I1(x3208), .I2(x3209), .I3(n11847), .I4(n11848), .O(n11851));
  LUT5 #(.INIT(32'hFF969600)) lut_n11852 (.I0(x3213), .I1(x3214), .I2(x3215), .I3(n11850), .I4(n11851), .O(n11852));
  LUT3 #(.INIT(8'h96)) lut_n11853 (.I0(n11841), .I1(n11844), .I2(n11845), .O(n11853));
  LUT3 #(.INIT(8'hE8)) lut_n11854 (.I0(n11849), .I1(n11852), .I2(n11853), .O(n11854));
  LUT3 #(.INIT(8'h96)) lut_n11855 (.I0(n11822), .I1(n11830), .I2(n11831), .O(n11855));
  LUT3 #(.INIT(8'hE8)) lut_n11856 (.I0(n11846), .I1(n11854), .I2(n11855), .O(n11856));
  LUT3 #(.INIT(8'h96)) lut_n11857 (.I0(x3222), .I1(x3223), .I2(x3224), .O(n11857));
  LUT5 #(.INIT(32'h96696996)) lut_n11858 (.I0(x3213), .I1(x3214), .I2(x3215), .I3(n11850), .I4(n11851), .O(n11858));
  LUT5 #(.INIT(32'hFF969600)) lut_n11859 (.I0(x3219), .I1(x3220), .I2(x3221), .I3(n11857), .I4(n11858), .O(n11859));
  LUT3 #(.INIT(8'h96)) lut_n11860 (.I0(x3228), .I1(x3229), .I2(x3230), .O(n11860));
  LUT5 #(.INIT(32'h96696996)) lut_n11861 (.I0(x3219), .I1(x3220), .I2(x3221), .I3(n11857), .I4(n11858), .O(n11861));
  LUT5 #(.INIT(32'hFF969600)) lut_n11862 (.I0(x3225), .I1(x3226), .I2(x3227), .I3(n11860), .I4(n11861), .O(n11862));
  LUT3 #(.INIT(8'h96)) lut_n11863 (.I0(n11849), .I1(n11852), .I2(n11853), .O(n11863));
  LUT3 #(.INIT(8'hE8)) lut_n11864 (.I0(n11859), .I1(n11862), .I2(n11863), .O(n11864));
  LUT3 #(.INIT(8'h96)) lut_n11865 (.I0(x3234), .I1(x3235), .I2(x3236), .O(n11865));
  LUT5 #(.INIT(32'h96696996)) lut_n11866 (.I0(x3225), .I1(x3226), .I2(x3227), .I3(n11860), .I4(n11861), .O(n11866));
  LUT5 #(.INIT(32'hFF969600)) lut_n11867 (.I0(x3231), .I1(x3232), .I2(x3233), .I3(n11865), .I4(n11866), .O(n11867));
  LUT3 #(.INIT(8'h96)) lut_n11868 (.I0(x3240), .I1(x3241), .I2(x3242), .O(n11868));
  LUT5 #(.INIT(32'h96696996)) lut_n11869 (.I0(x3231), .I1(x3232), .I2(x3233), .I3(n11865), .I4(n11866), .O(n11869));
  LUT5 #(.INIT(32'hFF969600)) lut_n11870 (.I0(x3237), .I1(x3238), .I2(x3239), .I3(n11868), .I4(n11869), .O(n11870));
  LUT3 #(.INIT(8'h96)) lut_n11871 (.I0(n11859), .I1(n11862), .I2(n11863), .O(n11871));
  LUT3 #(.INIT(8'hE8)) lut_n11872 (.I0(n11867), .I1(n11870), .I2(n11871), .O(n11872));
  LUT3 #(.INIT(8'h96)) lut_n11873 (.I0(n11846), .I1(n11854), .I2(n11855), .O(n11873));
  LUT3 #(.INIT(8'hE8)) lut_n11874 (.I0(n11864), .I1(n11872), .I2(n11873), .O(n11874));
  LUT3 #(.INIT(8'h96)) lut_n11875 (.I0(n11814), .I1(n11832), .I2(n11833), .O(n11875));
  LUT3 #(.INIT(8'hE8)) lut_n11876 (.I0(n11856), .I1(n11874), .I2(n11875), .O(n11876));
  LUT3 #(.INIT(8'h96)) lut_n11877 (.I0(x3246), .I1(x3247), .I2(x3248), .O(n11877));
  LUT5 #(.INIT(32'h96696996)) lut_n11878 (.I0(x3237), .I1(x3238), .I2(x3239), .I3(n11868), .I4(n11869), .O(n11878));
  LUT5 #(.INIT(32'hFF969600)) lut_n11879 (.I0(x3243), .I1(x3244), .I2(x3245), .I3(n11877), .I4(n11878), .O(n11879));
  LUT3 #(.INIT(8'h96)) lut_n11880 (.I0(x3252), .I1(x3253), .I2(x3254), .O(n11880));
  LUT5 #(.INIT(32'h96696996)) lut_n11881 (.I0(x3243), .I1(x3244), .I2(x3245), .I3(n11877), .I4(n11878), .O(n11881));
  LUT5 #(.INIT(32'hFF969600)) lut_n11882 (.I0(x3249), .I1(x3250), .I2(x3251), .I3(n11880), .I4(n11881), .O(n11882));
  LUT3 #(.INIT(8'h96)) lut_n11883 (.I0(n11867), .I1(n11870), .I2(n11871), .O(n11883));
  LUT3 #(.INIT(8'hE8)) lut_n11884 (.I0(n11879), .I1(n11882), .I2(n11883), .O(n11884));
  LUT3 #(.INIT(8'h96)) lut_n11885 (.I0(x3258), .I1(x3259), .I2(x3260), .O(n11885));
  LUT5 #(.INIT(32'h96696996)) lut_n11886 (.I0(x3249), .I1(x3250), .I2(x3251), .I3(n11880), .I4(n11881), .O(n11886));
  LUT5 #(.INIT(32'hFF969600)) lut_n11887 (.I0(x3255), .I1(x3256), .I2(x3257), .I3(n11885), .I4(n11886), .O(n11887));
  LUT3 #(.INIT(8'h96)) lut_n11888 (.I0(x3264), .I1(x3265), .I2(x3266), .O(n11888));
  LUT5 #(.INIT(32'h96696996)) lut_n11889 (.I0(x3255), .I1(x3256), .I2(x3257), .I3(n11885), .I4(n11886), .O(n11889));
  LUT5 #(.INIT(32'hFF969600)) lut_n11890 (.I0(x3261), .I1(x3262), .I2(x3263), .I3(n11888), .I4(n11889), .O(n11890));
  LUT3 #(.INIT(8'h96)) lut_n11891 (.I0(n11879), .I1(n11882), .I2(n11883), .O(n11891));
  LUT3 #(.INIT(8'hE8)) lut_n11892 (.I0(n11887), .I1(n11890), .I2(n11891), .O(n11892));
  LUT3 #(.INIT(8'h96)) lut_n11893 (.I0(n11864), .I1(n11872), .I2(n11873), .O(n11893));
  LUT3 #(.INIT(8'hE8)) lut_n11894 (.I0(n11884), .I1(n11892), .I2(n11893), .O(n11894));
  LUT3 #(.INIT(8'h96)) lut_n11895 (.I0(x3270), .I1(x3271), .I2(x3272), .O(n11895));
  LUT5 #(.INIT(32'h96696996)) lut_n11896 (.I0(x3261), .I1(x3262), .I2(x3263), .I3(n11888), .I4(n11889), .O(n11896));
  LUT5 #(.INIT(32'hFF969600)) lut_n11897 (.I0(x3267), .I1(x3268), .I2(x3269), .I3(n11895), .I4(n11896), .O(n11897));
  LUT3 #(.INIT(8'h96)) lut_n11898 (.I0(x3276), .I1(x3277), .I2(x3278), .O(n11898));
  LUT5 #(.INIT(32'h96696996)) lut_n11899 (.I0(x3267), .I1(x3268), .I2(x3269), .I3(n11895), .I4(n11896), .O(n11899));
  LUT5 #(.INIT(32'hFF969600)) lut_n11900 (.I0(x3273), .I1(x3274), .I2(x3275), .I3(n11898), .I4(n11899), .O(n11900));
  LUT3 #(.INIT(8'h96)) lut_n11901 (.I0(n11887), .I1(n11890), .I2(n11891), .O(n11901));
  LUT3 #(.INIT(8'hE8)) lut_n11902 (.I0(n11897), .I1(n11900), .I2(n11901), .O(n11902));
  LUT3 #(.INIT(8'h96)) lut_n11903 (.I0(x3282), .I1(x3283), .I2(x3284), .O(n11903));
  LUT5 #(.INIT(32'h96696996)) lut_n11904 (.I0(x3273), .I1(x3274), .I2(x3275), .I3(n11898), .I4(n11899), .O(n11904));
  LUT5 #(.INIT(32'hFF969600)) lut_n11905 (.I0(x3279), .I1(x3280), .I2(x3281), .I3(n11903), .I4(n11904), .O(n11905));
  LUT3 #(.INIT(8'h96)) lut_n11906 (.I0(x3288), .I1(x3289), .I2(x3290), .O(n11906));
  LUT5 #(.INIT(32'h96696996)) lut_n11907 (.I0(x3279), .I1(x3280), .I2(x3281), .I3(n11903), .I4(n11904), .O(n11907));
  LUT5 #(.INIT(32'hFF969600)) lut_n11908 (.I0(x3285), .I1(x3286), .I2(x3287), .I3(n11906), .I4(n11907), .O(n11908));
  LUT3 #(.INIT(8'h96)) lut_n11909 (.I0(n11897), .I1(n11900), .I2(n11901), .O(n11909));
  LUT3 #(.INIT(8'hE8)) lut_n11910 (.I0(n11905), .I1(n11908), .I2(n11909), .O(n11910));
  LUT3 #(.INIT(8'h96)) lut_n11911 (.I0(n11884), .I1(n11892), .I2(n11893), .O(n11911));
  LUT3 #(.INIT(8'hE8)) lut_n11912 (.I0(n11902), .I1(n11910), .I2(n11911), .O(n11912));
  LUT3 #(.INIT(8'h96)) lut_n11913 (.I0(n11856), .I1(n11874), .I2(n11875), .O(n11913));
  LUT3 #(.INIT(8'hE8)) lut_n11914 (.I0(n11894), .I1(n11912), .I2(n11913), .O(n11914));
  LUT3 #(.INIT(8'h96)) lut_n11915 (.I0(n11796), .I1(n11834), .I2(n11835), .O(n11915));
  LUT3 #(.INIT(8'hE8)) lut_n11916 (.I0(n11876), .I1(n11914), .I2(n11915), .O(n11916));
  LUT3 #(.INIT(8'h96)) lut_n11917 (.I0(x3294), .I1(x3295), .I2(x3296), .O(n11917));
  LUT5 #(.INIT(32'h96696996)) lut_n11918 (.I0(x3285), .I1(x3286), .I2(x3287), .I3(n11906), .I4(n11907), .O(n11918));
  LUT5 #(.INIT(32'hFF969600)) lut_n11919 (.I0(x3291), .I1(x3292), .I2(x3293), .I3(n11917), .I4(n11918), .O(n11919));
  LUT3 #(.INIT(8'h96)) lut_n11920 (.I0(x3300), .I1(x3301), .I2(x3302), .O(n11920));
  LUT5 #(.INIT(32'h96696996)) lut_n11921 (.I0(x3291), .I1(x3292), .I2(x3293), .I3(n11917), .I4(n11918), .O(n11921));
  LUT5 #(.INIT(32'hFF969600)) lut_n11922 (.I0(x3297), .I1(x3298), .I2(x3299), .I3(n11920), .I4(n11921), .O(n11922));
  LUT3 #(.INIT(8'h96)) lut_n11923 (.I0(n11905), .I1(n11908), .I2(n11909), .O(n11923));
  LUT3 #(.INIT(8'hE8)) lut_n11924 (.I0(n11919), .I1(n11922), .I2(n11923), .O(n11924));
  LUT3 #(.INIT(8'h96)) lut_n11925 (.I0(x3306), .I1(x3307), .I2(x3308), .O(n11925));
  LUT5 #(.INIT(32'h96696996)) lut_n11926 (.I0(x3297), .I1(x3298), .I2(x3299), .I3(n11920), .I4(n11921), .O(n11926));
  LUT5 #(.INIT(32'hFF969600)) lut_n11927 (.I0(x3303), .I1(x3304), .I2(x3305), .I3(n11925), .I4(n11926), .O(n11927));
  LUT3 #(.INIT(8'h96)) lut_n11928 (.I0(x3312), .I1(x3313), .I2(x3314), .O(n11928));
  LUT5 #(.INIT(32'h96696996)) lut_n11929 (.I0(x3303), .I1(x3304), .I2(x3305), .I3(n11925), .I4(n11926), .O(n11929));
  LUT5 #(.INIT(32'hFF969600)) lut_n11930 (.I0(x3309), .I1(x3310), .I2(x3311), .I3(n11928), .I4(n11929), .O(n11930));
  LUT3 #(.INIT(8'h96)) lut_n11931 (.I0(n11919), .I1(n11922), .I2(n11923), .O(n11931));
  LUT3 #(.INIT(8'hE8)) lut_n11932 (.I0(n11927), .I1(n11930), .I2(n11931), .O(n11932));
  LUT3 #(.INIT(8'h96)) lut_n11933 (.I0(n11902), .I1(n11910), .I2(n11911), .O(n11933));
  LUT3 #(.INIT(8'hE8)) lut_n11934 (.I0(n11924), .I1(n11932), .I2(n11933), .O(n11934));
  LUT3 #(.INIT(8'h96)) lut_n11935 (.I0(x3318), .I1(x3319), .I2(x3320), .O(n11935));
  LUT5 #(.INIT(32'h96696996)) lut_n11936 (.I0(x3309), .I1(x3310), .I2(x3311), .I3(n11928), .I4(n11929), .O(n11936));
  LUT5 #(.INIT(32'hFF969600)) lut_n11937 (.I0(x3315), .I1(x3316), .I2(x3317), .I3(n11935), .I4(n11936), .O(n11937));
  LUT3 #(.INIT(8'h96)) lut_n11938 (.I0(x3324), .I1(x3325), .I2(x3326), .O(n11938));
  LUT5 #(.INIT(32'h96696996)) lut_n11939 (.I0(x3315), .I1(x3316), .I2(x3317), .I3(n11935), .I4(n11936), .O(n11939));
  LUT5 #(.INIT(32'hFF969600)) lut_n11940 (.I0(x3321), .I1(x3322), .I2(x3323), .I3(n11938), .I4(n11939), .O(n11940));
  LUT3 #(.INIT(8'h96)) lut_n11941 (.I0(n11927), .I1(n11930), .I2(n11931), .O(n11941));
  LUT3 #(.INIT(8'hE8)) lut_n11942 (.I0(n11937), .I1(n11940), .I2(n11941), .O(n11942));
  LUT3 #(.INIT(8'h96)) lut_n11943 (.I0(x3330), .I1(x3331), .I2(x3332), .O(n11943));
  LUT5 #(.INIT(32'h96696996)) lut_n11944 (.I0(x3321), .I1(x3322), .I2(x3323), .I3(n11938), .I4(n11939), .O(n11944));
  LUT5 #(.INIT(32'hFF969600)) lut_n11945 (.I0(x3327), .I1(x3328), .I2(x3329), .I3(n11943), .I4(n11944), .O(n11945));
  LUT3 #(.INIT(8'h96)) lut_n11946 (.I0(x3336), .I1(x3337), .I2(x3338), .O(n11946));
  LUT5 #(.INIT(32'h96696996)) lut_n11947 (.I0(x3327), .I1(x3328), .I2(x3329), .I3(n11943), .I4(n11944), .O(n11947));
  LUT5 #(.INIT(32'hFF969600)) lut_n11948 (.I0(x3333), .I1(x3334), .I2(x3335), .I3(n11946), .I4(n11947), .O(n11948));
  LUT3 #(.INIT(8'h96)) lut_n11949 (.I0(n11937), .I1(n11940), .I2(n11941), .O(n11949));
  LUT3 #(.INIT(8'hE8)) lut_n11950 (.I0(n11945), .I1(n11948), .I2(n11949), .O(n11950));
  LUT3 #(.INIT(8'h96)) lut_n11951 (.I0(n11924), .I1(n11932), .I2(n11933), .O(n11951));
  LUT3 #(.INIT(8'hE8)) lut_n11952 (.I0(n11942), .I1(n11950), .I2(n11951), .O(n11952));
  LUT3 #(.INIT(8'h96)) lut_n11953 (.I0(n11894), .I1(n11912), .I2(n11913), .O(n11953));
  LUT3 #(.INIT(8'hE8)) lut_n11954 (.I0(n11934), .I1(n11952), .I2(n11953), .O(n11954));
  LUT3 #(.INIT(8'h96)) lut_n11955 (.I0(x3342), .I1(x3343), .I2(x3344), .O(n11955));
  LUT5 #(.INIT(32'h96696996)) lut_n11956 (.I0(x3333), .I1(x3334), .I2(x3335), .I3(n11946), .I4(n11947), .O(n11956));
  LUT5 #(.INIT(32'hFF969600)) lut_n11957 (.I0(x3339), .I1(x3340), .I2(x3341), .I3(n11955), .I4(n11956), .O(n11957));
  LUT3 #(.INIT(8'h96)) lut_n11958 (.I0(x3348), .I1(x3349), .I2(x3350), .O(n11958));
  LUT5 #(.INIT(32'h96696996)) lut_n11959 (.I0(x3339), .I1(x3340), .I2(x3341), .I3(n11955), .I4(n11956), .O(n11959));
  LUT5 #(.INIT(32'hFF969600)) lut_n11960 (.I0(x3345), .I1(x3346), .I2(x3347), .I3(n11958), .I4(n11959), .O(n11960));
  LUT3 #(.INIT(8'h96)) lut_n11961 (.I0(n11945), .I1(n11948), .I2(n11949), .O(n11961));
  LUT3 #(.INIT(8'hE8)) lut_n11962 (.I0(n11957), .I1(n11960), .I2(n11961), .O(n11962));
  LUT3 #(.INIT(8'h96)) lut_n11963 (.I0(x3354), .I1(x3355), .I2(x3356), .O(n11963));
  LUT5 #(.INIT(32'h96696996)) lut_n11964 (.I0(x3345), .I1(x3346), .I2(x3347), .I3(n11958), .I4(n11959), .O(n11964));
  LUT5 #(.INIT(32'hFF969600)) lut_n11965 (.I0(x3351), .I1(x3352), .I2(x3353), .I3(n11963), .I4(n11964), .O(n11965));
  LUT3 #(.INIT(8'h96)) lut_n11966 (.I0(x3360), .I1(x3361), .I2(x3362), .O(n11966));
  LUT5 #(.INIT(32'h96696996)) lut_n11967 (.I0(x3351), .I1(x3352), .I2(x3353), .I3(n11963), .I4(n11964), .O(n11967));
  LUT5 #(.INIT(32'hFF969600)) lut_n11968 (.I0(x3357), .I1(x3358), .I2(x3359), .I3(n11966), .I4(n11967), .O(n11968));
  LUT3 #(.INIT(8'h96)) lut_n11969 (.I0(n11957), .I1(n11960), .I2(n11961), .O(n11969));
  LUT3 #(.INIT(8'hE8)) lut_n11970 (.I0(n11965), .I1(n11968), .I2(n11969), .O(n11970));
  LUT3 #(.INIT(8'h96)) lut_n11971 (.I0(n11942), .I1(n11950), .I2(n11951), .O(n11971));
  LUT3 #(.INIT(8'hE8)) lut_n11972 (.I0(n11962), .I1(n11970), .I2(n11971), .O(n11972));
  LUT3 #(.INIT(8'h96)) lut_n11973 (.I0(x3366), .I1(x3367), .I2(x3368), .O(n11973));
  LUT5 #(.INIT(32'h96696996)) lut_n11974 (.I0(x3357), .I1(x3358), .I2(x3359), .I3(n11966), .I4(n11967), .O(n11974));
  LUT5 #(.INIT(32'hFF969600)) lut_n11975 (.I0(x3363), .I1(x3364), .I2(x3365), .I3(n11973), .I4(n11974), .O(n11975));
  LUT3 #(.INIT(8'h96)) lut_n11976 (.I0(x3372), .I1(x3373), .I2(x3374), .O(n11976));
  LUT5 #(.INIT(32'h96696996)) lut_n11977 (.I0(x3363), .I1(x3364), .I2(x3365), .I3(n11973), .I4(n11974), .O(n11977));
  LUT5 #(.INIT(32'hFF969600)) lut_n11978 (.I0(x3369), .I1(x3370), .I2(x3371), .I3(n11976), .I4(n11977), .O(n11978));
  LUT3 #(.INIT(8'h96)) lut_n11979 (.I0(n11965), .I1(n11968), .I2(n11969), .O(n11979));
  LUT3 #(.INIT(8'hE8)) lut_n11980 (.I0(n11975), .I1(n11978), .I2(n11979), .O(n11980));
  LUT3 #(.INIT(8'h96)) lut_n11981 (.I0(x3378), .I1(x3379), .I2(x3380), .O(n11981));
  LUT5 #(.INIT(32'h96696996)) lut_n11982 (.I0(x3369), .I1(x3370), .I2(x3371), .I3(n11976), .I4(n11977), .O(n11982));
  LUT5 #(.INIT(32'hFF969600)) lut_n11983 (.I0(x3375), .I1(x3376), .I2(x3377), .I3(n11981), .I4(n11982), .O(n11983));
  LUT3 #(.INIT(8'h96)) lut_n11984 (.I0(x3384), .I1(x3385), .I2(x3386), .O(n11984));
  LUT5 #(.INIT(32'h96696996)) lut_n11985 (.I0(x3375), .I1(x3376), .I2(x3377), .I3(n11981), .I4(n11982), .O(n11985));
  LUT5 #(.INIT(32'hFF969600)) lut_n11986 (.I0(x3381), .I1(x3382), .I2(x3383), .I3(n11984), .I4(n11985), .O(n11986));
  LUT3 #(.INIT(8'h96)) lut_n11987 (.I0(n11975), .I1(n11978), .I2(n11979), .O(n11987));
  LUT3 #(.INIT(8'hE8)) lut_n11988 (.I0(n11983), .I1(n11986), .I2(n11987), .O(n11988));
  LUT3 #(.INIT(8'h96)) lut_n11989 (.I0(n11962), .I1(n11970), .I2(n11971), .O(n11989));
  LUT3 #(.INIT(8'hE8)) lut_n11990 (.I0(n11980), .I1(n11988), .I2(n11989), .O(n11990));
  LUT3 #(.INIT(8'h96)) lut_n11991 (.I0(n11934), .I1(n11952), .I2(n11953), .O(n11991));
  LUT3 #(.INIT(8'hE8)) lut_n11992 (.I0(n11972), .I1(n11990), .I2(n11991), .O(n11992));
  LUT3 #(.INIT(8'h96)) lut_n11993 (.I0(n11876), .I1(n11914), .I2(n11915), .O(n11993));
  LUT3 #(.INIT(8'hE8)) lut_n11994 (.I0(n11954), .I1(n11992), .I2(n11993), .O(n11994));
  LUT3 #(.INIT(8'h96)) lut_n11995 (.I0(n11758), .I1(n11836), .I2(n11837), .O(n11995));
  LUT3 #(.INIT(8'hE8)) lut_n11996 (.I0(n11916), .I1(n11994), .I2(n11995), .O(n11996));
  LUT3 #(.INIT(8'h96)) lut_n11997 (.I0(n11518), .I1(n11676), .I2(n11677), .O(n11997));
  LUT3 #(.INIT(8'hE8)) lut_n11998 (.I0(n11838), .I1(n11996), .I2(n11997), .O(n11998));
  LUT3 #(.INIT(8'h96)) lut_n11999 (.I0(x3390), .I1(x3391), .I2(x3392), .O(n11999));
  LUT5 #(.INIT(32'h96696996)) lut_n12000 (.I0(x3381), .I1(x3382), .I2(x3383), .I3(n11984), .I4(n11985), .O(n12000));
  LUT5 #(.INIT(32'hFF969600)) lut_n12001 (.I0(x3387), .I1(x3388), .I2(x3389), .I3(n11999), .I4(n12000), .O(n12001));
  LUT3 #(.INIT(8'h96)) lut_n12002 (.I0(x3396), .I1(x3397), .I2(x3398), .O(n12002));
  LUT5 #(.INIT(32'h96696996)) lut_n12003 (.I0(x3387), .I1(x3388), .I2(x3389), .I3(n11999), .I4(n12000), .O(n12003));
  LUT5 #(.INIT(32'hFF969600)) lut_n12004 (.I0(x3393), .I1(x3394), .I2(x3395), .I3(n12002), .I4(n12003), .O(n12004));
  LUT3 #(.INIT(8'h96)) lut_n12005 (.I0(n11983), .I1(n11986), .I2(n11987), .O(n12005));
  LUT3 #(.INIT(8'hE8)) lut_n12006 (.I0(n12001), .I1(n12004), .I2(n12005), .O(n12006));
  LUT3 #(.INIT(8'h96)) lut_n12007 (.I0(x3402), .I1(x3403), .I2(x3404), .O(n12007));
  LUT5 #(.INIT(32'h96696996)) lut_n12008 (.I0(x3393), .I1(x3394), .I2(x3395), .I3(n12002), .I4(n12003), .O(n12008));
  LUT5 #(.INIT(32'hFF969600)) lut_n12009 (.I0(x3399), .I1(x3400), .I2(x3401), .I3(n12007), .I4(n12008), .O(n12009));
  LUT3 #(.INIT(8'h96)) lut_n12010 (.I0(x3408), .I1(x3409), .I2(x3410), .O(n12010));
  LUT5 #(.INIT(32'h96696996)) lut_n12011 (.I0(x3399), .I1(x3400), .I2(x3401), .I3(n12007), .I4(n12008), .O(n12011));
  LUT5 #(.INIT(32'hFF969600)) lut_n12012 (.I0(x3405), .I1(x3406), .I2(x3407), .I3(n12010), .I4(n12011), .O(n12012));
  LUT3 #(.INIT(8'h96)) lut_n12013 (.I0(n12001), .I1(n12004), .I2(n12005), .O(n12013));
  LUT3 #(.INIT(8'hE8)) lut_n12014 (.I0(n12009), .I1(n12012), .I2(n12013), .O(n12014));
  LUT3 #(.INIT(8'h96)) lut_n12015 (.I0(n11980), .I1(n11988), .I2(n11989), .O(n12015));
  LUT3 #(.INIT(8'hE8)) lut_n12016 (.I0(n12006), .I1(n12014), .I2(n12015), .O(n12016));
  LUT3 #(.INIT(8'h96)) lut_n12017 (.I0(x3414), .I1(x3415), .I2(x3416), .O(n12017));
  LUT5 #(.INIT(32'h96696996)) lut_n12018 (.I0(x3405), .I1(x3406), .I2(x3407), .I3(n12010), .I4(n12011), .O(n12018));
  LUT5 #(.INIT(32'hFF969600)) lut_n12019 (.I0(x3411), .I1(x3412), .I2(x3413), .I3(n12017), .I4(n12018), .O(n12019));
  LUT3 #(.INIT(8'h96)) lut_n12020 (.I0(x3420), .I1(x3421), .I2(x3422), .O(n12020));
  LUT5 #(.INIT(32'h96696996)) lut_n12021 (.I0(x3411), .I1(x3412), .I2(x3413), .I3(n12017), .I4(n12018), .O(n12021));
  LUT5 #(.INIT(32'hFF969600)) lut_n12022 (.I0(x3417), .I1(x3418), .I2(x3419), .I3(n12020), .I4(n12021), .O(n12022));
  LUT3 #(.INIT(8'h96)) lut_n12023 (.I0(n12009), .I1(n12012), .I2(n12013), .O(n12023));
  LUT3 #(.INIT(8'hE8)) lut_n12024 (.I0(n12019), .I1(n12022), .I2(n12023), .O(n12024));
  LUT3 #(.INIT(8'h96)) lut_n12025 (.I0(x3426), .I1(x3427), .I2(x3428), .O(n12025));
  LUT5 #(.INIT(32'h96696996)) lut_n12026 (.I0(x3417), .I1(x3418), .I2(x3419), .I3(n12020), .I4(n12021), .O(n12026));
  LUT5 #(.INIT(32'hFF969600)) lut_n12027 (.I0(x3423), .I1(x3424), .I2(x3425), .I3(n12025), .I4(n12026), .O(n12027));
  LUT3 #(.INIT(8'h96)) lut_n12028 (.I0(x3432), .I1(x3433), .I2(x3434), .O(n12028));
  LUT5 #(.INIT(32'h96696996)) lut_n12029 (.I0(x3423), .I1(x3424), .I2(x3425), .I3(n12025), .I4(n12026), .O(n12029));
  LUT5 #(.INIT(32'hFF969600)) lut_n12030 (.I0(x3429), .I1(x3430), .I2(x3431), .I3(n12028), .I4(n12029), .O(n12030));
  LUT3 #(.INIT(8'h96)) lut_n12031 (.I0(n12019), .I1(n12022), .I2(n12023), .O(n12031));
  LUT3 #(.INIT(8'hE8)) lut_n12032 (.I0(n12027), .I1(n12030), .I2(n12031), .O(n12032));
  LUT3 #(.INIT(8'h96)) lut_n12033 (.I0(n12006), .I1(n12014), .I2(n12015), .O(n12033));
  LUT3 #(.INIT(8'hE8)) lut_n12034 (.I0(n12024), .I1(n12032), .I2(n12033), .O(n12034));
  LUT3 #(.INIT(8'h96)) lut_n12035 (.I0(n11972), .I1(n11990), .I2(n11991), .O(n12035));
  LUT3 #(.INIT(8'hE8)) lut_n12036 (.I0(n12016), .I1(n12034), .I2(n12035), .O(n12036));
  LUT3 #(.INIT(8'h96)) lut_n12037 (.I0(x3438), .I1(x3439), .I2(x3440), .O(n12037));
  LUT5 #(.INIT(32'h96696996)) lut_n12038 (.I0(x3429), .I1(x3430), .I2(x3431), .I3(n12028), .I4(n12029), .O(n12038));
  LUT5 #(.INIT(32'hFF969600)) lut_n12039 (.I0(x3435), .I1(x3436), .I2(x3437), .I3(n12037), .I4(n12038), .O(n12039));
  LUT3 #(.INIT(8'h96)) lut_n12040 (.I0(x3444), .I1(x3445), .I2(x3446), .O(n12040));
  LUT5 #(.INIT(32'h96696996)) lut_n12041 (.I0(x3435), .I1(x3436), .I2(x3437), .I3(n12037), .I4(n12038), .O(n12041));
  LUT5 #(.INIT(32'hFF969600)) lut_n12042 (.I0(x3441), .I1(x3442), .I2(x3443), .I3(n12040), .I4(n12041), .O(n12042));
  LUT3 #(.INIT(8'h96)) lut_n12043 (.I0(n12027), .I1(n12030), .I2(n12031), .O(n12043));
  LUT3 #(.INIT(8'hE8)) lut_n12044 (.I0(n12039), .I1(n12042), .I2(n12043), .O(n12044));
  LUT3 #(.INIT(8'h96)) lut_n12045 (.I0(x3450), .I1(x3451), .I2(x3452), .O(n12045));
  LUT5 #(.INIT(32'h96696996)) lut_n12046 (.I0(x3441), .I1(x3442), .I2(x3443), .I3(n12040), .I4(n12041), .O(n12046));
  LUT5 #(.INIT(32'hFF969600)) lut_n12047 (.I0(x3447), .I1(x3448), .I2(x3449), .I3(n12045), .I4(n12046), .O(n12047));
  LUT3 #(.INIT(8'h96)) lut_n12048 (.I0(x3456), .I1(x3457), .I2(x3458), .O(n12048));
  LUT5 #(.INIT(32'h96696996)) lut_n12049 (.I0(x3447), .I1(x3448), .I2(x3449), .I3(n12045), .I4(n12046), .O(n12049));
  LUT5 #(.INIT(32'hFF969600)) lut_n12050 (.I0(x3453), .I1(x3454), .I2(x3455), .I3(n12048), .I4(n12049), .O(n12050));
  LUT3 #(.INIT(8'h96)) lut_n12051 (.I0(n12039), .I1(n12042), .I2(n12043), .O(n12051));
  LUT3 #(.INIT(8'hE8)) lut_n12052 (.I0(n12047), .I1(n12050), .I2(n12051), .O(n12052));
  LUT3 #(.INIT(8'h96)) lut_n12053 (.I0(n12024), .I1(n12032), .I2(n12033), .O(n12053));
  LUT3 #(.INIT(8'hE8)) lut_n12054 (.I0(n12044), .I1(n12052), .I2(n12053), .O(n12054));
  LUT3 #(.INIT(8'h96)) lut_n12055 (.I0(x3462), .I1(x3463), .I2(x3464), .O(n12055));
  LUT5 #(.INIT(32'h96696996)) lut_n12056 (.I0(x3453), .I1(x3454), .I2(x3455), .I3(n12048), .I4(n12049), .O(n12056));
  LUT5 #(.INIT(32'hFF969600)) lut_n12057 (.I0(x3459), .I1(x3460), .I2(x3461), .I3(n12055), .I4(n12056), .O(n12057));
  LUT3 #(.INIT(8'h96)) lut_n12058 (.I0(x3468), .I1(x3469), .I2(x3470), .O(n12058));
  LUT5 #(.INIT(32'h96696996)) lut_n12059 (.I0(x3459), .I1(x3460), .I2(x3461), .I3(n12055), .I4(n12056), .O(n12059));
  LUT5 #(.INIT(32'hFF969600)) lut_n12060 (.I0(x3465), .I1(x3466), .I2(x3467), .I3(n12058), .I4(n12059), .O(n12060));
  LUT3 #(.INIT(8'h96)) lut_n12061 (.I0(n12047), .I1(n12050), .I2(n12051), .O(n12061));
  LUT3 #(.INIT(8'hE8)) lut_n12062 (.I0(n12057), .I1(n12060), .I2(n12061), .O(n12062));
  LUT3 #(.INIT(8'h96)) lut_n12063 (.I0(x3474), .I1(x3475), .I2(x3476), .O(n12063));
  LUT5 #(.INIT(32'h96696996)) lut_n12064 (.I0(x3465), .I1(x3466), .I2(x3467), .I3(n12058), .I4(n12059), .O(n12064));
  LUT5 #(.INIT(32'hFF969600)) lut_n12065 (.I0(x3471), .I1(x3472), .I2(x3473), .I3(n12063), .I4(n12064), .O(n12065));
  LUT3 #(.INIT(8'h96)) lut_n12066 (.I0(x3480), .I1(x3481), .I2(x3482), .O(n12066));
  LUT5 #(.INIT(32'h96696996)) lut_n12067 (.I0(x3471), .I1(x3472), .I2(x3473), .I3(n12063), .I4(n12064), .O(n12067));
  LUT5 #(.INIT(32'hFF969600)) lut_n12068 (.I0(x3477), .I1(x3478), .I2(x3479), .I3(n12066), .I4(n12067), .O(n12068));
  LUT3 #(.INIT(8'h96)) lut_n12069 (.I0(n12057), .I1(n12060), .I2(n12061), .O(n12069));
  LUT3 #(.INIT(8'hE8)) lut_n12070 (.I0(n12065), .I1(n12068), .I2(n12069), .O(n12070));
  LUT3 #(.INIT(8'h96)) lut_n12071 (.I0(n12044), .I1(n12052), .I2(n12053), .O(n12071));
  LUT3 #(.INIT(8'hE8)) lut_n12072 (.I0(n12062), .I1(n12070), .I2(n12071), .O(n12072));
  LUT3 #(.INIT(8'h96)) lut_n12073 (.I0(n12016), .I1(n12034), .I2(n12035), .O(n12073));
  LUT3 #(.INIT(8'hE8)) lut_n12074 (.I0(n12054), .I1(n12072), .I2(n12073), .O(n12074));
  LUT3 #(.INIT(8'h96)) lut_n12075 (.I0(n11954), .I1(n11992), .I2(n11993), .O(n12075));
  LUT3 #(.INIT(8'hE8)) lut_n12076 (.I0(n12036), .I1(n12074), .I2(n12075), .O(n12076));
  LUT3 #(.INIT(8'h96)) lut_n12077 (.I0(x3486), .I1(x3487), .I2(x3488), .O(n12077));
  LUT5 #(.INIT(32'h96696996)) lut_n12078 (.I0(x3477), .I1(x3478), .I2(x3479), .I3(n12066), .I4(n12067), .O(n12078));
  LUT5 #(.INIT(32'hFF969600)) lut_n12079 (.I0(x3483), .I1(x3484), .I2(x3485), .I3(n12077), .I4(n12078), .O(n12079));
  LUT3 #(.INIT(8'h96)) lut_n12080 (.I0(x3492), .I1(x3493), .I2(x3494), .O(n12080));
  LUT5 #(.INIT(32'h96696996)) lut_n12081 (.I0(x3483), .I1(x3484), .I2(x3485), .I3(n12077), .I4(n12078), .O(n12081));
  LUT5 #(.INIT(32'hFF969600)) lut_n12082 (.I0(x3489), .I1(x3490), .I2(x3491), .I3(n12080), .I4(n12081), .O(n12082));
  LUT3 #(.INIT(8'h96)) lut_n12083 (.I0(n12065), .I1(n12068), .I2(n12069), .O(n12083));
  LUT3 #(.INIT(8'hE8)) lut_n12084 (.I0(n12079), .I1(n12082), .I2(n12083), .O(n12084));
  LUT3 #(.INIT(8'h96)) lut_n12085 (.I0(x3498), .I1(x3499), .I2(x3500), .O(n12085));
  LUT5 #(.INIT(32'h96696996)) lut_n12086 (.I0(x3489), .I1(x3490), .I2(x3491), .I3(n12080), .I4(n12081), .O(n12086));
  LUT5 #(.INIT(32'hFF969600)) lut_n12087 (.I0(x3495), .I1(x3496), .I2(x3497), .I3(n12085), .I4(n12086), .O(n12087));
  LUT3 #(.INIT(8'h96)) lut_n12088 (.I0(x3504), .I1(x3505), .I2(x3506), .O(n12088));
  LUT5 #(.INIT(32'h96696996)) lut_n12089 (.I0(x3495), .I1(x3496), .I2(x3497), .I3(n12085), .I4(n12086), .O(n12089));
  LUT5 #(.INIT(32'hFF969600)) lut_n12090 (.I0(x3501), .I1(x3502), .I2(x3503), .I3(n12088), .I4(n12089), .O(n12090));
  LUT3 #(.INIT(8'h96)) lut_n12091 (.I0(n12079), .I1(n12082), .I2(n12083), .O(n12091));
  LUT3 #(.INIT(8'hE8)) lut_n12092 (.I0(n12087), .I1(n12090), .I2(n12091), .O(n12092));
  LUT3 #(.INIT(8'h96)) lut_n12093 (.I0(n12062), .I1(n12070), .I2(n12071), .O(n12093));
  LUT3 #(.INIT(8'hE8)) lut_n12094 (.I0(n12084), .I1(n12092), .I2(n12093), .O(n12094));
  LUT3 #(.INIT(8'h96)) lut_n12095 (.I0(x3510), .I1(x3511), .I2(x3512), .O(n12095));
  LUT5 #(.INIT(32'h96696996)) lut_n12096 (.I0(x3501), .I1(x3502), .I2(x3503), .I3(n12088), .I4(n12089), .O(n12096));
  LUT5 #(.INIT(32'hFF969600)) lut_n12097 (.I0(x3507), .I1(x3508), .I2(x3509), .I3(n12095), .I4(n12096), .O(n12097));
  LUT3 #(.INIT(8'h96)) lut_n12098 (.I0(x3516), .I1(x3517), .I2(x3518), .O(n12098));
  LUT5 #(.INIT(32'h96696996)) lut_n12099 (.I0(x3507), .I1(x3508), .I2(x3509), .I3(n12095), .I4(n12096), .O(n12099));
  LUT5 #(.INIT(32'hFF969600)) lut_n12100 (.I0(x3513), .I1(x3514), .I2(x3515), .I3(n12098), .I4(n12099), .O(n12100));
  LUT3 #(.INIT(8'h96)) lut_n12101 (.I0(n12087), .I1(n12090), .I2(n12091), .O(n12101));
  LUT3 #(.INIT(8'hE8)) lut_n12102 (.I0(n12097), .I1(n12100), .I2(n12101), .O(n12102));
  LUT3 #(.INIT(8'h96)) lut_n12103 (.I0(x3522), .I1(x3523), .I2(x3524), .O(n12103));
  LUT5 #(.INIT(32'h96696996)) lut_n12104 (.I0(x3513), .I1(x3514), .I2(x3515), .I3(n12098), .I4(n12099), .O(n12104));
  LUT5 #(.INIT(32'hFF969600)) lut_n12105 (.I0(x3519), .I1(x3520), .I2(x3521), .I3(n12103), .I4(n12104), .O(n12105));
  LUT3 #(.INIT(8'h96)) lut_n12106 (.I0(x3528), .I1(x3529), .I2(x3530), .O(n12106));
  LUT5 #(.INIT(32'h96696996)) lut_n12107 (.I0(x3519), .I1(x3520), .I2(x3521), .I3(n12103), .I4(n12104), .O(n12107));
  LUT5 #(.INIT(32'hFF969600)) lut_n12108 (.I0(x3525), .I1(x3526), .I2(x3527), .I3(n12106), .I4(n12107), .O(n12108));
  LUT3 #(.INIT(8'h96)) lut_n12109 (.I0(n12097), .I1(n12100), .I2(n12101), .O(n12109));
  LUT3 #(.INIT(8'hE8)) lut_n12110 (.I0(n12105), .I1(n12108), .I2(n12109), .O(n12110));
  LUT3 #(.INIT(8'h96)) lut_n12111 (.I0(n12084), .I1(n12092), .I2(n12093), .O(n12111));
  LUT3 #(.INIT(8'hE8)) lut_n12112 (.I0(n12102), .I1(n12110), .I2(n12111), .O(n12112));
  LUT3 #(.INIT(8'h96)) lut_n12113 (.I0(n12054), .I1(n12072), .I2(n12073), .O(n12113));
  LUT3 #(.INIT(8'hE8)) lut_n12114 (.I0(n12094), .I1(n12112), .I2(n12113), .O(n12114));
  LUT3 #(.INIT(8'h96)) lut_n12115 (.I0(x3534), .I1(x3535), .I2(x3536), .O(n12115));
  LUT5 #(.INIT(32'h96696996)) lut_n12116 (.I0(x3525), .I1(x3526), .I2(x3527), .I3(n12106), .I4(n12107), .O(n12116));
  LUT5 #(.INIT(32'hFF969600)) lut_n12117 (.I0(x3531), .I1(x3532), .I2(x3533), .I3(n12115), .I4(n12116), .O(n12117));
  LUT3 #(.INIT(8'h96)) lut_n12118 (.I0(x3540), .I1(x3541), .I2(x3542), .O(n12118));
  LUT5 #(.INIT(32'h96696996)) lut_n12119 (.I0(x3531), .I1(x3532), .I2(x3533), .I3(n12115), .I4(n12116), .O(n12119));
  LUT5 #(.INIT(32'hFF969600)) lut_n12120 (.I0(x3537), .I1(x3538), .I2(x3539), .I3(n12118), .I4(n12119), .O(n12120));
  LUT3 #(.INIT(8'h96)) lut_n12121 (.I0(n12105), .I1(n12108), .I2(n12109), .O(n12121));
  LUT3 #(.INIT(8'hE8)) lut_n12122 (.I0(n12117), .I1(n12120), .I2(n12121), .O(n12122));
  LUT3 #(.INIT(8'h96)) lut_n12123 (.I0(x3546), .I1(x3547), .I2(x3548), .O(n12123));
  LUT5 #(.INIT(32'h96696996)) lut_n12124 (.I0(x3537), .I1(x3538), .I2(x3539), .I3(n12118), .I4(n12119), .O(n12124));
  LUT5 #(.INIT(32'hFF969600)) lut_n12125 (.I0(x3543), .I1(x3544), .I2(x3545), .I3(n12123), .I4(n12124), .O(n12125));
  LUT3 #(.INIT(8'h96)) lut_n12126 (.I0(x3552), .I1(x3553), .I2(x3554), .O(n12126));
  LUT5 #(.INIT(32'h96696996)) lut_n12127 (.I0(x3543), .I1(x3544), .I2(x3545), .I3(n12123), .I4(n12124), .O(n12127));
  LUT5 #(.INIT(32'hFF969600)) lut_n12128 (.I0(x3549), .I1(x3550), .I2(x3551), .I3(n12126), .I4(n12127), .O(n12128));
  LUT3 #(.INIT(8'h96)) lut_n12129 (.I0(n12117), .I1(n12120), .I2(n12121), .O(n12129));
  LUT3 #(.INIT(8'hE8)) lut_n12130 (.I0(n12125), .I1(n12128), .I2(n12129), .O(n12130));
  LUT3 #(.INIT(8'h96)) lut_n12131 (.I0(n12102), .I1(n12110), .I2(n12111), .O(n12131));
  LUT3 #(.INIT(8'hE8)) lut_n12132 (.I0(n12122), .I1(n12130), .I2(n12131), .O(n12132));
  LUT3 #(.INIT(8'h96)) lut_n12133 (.I0(x3558), .I1(x3559), .I2(x3560), .O(n12133));
  LUT5 #(.INIT(32'h96696996)) lut_n12134 (.I0(x3549), .I1(x3550), .I2(x3551), .I3(n12126), .I4(n12127), .O(n12134));
  LUT5 #(.INIT(32'hFF969600)) lut_n12135 (.I0(x3555), .I1(x3556), .I2(x3557), .I3(n12133), .I4(n12134), .O(n12135));
  LUT3 #(.INIT(8'h96)) lut_n12136 (.I0(x3564), .I1(x3565), .I2(x3566), .O(n12136));
  LUT5 #(.INIT(32'h96696996)) lut_n12137 (.I0(x3555), .I1(x3556), .I2(x3557), .I3(n12133), .I4(n12134), .O(n12137));
  LUT5 #(.INIT(32'hFF969600)) lut_n12138 (.I0(x3561), .I1(x3562), .I2(x3563), .I3(n12136), .I4(n12137), .O(n12138));
  LUT3 #(.INIT(8'h96)) lut_n12139 (.I0(n12125), .I1(n12128), .I2(n12129), .O(n12139));
  LUT3 #(.INIT(8'hE8)) lut_n12140 (.I0(n12135), .I1(n12138), .I2(n12139), .O(n12140));
  LUT3 #(.INIT(8'h96)) lut_n12141 (.I0(x3570), .I1(x3571), .I2(x3572), .O(n12141));
  LUT5 #(.INIT(32'h96696996)) lut_n12142 (.I0(x3561), .I1(x3562), .I2(x3563), .I3(n12136), .I4(n12137), .O(n12142));
  LUT5 #(.INIT(32'hFF969600)) lut_n12143 (.I0(x3567), .I1(x3568), .I2(x3569), .I3(n12141), .I4(n12142), .O(n12143));
  LUT3 #(.INIT(8'h96)) lut_n12144 (.I0(x3576), .I1(x3577), .I2(x3578), .O(n12144));
  LUT5 #(.INIT(32'h96696996)) lut_n12145 (.I0(x3567), .I1(x3568), .I2(x3569), .I3(n12141), .I4(n12142), .O(n12145));
  LUT5 #(.INIT(32'hFF969600)) lut_n12146 (.I0(x3573), .I1(x3574), .I2(x3575), .I3(n12144), .I4(n12145), .O(n12146));
  LUT3 #(.INIT(8'h96)) lut_n12147 (.I0(n12135), .I1(n12138), .I2(n12139), .O(n12147));
  LUT3 #(.INIT(8'hE8)) lut_n12148 (.I0(n12143), .I1(n12146), .I2(n12147), .O(n12148));
  LUT3 #(.INIT(8'h96)) lut_n12149 (.I0(n12122), .I1(n12130), .I2(n12131), .O(n12149));
  LUT3 #(.INIT(8'hE8)) lut_n12150 (.I0(n12140), .I1(n12148), .I2(n12149), .O(n12150));
  LUT3 #(.INIT(8'h96)) lut_n12151 (.I0(n12094), .I1(n12112), .I2(n12113), .O(n12151));
  LUT3 #(.INIT(8'hE8)) lut_n12152 (.I0(n12132), .I1(n12150), .I2(n12151), .O(n12152));
  LUT3 #(.INIT(8'h96)) lut_n12153 (.I0(n12036), .I1(n12074), .I2(n12075), .O(n12153));
  LUT3 #(.INIT(8'hE8)) lut_n12154 (.I0(n12114), .I1(n12152), .I2(n12153), .O(n12154));
  LUT3 #(.INIT(8'h96)) lut_n12155 (.I0(n11916), .I1(n11994), .I2(n11995), .O(n12155));
  LUT3 #(.INIT(8'hE8)) lut_n12156 (.I0(n12076), .I1(n12154), .I2(n12155), .O(n12156));
  LUT3 #(.INIT(8'h96)) lut_n12157 (.I0(x3582), .I1(x3583), .I2(x3584), .O(n12157));
  LUT5 #(.INIT(32'h96696996)) lut_n12158 (.I0(x3573), .I1(x3574), .I2(x3575), .I3(n12144), .I4(n12145), .O(n12158));
  LUT5 #(.INIT(32'hFF969600)) lut_n12159 (.I0(x3579), .I1(x3580), .I2(x3581), .I3(n12157), .I4(n12158), .O(n12159));
  LUT3 #(.INIT(8'h96)) lut_n12160 (.I0(x3588), .I1(x3589), .I2(x3590), .O(n12160));
  LUT5 #(.INIT(32'h96696996)) lut_n12161 (.I0(x3579), .I1(x3580), .I2(x3581), .I3(n12157), .I4(n12158), .O(n12161));
  LUT5 #(.INIT(32'hFF969600)) lut_n12162 (.I0(x3585), .I1(x3586), .I2(x3587), .I3(n12160), .I4(n12161), .O(n12162));
  LUT3 #(.INIT(8'h96)) lut_n12163 (.I0(n12143), .I1(n12146), .I2(n12147), .O(n12163));
  LUT3 #(.INIT(8'hE8)) lut_n12164 (.I0(n12159), .I1(n12162), .I2(n12163), .O(n12164));
  LUT3 #(.INIT(8'h96)) lut_n12165 (.I0(x3594), .I1(x3595), .I2(x3596), .O(n12165));
  LUT5 #(.INIT(32'h96696996)) lut_n12166 (.I0(x3585), .I1(x3586), .I2(x3587), .I3(n12160), .I4(n12161), .O(n12166));
  LUT5 #(.INIT(32'hFF969600)) lut_n12167 (.I0(x3591), .I1(x3592), .I2(x3593), .I3(n12165), .I4(n12166), .O(n12167));
  LUT3 #(.INIT(8'h96)) lut_n12168 (.I0(x3600), .I1(x3601), .I2(x3602), .O(n12168));
  LUT5 #(.INIT(32'h96696996)) lut_n12169 (.I0(x3591), .I1(x3592), .I2(x3593), .I3(n12165), .I4(n12166), .O(n12169));
  LUT5 #(.INIT(32'hFF969600)) lut_n12170 (.I0(x3597), .I1(x3598), .I2(x3599), .I3(n12168), .I4(n12169), .O(n12170));
  LUT3 #(.INIT(8'h96)) lut_n12171 (.I0(n12159), .I1(n12162), .I2(n12163), .O(n12171));
  LUT3 #(.INIT(8'hE8)) lut_n12172 (.I0(n12167), .I1(n12170), .I2(n12171), .O(n12172));
  LUT3 #(.INIT(8'h96)) lut_n12173 (.I0(n12140), .I1(n12148), .I2(n12149), .O(n12173));
  LUT3 #(.INIT(8'hE8)) lut_n12174 (.I0(n12164), .I1(n12172), .I2(n12173), .O(n12174));
  LUT3 #(.INIT(8'h96)) lut_n12175 (.I0(x3606), .I1(x3607), .I2(x3608), .O(n12175));
  LUT5 #(.INIT(32'h96696996)) lut_n12176 (.I0(x3597), .I1(x3598), .I2(x3599), .I3(n12168), .I4(n12169), .O(n12176));
  LUT5 #(.INIT(32'hFF969600)) lut_n12177 (.I0(x3603), .I1(x3604), .I2(x3605), .I3(n12175), .I4(n12176), .O(n12177));
  LUT3 #(.INIT(8'h96)) lut_n12178 (.I0(x3612), .I1(x3613), .I2(x3614), .O(n12178));
  LUT5 #(.INIT(32'h96696996)) lut_n12179 (.I0(x3603), .I1(x3604), .I2(x3605), .I3(n12175), .I4(n12176), .O(n12179));
  LUT5 #(.INIT(32'hFF969600)) lut_n12180 (.I0(x3609), .I1(x3610), .I2(x3611), .I3(n12178), .I4(n12179), .O(n12180));
  LUT3 #(.INIT(8'h96)) lut_n12181 (.I0(n12167), .I1(n12170), .I2(n12171), .O(n12181));
  LUT3 #(.INIT(8'hE8)) lut_n12182 (.I0(n12177), .I1(n12180), .I2(n12181), .O(n12182));
  LUT3 #(.INIT(8'h96)) lut_n12183 (.I0(x3618), .I1(x3619), .I2(x3620), .O(n12183));
  LUT5 #(.INIT(32'h96696996)) lut_n12184 (.I0(x3609), .I1(x3610), .I2(x3611), .I3(n12178), .I4(n12179), .O(n12184));
  LUT5 #(.INIT(32'hFF969600)) lut_n12185 (.I0(x3615), .I1(x3616), .I2(x3617), .I3(n12183), .I4(n12184), .O(n12185));
  LUT3 #(.INIT(8'h96)) lut_n12186 (.I0(x3624), .I1(x3625), .I2(x3626), .O(n12186));
  LUT5 #(.INIT(32'h96696996)) lut_n12187 (.I0(x3615), .I1(x3616), .I2(x3617), .I3(n12183), .I4(n12184), .O(n12187));
  LUT5 #(.INIT(32'hFF969600)) lut_n12188 (.I0(x3621), .I1(x3622), .I2(x3623), .I3(n12186), .I4(n12187), .O(n12188));
  LUT3 #(.INIT(8'h96)) lut_n12189 (.I0(n12177), .I1(n12180), .I2(n12181), .O(n12189));
  LUT3 #(.INIT(8'hE8)) lut_n12190 (.I0(n12185), .I1(n12188), .I2(n12189), .O(n12190));
  LUT3 #(.INIT(8'h96)) lut_n12191 (.I0(n12164), .I1(n12172), .I2(n12173), .O(n12191));
  LUT3 #(.INIT(8'hE8)) lut_n12192 (.I0(n12182), .I1(n12190), .I2(n12191), .O(n12192));
  LUT3 #(.INIT(8'h96)) lut_n12193 (.I0(n12132), .I1(n12150), .I2(n12151), .O(n12193));
  LUT3 #(.INIT(8'hE8)) lut_n12194 (.I0(n12174), .I1(n12192), .I2(n12193), .O(n12194));
  LUT3 #(.INIT(8'h96)) lut_n12195 (.I0(x3630), .I1(x3631), .I2(x3632), .O(n12195));
  LUT5 #(.INIT(32'h96696996)) lut_n12196 (.I0(x3621), .I1(x3622), .I2(x3623), .I3(n12186), .I4(n12187), .O(n12196));
  LUT5 #(.INIT(32'hFF969600)) lut_n12197 (.I0(x3627), .I1(x3628), .I2(x3629), .I3(n12195), .I4(n12196), .O(n12197));
  LUT3 #(.INIT(8'h96)) lut_n12198 (.I0(x3636), .I1(x3637), .I2(x3638), .O(n12198));
  LUT5 #(.INIT(32'h96696996)) lut_n12199 (.I0(x3627), .I1(x3628), .I2(x3629), .I3(n12195), .I4(n12196), .O(n12199));
  LUT5 #(.INIT(32'hFF969600)) lut_n12200 (.I0(x3633), .I1(x3634), .I2(x3635), .I3(n12198), .I4(n12199), .O(n12200));
  LUT3 #(.INIT(8'h96)) lut_n12201 (.I0(n12185), .I1(n12188), .I2(n12189), .O(n12201));
  LUT3 #(.INIT(8'hE8)) lut_n12202 (.I0(n12197), .I1(n12200), .I2(n12201), .O(n12202));
  LUT3 #(.INIT(8'h96)) lut_n12203 (.I0(x3642), .I1(x3643), .I2(x3644), .O(n12203));
  LUT5 #(.INIT(32'h96696996)) lut_n12204 (.I0(x3633), .I1(x3634), .I2(x3635), .I3(n12198), .I4(n12199), .O(n12204));
  LUT5 #(.INIT(32'hFF969600)) lut_n12205 (.I0(x3639), .I1(x3640), .I2(x3641), .I3(n12203), .I4(n12204), .O(n12205));
  LUT3 #(.INIT(8'h96)) lut_n12206 (.I0(x3648), .I1(x3649), .I2(x3650), .O(n12206));
  LUT5 #(.INIT(32'h96696996)) lut_n12207 (.I0(x3639), .I1(x3640), .I2(x3641), .I3(n12203), .I4(n12204), .O(n12207));
  LUT5 #(.INIT(32'hFF969600)) lut_n12208 (.I0(x3645), .I1(x3646), .I2(x3647), .I3(n12206), .I4(n12207), .O(n12208));
  LUT3 #(.INIT(8'h96)) lut_n12209 (.I0(n12197), .I1(n12200), .I2(n12201), .O(n12209));
  LUT3 #(.INIT(8'hE8)) lut_n12210 (.I0(n12205), .I1(n12208), .I2(n12209), .O(n12210));
  LUT3 #(.INIT(8'h96)) lut_n12211 (.I0(n12182), .I1(n12190), .I2(n12191), .O(n12211));
  LUT3 #(.INIT(8'hE8)) lut_n12212 (.I0(n12202), .I1(n12210), .I2(n12211), .O(n12212));
  LUT3 #(.INIT(8'h96)) lut_n12213 (.I0(x3654), .I1(x3655), .I2(x3656), .O(n12213));
  LUT5 #(.INIT(32'h96696996)) lut_n12214 (.I0(x3645), .I1(x3646), .I2(x3647), .I3(n12206), .I4(n12207), .O(n12214));
  LUT5 #(.INIT(32'hFF969600)) lut_n12215 (.I0(x3651), .I1(x3652), .I2(x3653), .I3(n12213), .I4(n12214), .O(n12215));
  LUT3 #(.INIT(8'h96)) lut_n12216 (.I0(x3660), .I1(x3661), .I2(x3662), .O(n12216));
  LUT5 #(.INIT(32'h96696996)) lut_n12217 (.I0(x3651), .I1(x3652), .I2(x3653), .I3(n12213), .I4(n12214), .O(n12217));
  LUT5 #(.INIT(32'hFF969600)) lut_n12218 (.I0(x3657), .I1(x3658), .I2(x3659), .I3(n12216), .I4(n12217), .O(n12218));
  LUT3 #(.INIT(8'h96)) lut_n12219 (.I0(n12205), .I1(n12208), .I2(n12209), .O(n12219));
  LUT3 #(.INIT(8'hE8)) lut_n12220 (.I0(n12215), .I1(n12218), .I2(n12219), .O(n12220));
  LUT3 #(.INIT(8'h96)) lut_n12221 (.I0(x3666), .I1(x3667), .I2(x3668), .O(n12221));
  LUT5 #(.INIT(32'h96696996)) lut_n12222 (.I0(x3657), .I1(x3658), .I2(x3659), .I3(n12216), .I4(n12217), .O(n12222));
  LUT5 #(.INIT(32'hFF969600)) lut_n12223 (.I0(x3663), .I1(x3664), .I2(x3665), .I3(n12221), .I4(n12222), .O(n12223));
  LUT3 #(.INIT(8'h96)) lut_n12224 (.I0(x3672), .I1(x3673), .I2(x3674), .O(n12224));
  LUT5 #(.INIT(32'h96696996)) lut_n12225 (.I0(x3663), .I1(x3664), .I2(x3665), .I3(n12221), .I4(n12222), .O(n12225));
  LUT5 #(.INIT(32'hFF969600)) lut_n12226 (.I0(x3669), .I1(x3670), .I2(x3671), .I3(n12224), .I4(n12225), .O(n12226));
  LUT3 #(.INIT(8'h96)) lut_n12227 (.I0(n12215), .I1(n12218), .I2(n12219), .O(n12227));
  LUT3 #(.INIT(8'hE8)) lut_n12228 (.I0(n12223), .I1(n12226), .I2(n12227), .O(n12228));
  LUT3 #(.INIT(8'h96)) lut_n12229 (.I0(n12202), .I1(n12210), .I2(n12211), .O(n12229));
  LUT3 #(.INIT(8'hE8)) lut_n12230 (.I0(n12220), .I1(n12228), .I2(n12229), .O(n12230));
  LUT3 #(.INIT(8'h96)) lut_n12231 (.I0(n12174), .I1(n12192), .I2(n12193), .O(n12231));
  LUT3 #(.INIT(8'hE8)) lut_n12232 (.I0(n12212), .I1(n12230), .I2(n12231), .O(n12232));
  LUT3 #(.INIT(8'h96)) lut_n12233 (.I0(n12114), .I1(n12152), .I2(n12153), .O(n12233));
  LUT3 #(.INIT(8'hE8)) lut_n12234 (.I0(n12194), .I1(n12232), .I2(n12233), .O(n12234));
  LUT3 #(.INIT(8'h96)) lut_n12235 (.I0(x3678), .I1(x3679), .I2(x3680), .O(n12235));
  LUT5 #(.INIT(32'h96696996)) lut_n12236 (.I0(x3669), .I1(x3670), .I2(x3671), .I3(n12224), .I4(n12225), .O(n12236));
  LUT5 #(.INIT(32'hFF969600)) lut_n12237 (.I0(x3675), .I1(x3676), .I2(x3677), .I3(n12235), .I4(n12236), .O(n12237));
  LUT3 #(.INIT(8'h96)) lut_n12238 (.I0(x3684), .I1(x3685), .I2(x3686), .O(n12238));
  LUT5 #(.INIT(32'h96696996)) lut_n12239 (.I0(x3675), .I1(x3676), .I2(x3677), .I3(n12235), .I4(n12236), .O(n12239));
  LUT5 #(.INIT(32'hFF969600)) lut_n12240 (.I0(x3681), .I1(x3682), .I2(x3683), .I3(n12238), .I4(n12239), .O(n12240));
  LUT3 #(.INIT(8'h96)) lut_n12241 (.I0(n12223), .I1(n12226), .I2(n12227), .O(n12241));
  LUT3 #(.INIT(8'hE8)) lut_n12242 (.I0(n12237), .I1(n12240), .I2(n12241), .O(n12242));
  LUT3 #(.INIT(8'h96)) lut_n12243 (.I0(x3690), .I1(x3691), .I2(x3692), .O(n12243));
  LUT5 #(.INIT(32'h96696996)) lut_n12244 (.I0(x3681), .I1(x3682), .I2(x3683), .I3(n12238), .I4(n12239), .O(n12244));
  LUT5 #(.INIT(32'hFF969600)) lut_n12245 (.I0(x3687), .I1(x3688), .I2(x3689), .I3(n12243), .I4(n12244), .O(n12245));
  LUT3 #(.INIT(8'h96)) lut_n12246 (.I0(x3696), .I1(x3697), .I2(x3698), .O(n12246));
  LUT5 #(.INIT(32'h96696996)) lut_n12247 (.I0(x3687), .I1(x3688), .I2(x3689), .I3(n12243), .I4(n12244), .O(n12247));
  LUT5 #(.INIT(32'hFF969600)) lut_n12248 (.I0(x3693), .I1(x3694), .I2(x3695), .I3(n12246), .I4(n12247), .O(n12248));
  LUT3 #(.INIT(8'h96)) lut_n12249 (.I0(n12237), .I1(n12240), .I2(n12241), .O(n12249));
  LUT3 #(.INIT(8'hE8)) lut_n12250 (.I0(n12245), .I1(n12248), .I2(n12249), .O(n12250));
  LUT3 #(.INIT(8'h96)) lut_n12251 (.I0(n12220), .I1(n12228), .I2(n12229), .O(n12251));
  LUT3 #(.INIT(8'hE8)) lut_n12252 (.I0(n12242), .I1(n12250), .I2(n12251), .O(n12252));
  LUT3 #(.INIT(8'h96)) lut_n12253 (.I0(x3702), .I1(x3703), .I2(x3704), .O(n12253));
  LUT5 #(.INIT(32'h96696996)) lut_n12254 (.I0(x3693), .I1(x3694), .I2(x3695), .I3(n12246), .I4(n12247), .O(n12254));
  LUT5 #(.INIT(32'hFF969600)) lut_n12255 (.I0(x3699), .I1(x3700), .I2(x3701), .I3(n12253), .I4(n12254), .O(n12255));
  LUT3 #(.INIT(8'h96)) lut_n12256 (.I0(x3708), .I1(x3709), .I2(x3710), .O(n12256));
  LUT5 #(.INIT(32'h96696996)) lut_n12257 (.I0(x3699), .I1(x3700), .I2(x3701), .I3(n12253), .I4(n12254), .O(n12257));
  LUT5 #(.INIT(32'hFF969600)) lut_n12258 (.I0(x3705), .I1(x3706), .I2(x3707), .I3(n12256), .I4(n12257), .O(n12258));
  LUT3 #(.INIT(8'h96)) lut_n12259 (.I0(n12245), .I1(n12248), .I2(n12249), .O(n12259));
  LUT3 #(.INIT(8'hE8)) lut_n12260 (.I0(n12255), .I1(n12258), .I2(n12259), .O(n12260));
  LUT3 #(.INIT(8'h96)) lut_n12261 (.I0(x3714), .I1(x3715), .I2(x3716), .O(n12261));
  LUT5 #(.INIT(32'h96696996)) lut_n12262 (.I0(x3705), .I1(x3706), .I2(x3707), .I3(n12256), .I4(n12257), .O(n12262));
  LUT5 #(.INIT(32'hFF969600)) lut_n12263 (.I0(x3711), .I1(x3712), .I2(x3713), .I3(n12261), .I4(n12262), .O(n12263));
  LUT3 #(.INIT(8'h96)) lut_n12264 (.I0(x3720), .I1(x3721), .I2(x3722), .O(n12264));
  LUT5 #(.INIT(32'h96696996)) lut_n12265 (.I0(x3711), .I1(x3712), .I2(x3713), .I3(n12261), .I4(n12262), .O(n12265));
  LUT5 #(.INIT(32'hFF969600)) lut_n12266 (.I0(x3717), .I1(x3718), .I2(x3719), .I3(n12264), .I4(n12265), .O(n12266));
  LUT3 #(.INIT(8'h96)) lut_n12267 (.I0(n12255), .I1(n12258), .I2(n12259), .O(n12267));
  LUT3 #(.INIT(8'hE8)) lut_n12268 (.I0(n12263), .I1(n12266), .I2(n12267), .O(n12268));
  LUT3 #(.INIT(8'h96)) lut_n12269 (.I0(n12242), .I1(n12250), .I2(n12251), .O(n12269));
  LUT3 #(.INIT(8'hE8)) lut_n12270 (.I0(n12260), .I1(n12268), .I2(n12269), .O(n12270));
  LUT3 #(.INIT(8'h96)) lut_n12271 (.I0(n12212), .I1(n12230), .I2(n12231), .O(n12271));
  LUT3 #(.INIT(8'hE8)) lut_n12272 (.I0(n12252), .I1(n12270), .I2(n12271), .O(n12272));
  LUT3 #(.INIT(8'h96)) lut_n12273 (.I0(x3726), .I1(x3727), .I2(x3728), .O(n12273));
  LUT5 #(.INIT(32'h96696996)) lut_n12274 (.I0(x3717), .I1(x3718), .I2(x3719), .I3(n12264), .I4(n12265), .O(n12274));
  LUT5 #(.INIT(32'hFF969600)) lut_n12275 (.I0(x3723), .I1(x3724), .I2(x3725), .I3(n12273), .I4(n12274), .O(n12275));
  LUT3 #(.INIT(8'h96)) lut_n12276 (.I0(x3732), .I1(x3733), .I2(x3734), .O(n12276));
  LUT5 #(.INIT(32'h96696996)) lut_n12277 (.I0(x3723), .I1(x3724), .I2(x3725), .I3(n12273), .I4(n12274), .O(n12277));
  LUT5 #(.INIT(32'hFF969600)) lut_n12278 (.I0(x3729), .I1(x3730), .I2(x3731), .I3(n12276), .I4(n12277), .O(n12278));
  LUT3 #(.INIT(8'h96)) lut_n12279 (.I0(n12263), .I1(n12266), .I2(n12267), .O(n12279));
  LUT3 #(.INIT(8'hE8)) lut_n12280 (.I0(n12275), .I1(n12278), .I2(n12279), .O(n12280));
  LUT3 #(.INIT(8'h96)) lut_n12281 (.I0(x3738), .I1(x3739), .I2(x3740), .O(n12281));
  LUT5 #(.INIT(32'h96696996)) lut_n12282 (.I0(x3729), .I1(x3730), .I2(x3731), .I3(n12276), .I4(n12277), .O(n12282));
  LUT5 #(.INIT(32'hFF969600)) lut_n12283 (.I0(x3735), .I1(x3736), .I2(x3737), .I3(n12281), .I4(n12282), .O(n12283));
  LUT3 #(.INIT(8'h96)) lut_n12284 (.I0(x3744), .I1(x3745), .I2(x3746), .O(n12284));
  LUT5 #(.INIT(32'h96696996)) lut_n12285 (.I0(x3735), .I1(x3736), .I2(x3737), .I3(n12281), .I4(n12282), .O(n12285));
  LUT5 #(.INIT(32'hFF969600)) lut_n12286 (.I0(x3741), .I1(x3742), .I2(x3743), .I3(n12284), .I4(n12285), .O(n12286));
  LUT3 #(.INIT(8'h96)) lut_n12287 (.I0(n12275), .I1(n12278), .I2(n12279), .O(n12287));
  LUT3 #(.INIT(8'hE8)) lut_n12288 (.I0(n12283), .I1(n12286), .I2(n12287), .O(n12288));
  LUT3 #(.INIT(8'h96)) lut_n12289 (.I0(n12260), .I1(n12268), .I2(n12269), .O(n12289));
  LUT3 #(.INIT(8'hE8)) lut_n12290 (.I0(n12280), .I1(n12288), .I2(n12289), .O(n12290));
  LUT3 #(.INIT(8'h96)) lut_n12291 (.I0(x3750), .I1(x3751), .I2(x3752), .O(n12291));
  LUT5 #(.INIT(32'h96696996)) lut_n12292 (.I0(x3741), .I1(x3742), .I2(x3743), .I3(n12284), .I4(n12285), .O(n12292));
  LUT5 #(.INIT(32'hFF969600)) lut_n12293 (.I0(x3747), .I1(x3748), .I2(x3749), .I3(n12291), .I4(n12292), .O(n12293));
  LUT3 #(.INIT(8'h96)) lut_n12294 (.I0(x3756), .I1(x3757), .I2(x3758), .O(n12294));
  LUT5 #(.INIT(32'h96696996)) lut_n12295 (.I0(x3747), .I1(x3748), .I2(x3749), .I3(n12291), .I4(n12292), .O(n12295));
  LUT5 #(.INIT(32'hFF969600)) lut_n12296 (.I0(x3753), .I1(x3754), .I2(x3755), .I3(n12294), .I4(n12295), .O(n12296));
  LUT3 #(.INIT(8'h96)) lut_n12297 (.I0(n12283), .I1(n12286), .I2(n12287), .O(n12297));
  LUT3 #(.INIT(8'hE8)) lut_n12298 (.I0(n12293), .I1(n12296), .I2(n12297), .O(n12298));
  LUT3 #(.INIT(8'h96)) lut_n12299 (.I0(x3762), .I1(x3763), .I2(x3764), .O(n12299));
  LUT5 #(.INIT(32'h96696996)) lut_n12300 (.I0(x3753), .I1(x3754), .I2(x3755), .I3(n12294), .I4(n12295), .O(n12300));
  LUT5 #(.INIT(32'hFF969600)) lut_n12301 (.I0(x3759), .I1(x3760), .I2(x3761), .I3(n12299), .I4(n12300), .O(n12301));
  LUT3 #(.INIT(8'h96)) lut_n12302 (.I0(x3768), .I1(x3769), .I2(x3770), .O(n12302));
  LUT5 #(.INIT(32'h96696996)) lut_n12303 (.I0(x3759), .I1(x3760), .I2(x3761), .I3(n12299), .I4(n12300), .O(n12303));
  LUT5 #(.INIT(32'hFF969600)) lut_n12304 (.I0(x3765), .I1(x3766), .I2(x3767), .I3(n12302), .I4(n12303), .O(n12304));
  LUT3 #(.INIT(8'h96)) lut_n12305 (.I0(n12293), .I1(n12296), .I2(n12297), .O(n12305));
  LUT3 #(.INIT(8'hE8)) lut_n12306 (.I0(n12301), .I1(n12304), .I2(n12305), .O(n12306));
  LUT3 #(.INIT(8'h96)) lut_n12307 (.I0(n12280), .I1(n12288), .I2(n12289), .O(n12307));
  LUT3 #(.INIT(8'hE8)) lut_n12308 (.I0(n12298), .I1(n12306), .I2(n12307), .O(n12308));
  LUT3 #(.INIT(8'h96)) lut_n12309 (.I0(n12252), .I1(n12270), .I2(n12271), .O(n12309));
  LUT3 #(.INIT(8'hE8)) lut_n12310 (.I0(n12290), .I1(n12308), .I2(n12309), .O(n12310));
  LUT3 #(.INIT(8'h96)) lut_n12311 (.I0(n12194), .I1(n12232), .I2(n12233), .O(n12311));
  LUT3 #(.INIT(8'hE8)) lut_n12312 (.I0(n12272), .I1(n12310), .I2(n12311), .O(n12312));
  LUT3 #(.INIT(8'h96)) lut_n12313 (.I0(n12076), .I1(n12154), .I2(n12155), .O(n12313));
  LUT3 #(.INIT(8'hE8)) lut_n12314 (.I0(n12234), .I1(n12312), .I2(n12313), .O(n12314));
  LUT3 #(.INIT(8'h96)) lut_n12315 (.I0(n11838), .I1(n11996), .I2(n11997), .O(n12315));
  LUT3 #(.INIT(8'hE8)) lut_n12316 (.I0(n12156), .I1(n12314), .I2(n12315), .O(n12316));
  LUT3 #(.INIT(8'h96)) lut_n12317 (.I0(n11360), .I1(n11678), .I2(n11679), .O(n12317));
  LUT3 #(.INIT(8'hE8)) lut_n12318 (.I0(n11998), .I1(n12316), .I2(n12317), .O(n12318));
  LUT3 #(.INIT(8'h96)) lut_n12319 (.I0(n10399), .I1(n11037), .I2(n11038), .O(n12319));
  LUT3 #(.INIT(8'hE8)) lut_n12320 (.I0(n11680), .I1(n12318), .I2(n12319), .O(n12320));
  LUT3 #(.INIT(8'h96)) lut_n12321 (.I0(x3774), .I1(x3775), .I2(x3776), .O(n12321));
  LUT5 #(.INIT(32'h96696996)) lut_n12322 (.I0(x3765), .I1(x3766), .I2(x3767), .I3(n12302), .I4(n12303), .O(n12322));
  LUT5 #(.INIT(32'hFF969600)) lut_n12323 (.I0(x3771), .I1(x3772), .I2(x3773), .I3(n12321), .I4(n12322), .O(n12323));
  LUT3 #(.INIT(8'h96)) lut_n12324 (.I0(x3780), .I1(x3781), .I2(x3782), .O(n12324));
  LUT5 #(.INIT(32'h96696996)) lut_n12325 (.I0(x3771), .I1(x3772), .I2(x3773), .I3(n12321), .I4(n12322), .O(n12325));
  LUT5 #(.INIT(32'hFF969600)) lut_n12326 (.I0(x3777), .I1(x3778), .I2(x3779), .I3(n12324), .I4(n12325), .O(n12326));
  LUT3 #(.INIT(8'h96)) lut_n12327 (.I0(n12301), .I1(n12304), .I2(n12305), .O(n12327));
  LUT3 #(.INIT(8'hE8)) lut_n12328 (.I0(n12323), .I1(n12326), .I2(n12327), .O(n12328));
  LUT3 #(.INIT(8'h96)) lut_n12329 (.I0(x3786), .I1(x3787), .I2(x3788), .O(n12329));
  LUT5 #(.INIT(32'h96696996)) lut_n12330 (.I0(x3777), .I1(x3778), .I2(x3779), .I3(n12324), .I4(n12325), .O(n12330));
  LUT5 #(.INIT(32'hFF969600)) lut_n12331 (.I0(x3783), .I1(x3784), .I2(x3785), .I3(n12329), .I4(n12330), .O(n12331));
  LUT3 #(.INIT(8'h96)) lut_n12332 (.I0(x3792), .I1(x3793), .I2(x3794), .O(n12332));
  LUT5 #(.INIT(32'h96696996)) lut_n12333 (.I0(x3783), .I1(x3784), .I2(x3785), .I3(n12329), .I4(n12330), .O(n12333));
  LUT5 #(.INIT(32'hFF969600)) lut_n12334 (.I0(x3789), .I1(x3790), .I2(x3791), .I3(n12332), .I4(n12333), .O(n12334));
  LUT3 #(.INIT(8'h96)) lut_n12335 (.I0(n12323), .I1(n12326), .I2(n12327), .O(n12335));
  LUT3 #(.INIT(8'hE8)) lut_n12336 (.I0(n12331), .I1(n12334), .I2(n12335), .O(n12336));
  LUT3 #(.INIT(8'h96)) lut_n12337 (.I0(n12298), .I1(n12306), .I2(n12307), .O(n12337));
  LUT3 #(.INIT(8'hE8)) lut_n12338 (.I0(n12328), .I1(n12336), .I2(n12337), .O(n12338));
  LUT3 #(.INIT(8'h96)) lut_n12339 (.I0(x3798), .I1(x3799), .I2(x3800), .O(n12339));
  LUT5 #(.INIT(32'h96696996)) lut_n12340 (.I0(x3789), .I1(x3790), .I2(x3791), .I3(n12332), .I4(n12333), .O(n12340));
  LUT5 #(.INIT(32'hFF969600)) lut_n12341 (.I0(x3795), .I1(x3796), .I2(x3797), .I3(n12339), .I4(n12340), .O(n12341));
  LUT3 #(.INIT(8'h96)) lut_n12342 (.I0(x3804), .I1(x3805), .I2(x3806), .O(n12342));
  LUT5 #(.INIT(32'h96696996)) lut_n12343 (.I0(x3795), .I1(x3796), .I2(x3797), .I3(n12339), .I4(n12340), .O(n12343));
  LUT5 #(.INIT(32'hFF969600)) lut_n12344 (.I0(x3801), .I1(x3802), .I2(x3803), .I3(n12342), .I4(n12343), .O(n12344));
  LUT3 #(.INIT(8'h96)) lut_n12345 (.I0(n12331), .I1(n12334), .I2(n12335), .O(n12345));
  LUT3 #(.INIT(8'hE8)) lut_n12346 (.I0(n12341), .I1(n12344), .I2(n12345), .O(n12346));
  LUT3 #(.INIT(8'h96)) lut_n12347 (.I0(x3810), .I1(x3811), .I2(x3812), .O(n12347));
  LUT5 #(.INIT(32'h96696996)) lut_n12348 (.I0(x3801), .I1(x3802), .I2(x3803), .I3(n12342), .I4(n12343), .O(n12348));
  LUT5 #(.INIT(32'hFF969600)) lut_n12349 (.I0(x3807), .I1(x3808), .I2(x3809), .I3(n12347), .I4(n12348), .O(n12349));
  LUT3 #(.INIT(8'h96)) lut_n12350 (.I0(x3816), .I1(x3817), .I2(x3818), .O(n12350));
  LUT5 #(.INIT(32'h96696996)) lut_n12351 (.I0(x3807), .I1(x3808), .I2(x3809), .I3(n12347), .I4(n12348), .O(n12351));
  LUT5 #(.INIT(32'hFF969600)) lut_n12352 (.I0(x3813), .I1(x3814), .I2(x3815), .I3(n12350), .I4(n12351), .O(n12352));
  LUT3 #(.INIT(8'h96)) lut_n12353 (.I0(n12341), .I1(n12344), .I2(n12345), .O(n12353));
  LUT3 #(.INIT(8'hE8)) lut_n12354 (.I0(n12349), .I1(n12352), .I2(n12353), .O(n12354));
  LUT3 #(.INIT(8'h96)) lut_n12355 (.I0(n12328), .I1(n12336), .I2(n12337), .O(n12355));
  LUT3 #(.INIT(8'hE8)) lut_n12356 (.I0(n12346), .I1(n12354), .I2(n12355), .O(n12356));
  LUT3 #(.INIT(8'h96)) lut_n12357 (.I0(n12290), .I1(n12308), .I2(n12309), .O(n12357));
  LUT3 #(.INIT(8'hE8)) lut_n12358 (.I0(n12338), .I1(n12356), .I2(n12357), .O(n12358));
  LUT3 #(.INIT(8'h96)) lut_n12359 (.I0(x3822), .I1(x3823), .I2(x3824), .O(n12359));
  LUT5 #(.INIT(32'h96696996)) lut_n12360 (.I0(x3813), .I1(x3814), .I2(x3815), .I3(n12350), .I4(n12351), .O(n12360));
  LUT5 #(.INIT(32'hFF969600)) lut_n12361 (.I0(x3819), .I1(x3820), .I2(x3821), .I3(n12359), .I4(n12360), .O(n12361));
  LUT3 #(.INIT(8'h96)) lut_n12362 (.I0(x3828), .I1(x3829), .I2(x3830), .O(n12362));
  LUT5 #(.INIT(32'h96696996)) lut_n12363 (.I0(x3819), .I1(x3820), .I2(x3821), .I3(n12359), .I4(n12360), .O(n12363));
  LUT5 #(.INIT(32'hFF969600)) lut_n12364 (.I0(x3825), .I1(x3826), .I2(x3827), .I3(n12362), .I4(n12363), .O(n12364));
  LUT3 #(.INIT(8'h96)) lut_n12365 (.I0(n12349), .I1(n12352), .I2(n12353), .O(n12365));
  LUT3 #(.INIT(8'hE8)) lut_n12366 (.I0(n12361), .I1(n12364), .I2(n12365), .O(n12366));
  LUT3 #(.INIT(8'h96)) lut_n12367 (.I0(x3834), .I1(x3835), .I2(x3836), .O(n12367));
  LUT5 #(.INIT(32'h96696996)) lut_n12368 (.I0(x3825), .I1(x3826), .I2(x3827), .I3(n12362), .I4(n12363), .O(n12368));
  LUT5 #(.INIT(32'hFF969600)) lut_n12369 (.I0(x3831), .I1(x3832), .I2(x3833), .I3(n12367), .I4(n12368), .O(n12369));
  LUT3 #(.INIT(8'h96)) lut_n12370 (.I0(x3840), .I1(x3841), .I2(x3842), .O(n12370));
  LUT5 #(.INIT(32'h96696996)) lut_n12371 (.I0(x3831), .I1(x3832), .I2(x3833), .I3(n12367), .I4(n12368), .O(n12371));
  LUT5 #(.INIT(32'hFF969600)) lut_n12372 (.I0(x3837), .I1(x3838), .I2(x3839), .I3(n12370), .I4(n12371), .O(n12372));
  LUT3 #(.INIT(8'h96)) lut_n12373 (.I0(n12361), .I1(n12364), .I2(n12365), .O(n12373));
  LUT3 #(.INIT(8'hE8)) lut_n12374 (.I0(n12369), .I1(n12372), .I2(n12373), .O(n12374));
  LUT3 #(.INIT(8'h96)) lut_n12375 (.I0(n12346), .I1(n12354), .I2(n12355), .O(n12375));
  LUT3 #(.INIT(8'hE8)) lut_n12376 (.I0(n12366), .I1(n12374), .I2(n12375), .O(n12376));
  LUT3 #(.INIT(8'h96)) lut_n12377 (.I0(x3846), .I1(x3847), .I2(x3848), .O(n12377));
  LUT5 #(.INIT(32'h96696996)) lut_n12378 (.I0(x3837), .I1(x3838), .I2(x3839), .I3(n12370), .I4(n12371), .O(n12378));
  LUT5 #(.INIT(32'hFF969600)) lut_n12379 (.I0(x3843), .I1(x3844), .I2(x3845), .I3(n12377), .I4(n12378), .O(n12379));
  LUT3 #(.INIT(8'h96)) lut_n12380 (.I0(x3852), .I1(x3853), .I2(x3854), .O(n12380));
  LUT5 #(.INIT(32'h96696996)) lut_n12381 (.I0(x3843), .I1(x3844), .I2(x3845), .I3(n12377), .I4(n12378), .O(n12381));
  LUT5 #(.INIT(32'hFF969600)) lut_n12382 (.I0(x3849), .I1(x3850), .I2(x3851), .I3(n12380), .I4(n12381), .O(n12382));
  LUT3 #(.INIT(8'h96)) lut_n12383 (.I0(n12369), .I1(n12372), .I2(n12373), .O(n12383));
  LUT3 #(.INIT(8'hE8)) lut_n12384 (.I0(n12379), .I1(n12382), .I2(n12383), .O(n12384));
  LUT3 #(.INIT(8'h96)) lut_n12385 (.I0(x3858), .I1(x3859), .I2(x3860), .O(n12385));
  LUT5 #(.INIT(32'h96696996)) lut_n12386 (.I0(x3849), .I1(x3850), .I2(x3851), .I3(n12380), .I4(n12381), .O(n12386));
  LUT5 #(.INIT(32'hFF969600)) lut_n12387 (.I0(x3855), .I1(x3856), .I2(x3857), .I3(n12385), .I4(n12386), .O(n12387));
  LUT3 #(.INIT(8'h96)) lut_n12388 (.I0(x3864), .I1(x3865), .I2(x3866), .O(n12388));
  LUT5 #(.INIT(32'h96696996)) lut_n12389 (.I0(x3855), .I1(x3856), .I2(x3857), .I3(n12385), .I4(n12386), .O(n12389));
  LUT5 #(.INIT(32'hFF969600)) lut_n12390 (.I0(x3861), .I1(x3862), .I2(x3863), .I3(n12388), .I4(n12389), .O(n12390));
  LUT3 #(.INIT(8'h96)) lut_n12391 (.I0(n12379), .I1(n12382), .I2(n12383), .O(n12391));
  LUT3 #(.INIT(8'hE8)) lut_n12392 (.I0(n12387), .I1(n12390), .I2(n12391), .O(n12392));
  LUT3 #(.INIT(8'h96)) lut_n12393 (.I0(n12366), .I1(n12374), .I2(n12375), .O(n12393));
  LUT3 #(.INIT(8'hE8)) lut_n12394 (.I0(n12384), .I1(n12392), .I2(n12393), .O(n12394));
  LUT3 #(.INIT(8'h96)) lut_n12395 (.I0(n12338), .I1(n12356), .I2(n12357), .O(n12395));
  LUT3 #(.INIT(8'hE8)) lut_n12396 (.I0(n12376), .I1(n12394), .I2(n12395), .O(n12396));
  LUT3 #(.INIT(8'h96)) lut_n12397 (.I0(n12272), .I1(n12310), .I2(n12311), .O(n12397));
  LUT3 #(.INIT(8'hE8)) lut_n12398 (.I0(n12358), .I1(n12396), .I2(n12397), .O(n12398));
  LUT3 #(.INIT(8'h96)) lut_n12399 (.I0(x3870), .I1(x3871), .I2(x3872), .O(n12399));
  LUT5 #(.INIT(32'h96696996)) lut_n12400 (.I0(x3861), .I1(x3862), .I2(x3863), .I3(n12388), .I4(n12389), .O(n12400));
  LUT5 #(.INIT(32'hFF969600)) lut_n12401 (.I0(x3867), .I1(x3868), .I2(x3869), .I3(n12399), .I4(n12400), .O(n12401));
  LUT3 #(.INIT(8'h96)) lut_n12402 (.I0(x3876), .I1(x3877), .I2(x3878), .O(n12402));
  LUT5 #(.INIT(32'h96696996)) lut_n12403 (.I0(x3867), .I1(x3868), .I2(x3869), .I3(n12399), .I4(n12400), .O(n12403));
  LUT5 #(.INIT(32'hFF969600)) lut_n12404 (.I0(x3873), .I1(x3874), .I2(x3875), .I3(n12402), .I4(n12403), .O(n12404));
  LUT3 #(.INIT(8'h96)) lut_n12405 (.I0(n12387), .I1(n12390), .I2(n12391), .O(n12405));
  LUT3 #(.INIT(8'hE8)) lut_n12406 (.I0(n12401), .I1(n12404), .I2(n12405), .O(n12406));
  LUT3 #(.INIT(8'h96)) lut_n12407 (.I0(x3882), .I1(x3883), .I2(x3884), .O(n12407));
  LUT5 #(.INIT(32'h96696996)) lut_n12408 (.I0(x3873), .I1(x3874), .I2(x3875), .I3(n12402), .I4(n12403), .O(n12408));
  LUT5 #(.INIT(32'hFF969600)) lut_n12409 (.I0(x3879), .I1(x3880), .I2(x3881), .I3(n12407), .I4(n12408), .O(n12409));
  LUT3 #(.INIT(8'h96)) lut_n12410 (.I0(x3888), .I1(x3889), .I2(x3890), .O(n12410));
  LUT5 #(.INIT(32'h96696996)) lut_n12411 (.I0(x3879), .I1(x3880), .I2(x3881), .I3(n12407), .I4(n12408), .O(n12411));
  LUT5 #(.INIT(32'hFF969600)) lut_n12412 (.I0(x3885), .I1(x3886), .I2(x3887), .I3(n12410), .I4(n12411), .O(n12412));
  LUT3 #(.INIT(8'h96)) lut_n12413 (.I0(n12401), .I1(n12404), .I2(n12405), .O(n12413));
  LUT3 #(.INIT(8'hE8)) lut_n12414 (.I0(n12409), .I1(n12412), .I2(n12413), .O(n12414));
  LUT3 #(.INIT(8'h96)) lut_n12415 (.I0(n12384), .I1(n12392), .I2(n12393), .O(n12415));
  LUT3 #(.INIT(8'hE8)) lut_n12416 (.I0(n12406), .I1(n12414), .I2(n12415), .O(n12416));
  LUT3 #(.INIT(8'h96)) lut_n12417 (.I0(x3894), .I1(x3895), .I2(x3896), .O(n12417));
  LUT5 #(.INIT(32'h96696996)) lut_n12418 (.I0(x3885), .I1(x3886), .I2(x3887), .I3(n12410), .I4(n12411), .O(n12418));
  LUT5 #(.INIT(32'hFF969600)) lut_n12419 (.I0(x3891), .I1(x3892), .I2(x3893), .I3(n12417), .I4(n12418), .O(n12419));
  LUT3 #(.INIT(8'h96)) lut_n12420 (.I0(x3900), .I1(x3901), .I2(x3902), .O(n12420));
  LUT5 #(.INIT(32'h96696996)) lut_n12421 (.I0(x3891), .I1(x3892), .I2(x3893), .I3(n12417), .I4(n12418), .O(n12421));
  LUT5 #(.INIT(32'hFF969600)) lut_n12422 (.I0(x3897), .I1(x3898), .I2(x3899), .I3(n12420), .I4(n12421), .O(n12422));
  LUT3 #(.INIT(8'h96)) lut_n12423 (.I0(n12409), .I1(n12412), .I2(n12413), .O(n12423));
  LUT3 #(.INIT(8'hE8)) lut_n12424 (.I0(n12419), .I1(n12422), .I2(n12423), .O(n12424));
  LUT3 #(.INIT(8'h96)) lut_n12425 (.I0(x3906), .I1(x3907), .I2(x3908), .O(n12425));
  LUT5 #(.INIT(32'h96696996)) lut_n12426 (.I0(x3897), .I1(x3898), .I2(x3899), .I3(n12420), .I4(n12421), .O(n12426));
  LUT5 #(.INIT(32'hFF969600)) lut_n12427 (.I0(x3903), .I1(x3904), .I2(x3905), .I3(n12425), .I4(n12426), .O(n12427));
  LUT3 #(.INIT(8'h96)) lut_n12428 (.I0(x3912), .I1(x3913), .I2(x3914), .O(n12428));
  LUT5 #(.INIT(32'h96696996)) lut_n12429 (.I0(x3903), .I1(x3904), .I2(x3905), .I3(n12425), .I4(n12426), .O(n12429));
  LUT5 #(.INIT(32'hFF969600)) lut_n12430 (.I0(x3909), .I1(x3910), .I2(x3911), .I3(n12428), .I4(n12429), .O(n12430));
  LUT3 #(.INIT(8'h96)) lut_n12431 (.I0(n12419), .I1(n12422), .I2(n12423), .O(n12431));
  LUT3 #(.INIT(8'hE8)) lut_n12432 (.I0(n12427), .I1(n12430), .I2(n12431), .O(n12432));
  LUT3 #(.INIT(8'h96)) lut_n12433 (.I0(n12406), .I1(n12414), .I2(n12415), .O(n12433));
  LUT3 #(.INIT(8'hE8)) lut_n12434 (.I0(n12424), .I1(n12432), .I2(n12433), .O(n12434));
  LUT3 #(.INIT(8'h96)) lut_n12435 (.I0(n12376), .I1(n12394), .I2(n12395), .O(n12435));
  LUT3 #(.INIT(8'hE8)) lut_n12436 (.I0(n12416), .I1(n12434), .I2(n12435), .O(n12436));
  LUT3 #(.INIT(8'h96)) lut_n12437 (.I0(x3918), .I1(x3919), .I2(x3920), .O(n12437));
  LUT5 #(.INIT(32'h96696996)) lut_n12438 (.I0(x3909), .I1(x3910), .I2(x3911), .I3(n12428), .I4(n12429), .O(n12438));
  LUT5 #(.INIT(32'hFF969600)) lut_n12439 (.I0(x3915), .I1(x3916), .I2(x3917), .I3(n12437), .I4(n12438), .O(n12439));
  LUT3 #(.INIT(8'h96)) lut_n12440 (.I0(x3924), .I1(x3925), .I2(x3926), .O(n12440));
  LUT5 #(.INIT(32'h96696996)) lut_n12441 (.I0(x3915), .I1(x3916), .I2(x3917), .I3(n12437), .I4(n12438), .O(n12441));
  LUT5 #(.INIT(32'hFF969600)) lut_n12442 (.I0(x3921), .I1(x3922), .I2(x3923), .I3(n12440), .I4(n12441), .O(n12442));
  LUT3 #(.INIT(8'h96)) lut_n12443 (.I0(n12427), .I1(n12430), .I2(n12431), .O(n12443));
  LUT3 #(.INIT(8'hE8)) lut_n12444 (.I0(n12439), .I1(n12442), .I2(n12443), .O(n12444));
  LUT3 #(.INIT(8'h96)) lut_n12445 (.I0(x3930), .I1(x3931), .I2(x3932), .O(n12445));
  LUT5 #(.INIT(32'h96696996)) lut_n12446 (.I0(x3921), .I1(x3922), .I2(x3923), .I3(n12440), .I4(n12441), .O(n12446));
  LUT5 #(.INIT(32'hFF969600)) lut_n12447 (.I0(x3927), .I1(x3928), .I2(x3929), .I3(n12445), .I4(n12446), .O(n12447));
  LUT3 #(.INIT(8'h96)) lut_n12448 (.I0(x3936), .I1(x3937), .I2(x3938), .O(n12448));
  LUT5 #(.INIT(32'h96696996)) lut_n12449 (.I0(x3927), .I1(x3928), .I2(x3929), .I3(n12445), .I4(n12446), .O(n12449));
  LUT5 #(.INIT(32'hFF969600)) lut_n12450 (.I0(x3933), .I1(x3934), .I2(x3935), .I3(n12448), .I4(n12449), .O(n12450));
  LUT3 #(.INIT(8'h96)) lut_n12451 (.I0(n12439), .I1(n12442), .I2(n12443), .O(n12451));
  LUT3 #(.INIT(8'hE8)) lut_n12452 (.I0(n12447), .I1(n12450), .I2(n12451), .O(n12452));
  LUT3 #(.INIT(8'h96)) lut_n12453 (.I0(n12424), .I1(n12432), .I2(n12433), .O(n12453));
  LUT3 #(.INIT(8'hE8)) lut_n12454 (.I0(n12444), .I1(n12452), .I2(n12453), .O(n12454));
  LUT3 #(.INIT(8'h96)) lut_n12455 (.I0(x3942), .I1(x3943), .I2(x3944), .O(n12455));
  LUT5 #(.INIT(32'h96696996)) lut_n12456 (.I0(x3933), .I1(x3934), .I2(x3935), .I3(n12448), .I4(n12449), .O(n12456));
  LUT5 #(.INIT(32'hFF969600)) lut_n12457 (.I0(x3939), .I1(x3940), .I2(x3941), .I3(n12455), .I4(n12456), .O(n12457));
  LUT3 #(.INIT(8'h96)) lut_n12458 (.I0(x3948), .I1(x3949), .I2(x3950), .O(n12458));
  LUT5 #(.INIT(32'h96696996)) lut_n12459 (.I0(x3939), .I1(x3940), .I2(x3941), .I3(n12455), .I4(n12456), .O(n12459));
  LUT5 #(.INIT(32'hFF969600)) lut_n12460 (.I0(x3945), .I1(x3946), .I2(x3947), .I3(n12458), .I4(n12459), .O(n12460));
  LUT3 #(.INIT(8'h96)) lut_n12461 (.I0(n12447), .I1(n12450), .I2(n12451), .O(n12461));
  LUT3 #(.INIT(8'hE8)) lut_n12462 (.I0(n12457), .I1(n12460), .I2(n12461), .O(n12462));
  LUT3 #(.INIT(8'h96)) lut_n12463 (.I0(x3954), .I1(x3955), .I2(x3956), .O(n12463));
  LUT5 #(.INIT(32'h96696996)) lut_n12464 (.I0(x3945), .I1(x3946), .I2(x3947), .I3(n12458), .I4(n12459), .O(n12464));
  LUT5 #(.INIT(32'hFF969600)) lut_n12465 (.I0(x3951), .I1(x3952), .I2(x3953), .I3(n12463), .I4(n12464), .O(n12465));
  LUT3 #(.INIT(8'h96)) lut_n12466 (.I0(x3960), .I1(x3961), .I2(x3962), .O(n12466));
  LUT5 #(.INIT(32'h96696996)) lut_n12467 (.I0(x3951), .I1(x3952), .I2(x3953), .I3(n12463), .I4(n12464), .O(n12467));
  LUT5 #(.INIT(32'hFF969600)) lut_n12468 (.I0(x3957), .I1(x3958), .I2(x3959), .I3(n12466), .I4(n12467), .O(n12468));
  LUT3 #(.INIT(8'h96)) lut_n12469 (.I0(n12457), .I1(n12460), .I2(n12461), .O(n12469));
  LUT3 #(.INIT(8'hE8)) lut_n12470 (.I0(n12465), .I1(n12468), .I2(n12469), .O(n12470));
  LUT3 #(.INIT(8'h96)) lut_n12471 (.I0(n12444), .I1(n12452), .I2(n12453), .O(n12471));
  LUT3 #(.INIT(8'hE8)) lut_n12472 (.I0(n12462), .I1(n12470), .I2(n12471), .O(n12472));
  LUT3 #(.INIT(8'h96)) lut_n12473 (.I0(n12416), .I1(n12434), .I2(n12435), .O(n12473));
  LUT3 #(.INIT(8'hE8)) lut_n12474 (.I0(n12454), .I1(n12472), .I2(n12473), .O(n12474));
  LUT3 #(.INIT(8'h96)) lut_n12475 (.I0(n12358), .I1(n12396), .I2(n12397), .O(n12475));
  LUT3 #(.INIT(8'hE8)) lut_n12476 (.I0(n12436), .I1(n12474), .I2(n12475), .O(n12476));
  LUT3 #(.INIT(8'h96)) lut_n12477 (.I0(n12234), .I1(n12312), .I2(n12313), .O(n12477));
  LUT3 #(.INIT(8'hE8)) lut_n12478 (.I0(n12398), .I1(n12476), .I2(n12477), .O(n12478));
  LUT3 #(.INIT(8'h96)) lut_n12479 (.I0(x3966), .I1(x3967), .I2(x3968), .O(n12479));
  LUT5 #(.INIT(32'h96696996)) lut_n12480 (.I0(x3957), .I1(x3958), .I2(x3959), .I3(n12466), .I4(n12467), .O(n12480));
  LUT5 #(.INIT(32'hFF969600)) lut_n12481 (.I0(x3963), .I1(x3964), .I2(x3965), .I3(n12479), .I4(n12480), .O(n12481));
  LUT3 #(.INIT(8'h96)) lut_n12482 (.I0(x3972), .I1(x3973), .I2(x3974), .O(n12482));
  LUT5 #(.INIT(32'h96696996)) lut_n12483 (.I0(x3963), .I1(x3964), .I2(x3965), .I3(n12479), .I4(n12480), .O(n12483));
  LUT5 #(.INIT(32'hFF969600)) lut_n12484 (.I0(x3969), .I1(x3970), .I2(x3971), .I3(n12482), .I4(n12483), .O(n12484));
  LUT3 #(.INIT(8'h96)) lut_n12485 (.I0(n12465), .I1(n12468), .I2(n12469), .O(n12485));
  LUT3 #(.INIT(8'hE8)) lut_n12486 (.I0(n12481), .I1(n12484), .I2(n12485), .O(n12486));
  LUT3 #(.INIT(8'h96)) lut_n12487 (.I0(x3978), .I1(x3979), .I2(x3980), .O(n12487));
  LUT5 #(.INIT(32'h96696996)) lut_n12488 (.I0(x3969), .I1(x3970), .I2(x3971), .I3(n12482), .I4(n12483), .O(n12488));
  LUT5 #(.INIT(32'hFF969600)) lut_n12489 (.I0(x3975), .I1(x3976), .I2(x3977), .I3(n12487), .I4(n12488), .O(n12489));
  LUT3 #(.INIT(8'h96)) lut_n12490 (.I0(x3984), .I1(x3985), .I2(x3986), .O(n12490));
  LUT5 #(.INIT(32'h96696996)) lut_n12491 (.I0(x3975), .I1(x3976), .I2(x3977), .I3(n12487), .I4(n12488), .O(n12491));
  LUT5 #(.INIT(32'hFF969600)) lut_n12492 (.I0(x3981), .I1(x3982), .I2(x3983), .I3(n12490), .I4(n12491), .O(n12492));
  LUT3 #(.INIT(8'h96)) lut_n12493 (.I0(n12481), .I1(n12484), .I2(n12485), .O(n12493));
  LUT3 #(.INIT(8'hE8)) lut_n12494 (.I0(n12489), .I1(n12492), .I2(n12493), .O(n12494));
  LUT3 #(.INIT(8'h96)) lut_n12495 (.I0(n12462), .I1(n12470), .I2(n12471), .O(n12495));
  LUT3 #(.INIT(8'hE8)) lut_n12496 (.I0(n12486), .I1(n12494), .I2(n12495), .O(n12496));
  LUT3 #(.INIT(8'h96)) lut_n12497 (.I0(x3990), .I1(x3991), .I2(x3992), .O(n12497));
  LUT5 #(.INIT(32'h96696996)) lut_n12498 (.I0(x3981), .I1(x3982), .I2(x3983), .I3(n12490), .I4(n12491), .O(n12498));
  LUT5 #(.INIT(32'hFF969600)) lut_n12499 (.I0(x3987), .I1(x3988), .I2(x3989), .I3(n12497), .I4(n12498), .O(n12499));
  LUT3 #(.INIT(8'h96)) lut_n12500 (.I0(x3996), .I1(x3997), .I2(x3998), .O(n12500));
  LUT5 #(.INIT(32'h96696996)) lut_n12501 (.I0(x3987), .I1(x3988), .I2(x3989), .I3(n12497), .I4(n12498), .O(n12501));
  LUT5 #(.INIT(32'hFF969600)) lut_n12502 (.I0(x3993), .I1(x3994), .I2(x3995), .I3(n12500), .I4(n12501), .O(n12502));
  LUT3 #(.INIT(8'h96)) lut_n12503 (.I0(n12489), .I1(n12492), .I2(n12493), .O(n12503));
  LUT3 #(.INIT(8'hE8)) lut_n12504 (.I0(n12499), .I1(n12502), .I2(n12503), .O(n12504));
  LUT3 #(.INIT(8'h96)) lut_n12505 (.I0(x4002), .I1(x4003), .I2(x4004), .O(n12505));
  LUT5 #(.INIT(32'h96696996)) lut_n12506 (.I0(x3993), .I1(x3994), .I2(x3995), .I3(n12500), .I4(n12501), .O(n12506));
  LUT5 #(.INIT(32'hFF969600)) lut_n12507 (.I0(x3999), .I1(x4000), .I2(x4001), .I3(n12505), .I4(n12506), .O(n12507));
  LUT3 #(.INIT(8'h96)) lut_n12508 (.I0(x4008), .I1(x4009), .I2(x4010), .O(n12508));
  LUT5 #(.INIT(32'h96696996)) lut_n12509 (.I0(x3999), .I1(x4000), .I2(x4001), .I3(n12505), .I4(n12506), .O(n12509));
  LUT5 #(.INIT(32'hFF969600)) lut_n12510 (.I0(x4005), .I1(x4006), .I2(x4007), .I3(n12508), .I4(n12509), .O(n12510));
  LUT3 #(.INIT(8'h96)) lut_n12511 (.I0(n12499), .I1(n12502), .I2(n12503), .O(n12511));
  LUT3 #(.INIT(8'hE8)) lut_n12512 (.I0(n12507), .I1(n12510), .I2(n12511), .O(n12512));
  LUT3 #(.INIT(8'h96)) lut_n12513 (.I0(n12486), .I1(n12494), .I2(n12495), .O(n12513));
  LUT3 #(.INIT(8'hE8)) lut_n12514 (.I0(n12504), .I1(n12512), .I2(n12513), .O(n12514));
  LUT3 #(.INIT(8'h96)) lut_n12515 (.I0(n12454), .I1(n12472), .I2(n12473), .O(n12515));
  LUT3 #(.INIT(8'hE8)) lut_n12516 (.I0(n12496), .I1(n12514), .I2(n12515), .O(n12516));
  LUT3 #(.INIT(8'h96)) lut_n12517 (.I0(x4014), .I1(x4015), .I2(x4016), .O(n12517));
  LUT5 #(.INIT(32'h96696996)) lut_n12518 (.I0(x4005), .I1(x4006), .I2(x4007), .I3(n12508), .I4(n12509), .O(n12518));
  LUT5 #(.INIT(32'hFF969600)) lut_n12519 (.I0(x4011), .I1(x4012), .I2(x4013), .I3(n12517), .I4(n12518), .O(n12519));
  LUT3 #(.INIT(8'h96)) lut_n12520 (.I0(x4020), .I1(x4021), .I2(x4022), .O(n12520));
  LUT5 #(.INIT(32'h96696996)) lut_n12521 (.I0(x4011), .I1(x4012), .I2(x4013), .I3(n12517), .I4(n12518), .O(n12521));
  LUT5 #(.INIT(32'hFF969600)) lut_n12522 (.I0(x4017), .I1(x4018), .I2(x4019), .I3(n12520), .I4(n12521), .O(n12522));
  LUT3 #(.INIT(8'h96)) lut_n12523 (.I0(n12507), .I1(n12510), .I2(n12511), .O(n12523));
  LUT3 #(.INIT(8'hE8)) lut_n12524 (.I0(n12519), .I1(n12522), .I2(n12523), .O(n12524));
  LUT3 #(.INIT(8'h96)) lut_n12525 (.I0(x4026), .I1(x4027), .I2(x4028), .O(n12525));
  LUT5 #(.INIT(32'h96696996)) lut_n12526 (.I0(x4017), .I1(x4018), .I2(x4019), .I3(n12520), .I4(n12521), .O(n12526));
  LUT5 #(.INIT(32'hFF969600)) lut_n12527 (.I0(x4023), .I1(x4024), .I2(x4025), .I3(n12525), .I4(n12526), .O(n12527));
  LUT3 #(.INIT(8'h96)) lut_n12528 (.I0(x4032), .I1(x4033), .I2(x4034), .O(n12528));
  LUT5 #(.INIT(32'h96696996)) lut_n12529 (.I0(x4023), .I1(x4024), .I2(x4025), .I3(n12525), .I4(n12526), .O(n12529));
  LUT5 #(.INIT(32'hFF969600)) lut_n12530 (.I0(x4029), .I1(x4030), .I2(x4031), .I3(n12528), .I4(n12529), .O(n12530));
  LUT3 #(.INIT(8'h96)) lut_n12531 (.I0(n12519), .I1(n12522), .I2(n12523), .O(n12531));
  LUT3 #(.INIT(8'hE8)) lut_n12532 (.I0(n12527), .I1(n12530), .I2(n12531), .O(n12532));
  LUT3 #(.INIT(8'h96)) lut_n12533 (.I0(n12504), .I1(n12512), .I2(n12513), .O(n12533));
  LUT3 #(.INIT(8'hE8)) lut_n12534 (.I0(n12524), .I1(n12532), .I2(n12533), .O(n12534));
  LUT3 #(.INIT(8'h96)) lut_n12535 (.I0(x4038), .I1(x4039), .I2(x4040), .O(n12535));
  LUT5 #(.INIT(32'h96696996)) lut_n12536 (.I0(x4029), .I1(x4030), .I2(x4031), .I3(n12528), .I4(n12529), .O(n12536));
  LUT5 #(.INIT(32'hFF969600)) lut_n12537 (.I0(x4035), .I1(x4036), .I2(x4037), .I3(n12535), .I4(n12536), .O(n12537));
  LUT3 #(.INIT(8'h96)) lut_n12538 (.I0(x4044), .I1(x4045), .I2(x4046), .O(n12538));
  LUT5 #(.INIT(32'h96696996)) lut_n12539 (.I0(x4035), .I1(x4036), .I2(x4037), .I3(n12535), .I4(n12536), .O(n12539));
  LUT5 #(.INIT(32'hFF969600)) lut_n12540 (.I0(x4041), .I1(x4042), .I2(x4043), .I3(n12538), .I4(n12539), .O(n12540));
  LUT3 #(.INIT(8'h96)) lut_n12541 (.I0(n12527), .I1(n12530), .I2(n12531), .O(n12541));
  LUT3 #(.INIT(8'hE8)) lut_n12542 (.I0(n12537), .I1(n12540), .I2(n12541), .O(n12542));
  LUT3 #(.INIT(8'h96)) lut_n12543 (.I0(x4050), .I1(x4051), .I2(x4052), .O(n12543));
  LUT5 #(.INIT(32'h96696996)) lut_n12544 (.I0(x4041), .I1(x4042), .I2(x4043), .I3(n12538), .I4(n12539), .O(n12544));
  LUT5 #(.INIT(32'hFF969600)) lut_n12545 (.I0(x4047), .I1(x4048), .I2(x4049), .I3(n12543), .I4(n12544), .O(n12545));
  LUT3 #(.INIT(8'h96)) lut_n12546 (.I0(x4056), .I1(x4057), .I2(x4058), .O(n12546));
  LUT5 #(.INIT(32'h96696996)) lut_n12547 (.I0(x4047), .I1(x4048), .I2(x4049), .I3(n12543), .I4(n12544), .O(n12547));
  LUT5 #(.INIT(32'hFF969600)) lut_n12548 (.I0(x4053), .I1(x4054), .I2(x4055), .I3(n12546), .I4(n12547), .O(n12548));
  LUT3 #(.INIT(8'h96)) lut_n12549 (.I0(n12537), .I1(n12540), .I2(n12541), .O(n12549));
  LUT3 #(.INIT(8'hE8)) lut_n12550 (.I0(n12545), .I1(n12548), .I2(n12549), .O(n12550));
  LUT3 #(.INIT(8'h96)) lut_n12551 (.I0(n12524), .I1(n12532), .I2(n12533), .O(n12551));
  LUT3 #(.INIT(8'hE8)) lut_n12552 (.I0(n12542), .I1(n12550), .I2(n12551), .O(n12552));
  LUT3 #(.INIT(8'h96)) lut_n12553 (.I0(n12496), .I1(n12514), .I2(n12515), .O(n12553));
  LUT3 #(.INIT(8'hE8)) lut_n12554 (.I0(n12534), .I1(n12552), .I2(n12553), .O(n12554));
  LUT3 #(.INIT(8'h96)) lut_n12555 (.I0(n12436), .I1(n12474), .I2(n12475), .O(n12555));
  LUT3 #(.INIT(8'hE8)) lut_n12556 (.I0(n12516), .I1(n12554), .I2(n12555), .O(n12556));
  LUT3 #(.INIT(8'h96)) lut_n12557 (.I0(x4062), .I1(x4063), .I2(x4064), .O(n12557));
  LUT5 #(.INIT(32'h96696996)) lut_n12558 (.I0(x4053), .I1(x4054), .I2(x4055), .I3(n12546), .I4(n12547), .O(n12558));
  LUT5 #(.INIT(32'hFF969600)) lut_n12559 (.I0(x4059), .I1(x4060), .I2(x4061), .I3(n12557), .I4(n12558), .O(n12559));
  LUT3 #(.INIT(8'h96)) lut_n12560 (.I0(x4068), .I1(x4069), .I2(x4070), .O(n12560));
  LUT5 #(.INIT(32'h96696996)) lut_n12561 (.I0(x4059), .I1(x4060), .I2(x4061), .I3(n12557), .I4(n12558), .O(n12561));
  LUT5 #(.INIT(32'hFF969600)) lut_n12562 (.I0(x4065), .I1(x4066), .I2(x4067), .I3(n12560), .I4(n12561), .O(n12562));
  LUT3 #(.INIT(8'h96)) lut_n12563 (.I0(n12545), .I1(n12548), .I2(n12549), .O(n12563));
  LUT3 #(.INIT(8'hE8)) lut_n12564 (.I0(n12559), .I1(n12562), .I2(n12563), .O(n12564));
  LUT3 #(.INIT(8'h96)) lut_n12565 (.I0(x4074), .I1(x4075), .I2(x4076), .O(n12565));
  LUT5 #(.INIT(32'h96696996)) lut_n12566 (.I0(x4065), .I1(x4066), .I2(x4067), .I3(n12560), .I4(n12561), .O(n12566));
  LUT5 #(.INIT(32'hFF969600)) lut_n12567 (.I0(x4071), .I1(x4072), .I2(x4073), .I3(n12565), .I4(n12566), .O(n12567));
  LUT3 #(.INIT(8'h96)) lut_n12568 (.I0(x4080), .I1(x4081), .I2(x4082), .O(n12568));
  LUT5 #(.INIT(32'h96696996)) lut_n12569 (.I0(x4071), .I1(x4072), .I2(x4073), .I3(n12565), .I4(n12566), .O(n12569));
  LUT5 #(.INIT(32'hFF969600)) lut_n12570 (.I0(x4077), .I1(x4078), .I2(x4079), .I3(n12568), .I4(n12569), .O(n12570));
  LUT3 #(.INIT(8'h96)) lut_n12571 (.I0(n12559), .I1(n12562), .I2(n12563), .O(n12571));
  LUT3 #(.INIT(8'hE8)) lut_n12572 (.I0(n12567), .I1(n12570), .I2(n12571), .O(n12572));
  LUT3 #(.INIT(8'h96)) lut_n12573 (.I0(n12542), .I1(n12550), .I2(n12551), .O(n12573));
  LUT3 #(.INIT(8'hE8)) lut_n12574 (.I0(n12564), .I1(n12572), .I2(n12573), .O(n12574));
  LUT3 #(.INIT(8'h96)) lut_n12575 (.I0(x4086), .I1(x4087), .I2(x4088), .O(n12575));
  LUT5 #(.INIT(32'h96696996)) lut_n12576 (.I0(x4077), .I1(x4078), .I2(x4079), .I3(n12568), .I4(n12569), .O(n12576));
  LUT5 #(.INIT(32'hFF969600)) lut_n12577 (.I0(x4083), .I1(x4084), .I2(x4085), .I3(n12575), .I4(n12576), .O(n12577));
  LUT3 #(.INIT(8'h96)) lut_n12578 (.I0(x4092), .I1(x4093), .I2(x4094), .O(n12578));
  LUT5 #(.INIT(32'h96696996)) lut_n12579 (.I0(x4083), .I1(x4084), .I2(x4085), .I3(n12575), .I4(n12576), .O(n12579));
  LUT5 #(.INIT(32'hFF969600)) lut_n12580 (.I0(x4089), .I1(x4090), .I2(x4091), .I3(n12578), .I4(n12579), .O(n12580));
  LUT3 #(.INIT(8'h96)) lut_n12581 (.I0(n12567), .I1(n12570), .I2(n12571), .O(n12581));
  LUT3 #(.INIT(8'hE8)) lut_n12582 (.I0(n12577), .I1(n12580), .I2(n12581), .O(n12582));
  LUT3 #(.INIT(8'h96)) lut_n12583 (.I0(x4098), .I1(x4099), .I2(x4100), .O(n12583));
  LUT5 #(.INIT(32'h96696996)) lut_n12584 (.I0(x4089), .I1(x4090), .I2(x4091), .I3(n12578), .I4(n12579), .O(n12584));
  LUT5 #(.INIT(32'hFF969600)) lut_n12585 (.I0(x4095), .I1(x4096), .I2(x4097), .I3(n12583), .I4(n12584), .O(n12585));
  LUT3 #(.INIT(8'h96)) lut_n12586 (.I0(x4104), .I1(x4105), .I2(x4106), .O(n12586));
  LUT5 #(.INIT(32'h96696996)) lut_n12587 (.I0(x4095), .I1(x4096), .I2(x4097), .I3(n12583), .I4(n12584), .O(n12587));
  LUT5 #(.INIT(32'hFF969600)) lut_n12588 (.I0(x4101), .I1(x4102), .I2(x4103), .I3(n12586), .I4(n12587), .O(n12588));
  LUT3 #(.INIT(8'h96)) lut_n12589 (.I0(n12577), .I1(n12580), .I2(n12581), .O(n12589));
  LUT3 #(.INIT(8'hE8)) lut_n12590 (.I0(n12585), .I1(n12588), .I2(n12589), .O(n12590));
  LUT3 #(.INIT(8'h96)) lut_n12591 (.I0(n12564), .I1(n12572), .I2(n12573), .O(n12591));
  LUT3 #(.INIT(8'hE8)) lut_n12592 (.I0(n12582), .I1(n12590), .I2(n12591), .O(n12592));
  LUT3 #(.INIT(8'h96)) lut_n12593 (.I0(n12534), .I1(n12552), .I2(n12553), .O(n12593));
  LUT3 #(.INIT(8'hE8)) lut_n12594 (.I0(n12574), .I1(n12592), .I2(n12593), .O(n12594));
  LUT3 #(.INIT(8'h96)) lut_n12595 (.I0(x4110), .I1(x4111), .I2(x4112), .O(n12595));
  LUT5 #(.INIT(32'h96696996)) lut_n12596 (.I0(x4101), .I1(x4102), .I2(x4103), .I3(n12586), .I4(n12587), .O(n12596));
  LUT5 #(.INIT(32'hFF969600)) lut_n12597 (.I0(x4107), .I1(x4108), .I2(x4109), .I3(n12595), .I4(n12596), .O(n12597));
  LUT3 #(.INIT(8'h96)) lut_n12598 (.I0(x4116), .I1(x4117), .I2(x4118), .O(n12598));
  LUT5 #(.INIT(32'h96696996)) lut_n12599 (.I0(x4107), .I1(x4108), .I2(x4109), .I3(n12595), .I4(n12596), .O(n12599));
  LUT5 #(.INIT(32'hFF969600)) lut_n12600 (.I0(x4113), .I1(x4114), .I2(x4115), .I3(n12598), .I4(n12599), .O(n12600));
  LUT3 #(.INIT(8'h96)) lut_n12601 (.I0(n12585), .I1(n12588), .I2(n12589), .O(n12601));
  LUT3 #(.INIT(8'hE8)) lut_n12602 (.I0(n12597), .I1(n12600), .I2(n12601), .O(n12602));
  LUT3 #(.INIT(8'h96)) lut_n12603 (.I0(x4122), .I1(x4123), .I2(x4124), .O(n12603));
  LUT5 #(.INIT(32'h96696996)) lut_n12604 (.I0(x4113), .I1(x4114), .I2(x4115), .I3(n12598), .I4(n12599), .O(n12604));
  LUT5 #(.INIT(32'hFF969600)) lut_n12605 (.I0(x4119), .I1(x4120), .I2(x4121), .I3(n12603), .I4(n12604), .O(n12605));
  LUT3 #(.INIT(8'h96)) lut_n12606 (.I0(x4128), .I1(x4129), .I2(x4130), .O(n12606));
  LUT5 #(.INIT(32'h96696996)) lut_n12607 (.I0(x4119), .I1(x4120), .I2(x4121), .I3(n12603), .I4(n12604), .O(n12607));
  LUT5 #(.INIT(32'hFF969600)) lut_n12608 (.I0(x4125), .I1(x4126), .I2(x4127), .I3(n12606), .I4(n12607), .O(n12608));
  LUT3 #(.INIT(8'h96)) lut_n12609 (.I0(n12597), .I1(n12600), .I2(n12601), .O(n12609));
  LUT3 #(.INIT(8'hE8)) lut_n12610 (.I0(n12605), .I1(n12608), .I2(n12609), .O(n12610));
  LUT3 #(.INIT(8'h96)) lut_n12611 (.I0(n12582), .I1(n12590), .I2(n12591), .O(n12611));
  LUT3 #(.INIT(8'hE8)) lut_n12612 (.I0(n12602), .I1(n12610), .I2(n12611), .O(n12612));
  LUT3 #(.INIT(8'h96)) lut_n12613 (.I0(x4134), .I1(x4135), .I2(x4136), .O(n12613));
  LUT5 #(.INIT(32'h96696996)) lut_n12614 (.I0(x4125), .I1(x4126), .I2(x4127), .I3(n12606), .I4(n12607), .O(n12614));
  LUT5 #(.INIT(32'hFF969600)) lut_n12615 (.I0(x4131), .I1(x4132), .I2(x4133), .I3(n12613), .I4(n12614), .O(n12615));
  LUT3 #(.INIT(8'h96)) lut_n12616 (.I0(x4140), .I1(x4141), .I2(x4142), .O(n12616));
  LUT5 #(.INIT(32'h96696996)) lut_n12617 (.I0(x4131), .I1(x4132), .I2(x4133), .I3(n12613), .I4(n12614), .O(n12617));
  LUT5 #(.INIT(32'hFF969600)) lut_n12618 (.I0(x4137), .I1(x4138), .I2(x4139), .I3(n12616), .I4(n12617), .O(n12618));
  LUT3 #(.INIT(8'h96)) lut_n12619 (.I0(n12605), .I1(n12608), .I2(n12609), .O(n12619));
  LUT3 #(.INIT(8'hE8)) lut_n12620 (.I0(n12615), .I1(n12618), .I2(n12619), .O(n12620));
  LUT3 #(.INIT(8'h96)) lut_n12621 (.I0(x4146), .I1(x4147), .I2(x4148), .O(n12621));
  LUT5 #(.INIT(32'h96696996)) lut_n12622 (.I0(x4137), .I1(x4138), .I2(x4139), .I3(n12616), .I4(n12617), .O(n12622));
  LUT5 #(.INIT(32'hFF969600)) lut_n12623 (.I0(x4143), .I1(x4144), .I2(x4145), .I3(n12621), .I4(n12622), .O(n12623));
  LUT3 #(.INIT(8'h96)) lut_n12624 (.I0(x4152), .I1(x4153), .I2(x4154), .O(n12624));
  LUT5 #(.INIT(32'h96696996)) lut_n12625 (.I0(x4143), .I1(x4144), .I2(x4145), .I3(n12621), .I4(n12622), .O(n12625));
  LUT5 #(.INIT(32'hFF969600)) lut_n12626 (.I0(x4149), .I1(x4150), .I2(x4151), .I3(n12624), .I4(n12625), .O(n12626));
  LUT3 #(.INIT(8'h96)) lut_n12627 (.I0(n12615), .I1(n12618), .I2(n12619), .O(n12627));
  LUT3 #(.INIT(8'hE8)) lut_n12628 (.I0(n12623), .I1(n12626), .I2(n12627), .O(n12628));
  LUT3 #(.INIT(8'h96)) lut_n12629 (.I0(n12602), .I1(n12610), .I2(n12611), .O(n12629));
  LUT3 #(.INIT(8'hE8)) lut_n12630 (.I0(n12620), .I1(n12628), .I2(n12629), .O(n12630));
  LUT3 #(.INIT(8'h96)) lut_n12631 (.I0(n12574), .I1(n12592), .I2(n12593), .O(n12631));
  LUT3 #(.INIT(8'hE8)) lut_n12632 (.I0(n12612), .I1(n12630), .I2(n12631), .O(n12632));
  LUT3 #(.INIT(8'h96)) lut_n12633 (.I0(n12516), .I1(n12554), .I2(n12555), .O(n12633));
  LUT3 #(.INIT(8'hE8)) lut_n12634 (.I0(n12594), .I1(n12632), .I2(n12633), .O(n12634));
  LUT3 #(.INIT(8'h96)) lut_n12635 (.I0(n12398), .I1(n12476), .I2(n12477), .O(n12635));
  LUT3 #(.INIT(8'hE8)) lut_n12636 (.I0(n12556), .I1(n12634), .I2(n12635), .O(n12636));
  LUT3 #(.INIT(8'h96)) lut_n12637 (.I0(n12156), .I1(n12314), .I2(n12315), .O(n12637));
  LUT3 #(.INIT(8'hE8)) lut_n12638 (.I0(n12478), .I1(n12636), .I2(n12637), .O(n12638));
  LUT3 #(.INIT(8'h96)) lut_n12639 (.I0(x4158), .I1(x4159), .I2(x4160), .O(n12639));
  LUT5 #(.INIT(32'h96696996)) lut_n12640 (.I0(x4149), .I1(x4150), .I2(x4151), .I3(n12624), .I4(n12625), .O(n12640));
  LUT5 #(.INIT(32'hFF969600)) lut_n12641 (.I0(x4155), .I1(x4156), .I2(x4157), .I3(n12639), .I4(n12640), .O(n12641));
  LUT3 #(.INIT(8'h96)) lut_n12642 (.I0(x4164), .I1(x4165), .I2(x4166), .O(n12642));
  LUT5 #(.INIT(32'h96696996)) lut_n12643 (.I0(x4155), .I1(x4156), .I2(x4157), .I3(n12639), .I4(n12640), .O(n12643));
  LUT5 #(.INIT(32'hFF969600)) lut_n12644 (.I0(x4161), .I1(x4162), .I2(x4163), .I3(n12642), .I4(n12643), .O(n12644));
  LUT3 #(.INIT(8'h96)) lut_n12645 (.I0(n12623), .I1(n12626), .I2(n12627), .O(n12645));
  LUT3 #(.INIT(8'hE8)) lut_n12646 (.I0(n12641), .I1(n12644), .I2(n12645), .O(n12646));
  LUT3 #(.INIT(8'h96)) lut_n12647 (.I0(x4170), .I1(x4171), .I2(x4172), .O(n12647));
  LUT5 #(.INIT(32'h96696996)) lut_n12648 (.I0(x4161), .I1(x4162), .I2(x4163), .I3(n12642), .I4(n12643), .O(n12648));
  LUT5 #(.INIT(32'hFF969600)) lut_n12649 (.I0(x4167), .I1(x4168), .I2(x4169), .I3(n12647), .I4(n12648), .O(n12649));
  LUT3 #(.INIT(8'h96)) lut_n12650 (.I0(x4176), .I1(x4177), .I2(x4178), .O(n12650));
  LUT5 #(.INIT(32'h96696996)) lut_n12651 (.I0(x4167), .I1(x4168), .I2(x4169), .I3(n12647), .I4(n12648), .O(n12651));
  LUT5 #(.INIT(32'hFF969600)) lut_n12652 (.I0(x4173), .I1(x4174), .I2(x4175), .I3(n12650), .I4(n12651), .O(n12652));
  LUT3 #(.INIT(8'h96)) lut_n12653 (.I0(n12641), .I1(n12644), .I2(n12645), .O(n12653));
  LUT3 #(.INIT(8'hE8)) lut_n12654 (.I0(n12649), .I1(n12652), .I2(n12653), .O(n12654));
  LUT3 #(.INIT(8'h96)) lut_n12655 (.I0(n12620), .I1(n12628), .I2(n12629), .O(n12655));
  LUT3 #(.INIT(8'hE8)) lut_n12656 (.I0(n12646), .I1(n12654), .I2(n12655), .O(n12656));
  LUT3 #(.INIT(8'h96)) lut_n12657 (.I0(x4182), .I1(x4183), .I2(x4184), .O(n12657));
  LUT5 #(.INIT(32'h96696996)) lut_n12658 (.I0(x4173), .I1(x4174), .I2(x4175), .I3(n12650), .I4(n12651), .O(n12658));
  LUT5 #(.INIT(32'hFF969600)) lut_n12659 (.I0(x4179), .I1(x4180), .I2(x4181), .I3(n12657), .I4(n12658), .O(n12659));
  LUT3 #(.INIT(8'h96)) lut_n12660 (.I0(x4188), .I1(x4189), .I2(x4190), .O(n12660));
  LUT5 #(.INIT(32'h96696996)) lut_n12661 (.I0(x4179), .I1(x4180), .I2(x4181), .I3(n12657), .I4(n12658), .O(n12661));
  LUT5 #(.INIT(32'hFF969600)) lut_n12662 (.I0(x4185), .I1(x4186), .I2(x4187), .I3(n12660), .I4(n12661), .O(n12662));
  LUT3 #(.INIT(8'h96)) lut_n12663 (.I0(n12649), .I1(n12652), .I2(n12653), .O(n12663));
  LUT3 #(.INIT(8'hE8)) lut_n12664 (.I0(n12659), .I1(n12662), .I2(n12663), .O(n12664));
  LUT3 #(.INIT(8'h96)) lut_n12665 (.I0(x4194), .I1(x4195), .I2(x4196), .O(n12665));
  LUT5 #(.INIT(32'h96696996)) lut_n12666 (.I0(x4185), .I1(x4186), .I2(x4187), .I3(n12660), .I4(n12661), .O(n12666));
  LUT5 #(.INIT(32'hFF969600)) lut_n12667 (.I0(x4191), .I1(x4192), .I2(x4193), .I3(n12665), .I4(n12666), .O(n12667));
  LUT3 #(.INIT(8'h96)) lut_n12668 (.I0(x4200), .I1(x4201), .I2(x4202), .O(n12668));
  LUT5 #(.INIT(32'h96696996)) lut_n12669 (.I0(x4191), .I1(x4192), .I2(x4193), .I3(n12665), .I4(n12666), .O(n12669));
  LUT5 #(.INIT(32'hFF969600)) lut_n12670 (.I0(x4197), .I1(x4198), .I2(x4199), .I3(n12668), .I4(n12669), .O(n12670));
  LUT3 #(.INIT(8'h96)) lut_n12671 (.I0(n12659), .I1(n12662), .I2(n12663), .O(n12671));
  LUT3 #(.INIT(8'hE8)) lut_n12672 (.I0(n12667), .I1(n12670), .I2(n12671), .O(n12672));
  LUT3 #(.INIT(8'h96)) lut_n12673 (.I0(n12646), .I1(n12654), .I2(n12655), .O(n12673));
  LUT3 #(.INIT(8'hE8)) lut_n12674 (.I0(n12664), .I1(n12672), .I2(n12673), .O(n12674));
  LUT3 #(.INIT(8'h96)) lut_n12675 (.I0(n12612), .I1(n12630), .I2(n12631), .O(n12675));
  LUT3 #(.INIT(8'hE8)) lut_n12676 (.I0(n12656), .I1(n12674), .I2(n12675), .O(n12676));
  LUT3 #(.INIT(8'h96)) lut_n12677 (.I0(x4206), .I1(x4207), .I2(x4208), .O(n12677));
  LUT5 #(.INIT(32'h96696996)) lut_n12678 (.I0(x4197), .I1(x4198), .I2(x4199), .I3(n12668), .I4(n12669), .O(n12678));
  LUT5 #(.INIT(32'hFF969600)) lut_n12679 (.I0(x4203), .I1(x4204), .I2(x4205), .I3(n12677), .I4(n12678), .O(n12679));
  LUT3 #(.INIT(8'h96)) lut_n12680 (.I0(x4212), .I1(x4213), .I2(x4214), .O(n12680));
  LUT5 #(.INIT(32'h96696996)) lut_n12681 (.I0(x4203), .I1(x4204), .I2(x4205), .I3(n12677), .I4(n12678), .O(n12681));
  LUT5 #(.INIT(32'hFF969600)) lut_n12682 (.I0(x4209), .I1(x4210), .I2(x4211), .I3(n12680), .I4(n12681), .O(n12682));
  LUT3 #(.INIT(8'h96)) lut_n12683 (.I0(n12667), .I1(n12670), .I2(n12671), .O(n12683));
  LUT3 #(.INIT(8'hE8)) lut_n12684 (.I0(n12679), .I1(n12682), .I2(n12683), .O(n12684));
  LUT3 #(.INIT(8'h96)) lut_n12685 (.I0(x4218), .I1(x4219), .I2(x4220), .O(n12685));
  LUT5 #(.INIT(32'h96696996)) lut_n12686 (.I0(x4209), .I1(x4210), .I2(x4211), .I3(n12680), .I4(n12681), .O(n12686));
  LUT5 #(.INIT(32'hFF969600)) lut_n12687 (.I0(x4215), .I1(x4216), .I2(x4217), .I3(n12685), .I4(n12686), .O(n12687));
  LUT3 #(.INIT(8'h96)) lut_n12688 (.I0(x4224), .I1(x4225), .I2(x4226), .O(n12688));
  LUT5 #(.INIT(32'h96696996)) lut_n12689 (.I0(x4215), .I1(x4216), .I2(x4217), .I3(n12685), .I4(n12686), .O(n12689));
  LUT5 #(.INIT(32'hFF969600)) lut_n12690 (.I0(x4221), .I1(x4222), .I2(x4223), .I3(n12688), .I4(n12689), .O(n12690));
  LUT3 #(.INIT(8'h96)) lut_n12691 (.I0(n12679), .I1(n12682), .I2(n12683), .O(n12691));
  LUT3 #(.INIT(8'hE8)) lut_n12692 (.I0(n12687), .I1(n12690), .I2(n12691), .O(n12692));
  LUT3 #(.INIT(8'h96)) lut_n12693 (.I0(n12664), .I1(n12672), .I2(n12673), .O(n12693));
  LUT3 #(.INIT(8'hE8)) lut_n12694 (.I0(n12684), .I1(n12692), .I2(n12693), .O(n12694));
  LUT3 #(.INIT(8'h96)) lut_n12695 (.I0(x4230), .I1(x4231), .I2(x4232), .O(n12695));
  LUT5 #(.INIT(32'h96696996)) lut_n12696 (.I0(x4221), .I1(x4222), .I2(x4223), .I3(n12688), .I4(n12689), .O(n12696));
  LUT5 #(.INIT(32'hFF969600)) lut_n12697 (.I0(x4227), .I1(x4228), .I2(x4229), .I3(n12695), .I4(n12696), .O(n12697));
  LUT3 #(.INIT(8'h96)) lut_n12698 (.I0(x4236), .I1(x4237), .I2(x4238), .O(n12698));
  LUT5 #(.INIT(32'h96696996)) lut_n12699 (.I0(x4227), .I1(x4228), .I2(x4229), .I3(n12695), .I4(n12696), .O(n12699));
  LUT5 #(.INIT(32'hFF969600)) lut_n12700 (.I0(x4233), .I1(x4234), .I2(x4235), .I3(n12698), .I4(n12699), .O(n12700));
  LUT3 #(.INIT(8'h96)) lut_n12701 (.I0(n12687), .I1(n12690), .I2(n12691), .O(n12701));
  LUT3 #(.INIT(8'hE8)) lut_n12702 (.I0(n12697), .I1(n12700), .I2(n12701), .O(n12702));
  LUT3 #(.INIT(8'h96)) lut_n12703 (.I0(x4242), .I1(x4243), .I2(x4244), .O(n12703));
  LUT5 #(.INIT(32'h96696996)) lut_n12704 (.I0(x4233), .I1(x4234), .I2(x4235), .I3(n12698), .I4(n12699), .O(n12704));
  LUT5 #(.INIT(32'hFF969600)) lut_n12705 (.I0(x4239), .I1(x4240), .I2(x4241), .I3(n12703), .I4(n12704), .O(n12705));
  LUT3 #(.INIT(8'h96)) lut_n12706 (.I0(x4248), .I1(x4249), .I2(x4250), .O(n12706));
  LUT5 #(.INIT(32'h96696996)) lut_n12707 (.I0(x4239), .I1(x4240), .I2(x4241), .I3(n12703), .I4(n12704), .O(n12707));
  LUT5 #(.INIT(32'hFF969600)) lut_n12708 (.I0(x4245), .I1(x4246), .I2(x4247), .I3(n12706), .I4(n12707), .O(n12708));
  LUT3 #(.INIT(8'h96)) lut_n12709 (.I0(n12697), .I1(n12700), .I2(n12701), .O(n12709));
  LUT3 #(.INIT(8'hE8)) lut_n12710 (.I0(n12705), .I1(n12708), .I2(n12709), .O(n12710));
  LUT3 #(.INIT(8'h96)) lut_n12711 (.I0(n12684), .I1(n12692), .I2(n12693), .O(n12711));
  LUT3 #(.INIT(8'hE8)) lut_n12712 (.I0(n12702), .I1(n12710), .I2(n12711), .O(n12712));
  LUT3 #(.INIT(8'h96)) lut_n12713 (.I0(n12656), .I1(n12674), .I2(n12675), .O(n12713));
  LUT3 #(.INIT(8'hE8)) lut_n12714 (.I0(n12694), .I1(n12712), .I2(n12713), .O(n12714));
  LUT3 #(.INIT(8'h96)) lut_n12715 (.I0(n12594), .I1(n12632), .I2(n12633), .O(n12715));
  LUT3 #(.INIT(8'hE8)) lut_n12716 (.I0(n12676), .I1(n12714), .I2(n12715), .O(n12716));
  LUT3 #(.INIT(8'h96)) lut_n12717 (.I0(x4254), .I1(x4255), .I2(x4256), .O(n12717));
  LUT5 #(.INIT(32'h96696996)) lut_n12718 (.I0(x4245), .I1(x4246), .I2(x4247), .I3(n12706), .I4(n12707), .O(n12718));
  LUT5 #(.INIT(32'hFF969600)) lut_n12719 (.I0(x4251), .I1(x4252), .I2(x4253), .I3(n12717), .I4(n12718), .O(n12719));
  LUT3 #(.INIT(8'h96)) lut_n12720 (.I0(x4260), .I1(x4261), .I2(x4262), .O(n12720));
  LUT5 #(.INIT(32'h96696996)) lut_n12721 (.I0(x4251), .I1(x4252), .I2(x4253), .I3(n12717), .I4(n12718), .O(n12721));
  LUT5 #(.INIT(32'hFF969600)) lut_n12722 (.I0(x4257), .I1(x4258), .I2(x4259), .I3(n12720), .I4(n12721), .O(n12722));
  LUT3 #(.INIT(8'h96)) lut_n12723 (.I0(n12705), .I1(n12708), .I2(n12709), .O(n12723));
  LUT3 #(.INIT(8'hE8)) lut_n12724 (.I0(n12719), .I1(n12722), .I2(n12723), .O(n12724));
  LUT3 #(.INIT(8'h96)) lut_n12725 (.I0(x4266), .I1(x4267), .I2(x4268), .O(n12725));
  LUT5 #(.INIT(32'h96696996)) lut_n12726 (.I0(x4257), .I1(x4258), .I2(x4259), .I3(n12720), .I4(n12721), .O(n12726));
  LUT5 #(.INIT(32'hFF969600)) lut_n12727 (.I0(x4263), .I1(x4264), .I2(x4265), .I3(n12725), .I4(n12726), .O(n12727));
  LUT3 #(.INIT(8'h96)) lut_n12728 (.I0(x4272), .I1(x4273), .I2(x4274), .O(n12728));
  LUT5 #(.INIT(32'h96696996)) lut_n12729 (.I0(x4263), .I1(x4264), .I2(x4265), .I3(n12725), .I4(n12726), .O(n12729));
  LUT5 #(.INIT(32'hFF969600)) lut_n12730 (.I0(x4269), .I1(x4270), .I2(x4271), .I3(n12728), .I4(n12729), .O(n12730));
  LUT3 #(.INIT(8'h96)) lut_n12731 (.I0(n12719), .I1(n12722), .I2(n12723), .O(n12731));
  LUT3 #(.INIT(8'hE8)) lut_n12732 (.I0(n12727), .I1(n12730), .I2(n12731), .O(n12732));
  LUT3 #(.INIT(8'h96)) lut_n12733 (.I0(n12702), .I1(n12710), .I2(n12711), .O(n12733));
  LUT3 #(.INIT(8'hE8)) lut_n12734 (.I0(n12724), .I1(n12732), .I2(n12733), .O(n12734));
  LUT3 #(.INIT(8'h96)) lut_n12735 (.I0(x4278), .I1(x4279), .I2(x4280), .O(n12735));
  LUT5 #(.INIT(32'h96696996)) lut_n12736 (.I0(x4269), .I1(x4270), .I2(x4271), .I3(n12728), .I4(n12729), .O(n12736));
  LUT5 #(.INIT(32'hFF969600)) lut_n12737 (.I0(x4275), .I1(x4276), .I2(x4277), .I3(n12735), .I4(n12736), .O(n12737));
  LUT3 #(.INIT(8'h96)) lut_n12738 (.I0(x4284), .I1(x4285), .I2(x4286), .O(n12738));
  LUT5 #(.INIT(32'h96696996)) lut_n12739 (.I0(x4275), .I1(x4276), .I2(x4277), .I3(n12735), .I4(n12736), .O(n12739));
  LUT5 #(.INIT(32'hFF969600)) lut_n12740 (.I0(x4281), .I1(x4282), .I2(x4283), .I3(n12738), .I4(n12739), .O(n12740));
  LUT3 #(.INIT(8'h96)) lut_n12741 (.I0(n12727), .I1(n12730), .I2(n12731), .O(n12741));
  LUT3 #(.INIT(8'hE8)) lut_n12742 (.I0(n12737), .I1(n12740), .I2(n12741), .O(n12742));
  LUT3 #(.INIT(8'h96)) lut_n12743 (.I0(x4290), .I1(x4291), .I2(x4292), .O(n12743));
  LUT5 #(.INIT(32'h96696996)) lut_n12744 (.I0(x4281), .I1(x4282), .I2(x4283), .I3(n12738), .I4(n12739), .O(n12744));
  LUT5 #(.INIT(32'hFF969600)) lut_n12745 (.I0(x4287), .I1(x4288), .I2(x4289), .I3(n12743), .I4(n12744), .O(n12745));
  LUT3 #(.INIT(8'h96)) lut_n12746 (.I0(x4296), .I1(x4297), .I2(x4298), .O(n12746));
  LUT5 #(.INIT(32'h96696996)) lut_n12747 (.I0(x4287), .I1(x4288), .I2(x4289), .I3(n12743), .I4(n12744), .O(n12747));
  LUT5 #(.INIT(32'hFF969600)) lut_n12748 (.I0(x4293), .I1(x4294), .I2(x4295), .I3(n12746), .I4(n12747), .O(n12748));
  LUT3 #(.INIT(8'h96)) lut_n12749 (.I0(n12737), .I1(n12740), .I2(n12741), .O(n12749));
  LUT3 #(.INIT(8'hE8)) lut_n12750 (.I0(n12745), .I1(n12748), .I2(n12749), .O(n12750));
  LUT3 #(.INIT(8'h96)) lut_n12751 (.I0(n12724), .I1(n12732), .I2(n12733), .O(n12751));
  LUT3 #(.INIT(8'hE8)) lut_n12752 (.I0(n12742), .I1(n12750), .I2(n12751), .O(n12752));
  LUT3 #(.INIT(8'h96)) lut_n12753 (.I0(n12694), .I1(n12712), .I2(n12713), .O(n12753));
  LUT3 #(.INIT(8'hE8)) lut_n12754 (.I0(n12734), .I1(n12752), .I2(n12753), .O(n12754));
  LUT3 #(.INIT(8'h96)) lut_n12755 (.I0(x4302), .I1(x4303), .I2(x4304), .O(n12755));
  LUT5 #(.INIT(32'h96696996)) lut_n12756 (.I0(x4293), .I1(x4294), .I2(x4295), .I3(n12746), .I4(n12747), .O(n12756));
  LUT5 #(.INIT(32'hFF969600)) lut_n12757 (.I0(x4299), .I1(x4300), .I2(x4301), .I3(n12755), .I4(n12756), .O(n12757));
  LUT3 #(.INIT(8'h96)) lut_n12758 (.I0(x4308), .I1(x4309), .I2(x4310), .O(n12758));
  LUT5 #(.INIT(32'h96696996)) lut_n12759 (.I0(x4299), .I1(x4300), .I2(x4301), .I3(n12755), .I4(n12756), .O(n12759));
  LUT5 #(.INIT(32'hFF969600)) lut_n12760 (.I0(x4305), .I1(x4306), .I2(x4307), .I3(n12758), .I4(n12759), .O(n12760));
  LUT3 #(.INIT(8'h96)) lut_n12761 (.I0(n12745), .I1(n12748), .I2(n12749), .O(n12761));
  LUT3 #(.INIT(8'hE8)) lut_n12762 (.I0(n12757), .I1(n12760), .I2(n12761), .O(n12762));
  LUT3 #(.INIT(8'h96)) lut_n12763 (.I0(x4314), .I1(x4315), .I2(x4316), .O(n12763));
  LUT5 #(.INIT(32'h96696996)) lut_n12764 (.I0(x4305), .I1(x4306), .I2(x4307), .I3(n12758), .I4(n12759), .O(n12764));
  LUT5 #(.INIT(32'hFF969600)) lut_n12765 (.I0(x4311), .I1(x4312), .I2(x4313), .I3(n12763), .I4(n12764), .O(n12765));
  LUT3 #(.INIT(8'h96)) lut_n12766 (.I0(x4320), .I1(x4321), .I2(x4322), .O(n12766));
  LUT5 #(.INIT(32'h96696996)) lut_n12767 (.I0(x4311), .I1(x4312), .I2(x4313), .I3(n12763), .I4(n12764), .O(n12767));
  LUT5 #(.INIT(32'hFF969600)) lut_n12768 (.I0(x4317), .I1(x4318), .I2(x4319), .I3(n12766), .I4(n12767), .O(n12768));
  LUT3 #(.INIT(8'h96)) lut_n12769 (.I0(n12757), .I1(n12760), .I2(n12761), .O(n12769));
  LUT3 #(.INIT(8'hE8)) lut_n12770 (.I0(n12765), .I1(n12768), .I2(n12769), .O(n12770));
  LUT3 #(.INIT(8'h96)) lut_n12771 (.I0(n12742), .I1(n12750), .I2(n12751), .O(n12771));
  LUT3 #(.INIT(8'hE8)) lut_n12772 (.I0(n12762), .I1(n12770), .I2(n12771), .O(n12772));
  LUT3 #(.INIT(8'h96)) lut_n12773 (.I0(x4326), .I1(x4327), .I2(x4328), .O(n12773));
  LUT5 #(.INIT(32'h96696996)) lut_n12774 (.I0(x4317), .I1(x4318), .I2(x4319), .I3(n12766), .I4(n12767), .O(n12774));
  LUT5 #(.INIT(32'hFF969600)) lut_n12775 (.I0(x4323), .I1(x4324), .I2(x4325), .I3(n12773), .I4(n12774), .O(n12775));
  LUT3 #(.INIT(8'h96)) lut_n12776 (.I0(x4332), .I1(x4333), .I2(x4334), .O(n12776));
  LUT5 #(.INIT(32'h96696996)) lut_n12777 (.I0(x4323), .I1(x4324), .I2(x4325), .I3(n12773), .I4(n12774), .O(n12777));
  LUT5 #(.INIT(32'hFF969600)) lut_n12778 (.I0(x4329), .I1(x4330), .I2(x4331), .I3(n12776), .I4(n12777), .O(n12778));
  LUT3 #(.INIT(8'h96)) lut_n12779 (.I0(n12765), .I1(n12768), .I2(n12769), .O(n12779));
  LUT3 #(.INIT(8'hE8)) lut_n12780 (.I0(n12775), .I1(n12778), .I2(n12779), .O(n12780));
  LUT3 #(.INIT(8'h96)) lut_n12781 (.I0(x4338), .I1(x4339), .I2(x4340), .O(n12781));
  LUT5 #(.INIT(32'h96696996)) lut_n12782 (.I0(x4329), .I1(x4330), .I2(x4331), .I3(n12776), .I4(n12777), .O(n12782));
  LUT5 #(.INIT(32'hFF969600)) lut_n12783 (.I0(x4335), .I1(x4336), .I2(x4337), .I3(n12781), .I4(n12782), .O(n12783));
  LUT3 #(.INIT(8'h96)) lut_n12784 (.I0(x4344), .I1(x4345), .I2(x4346), .O(n12784));
  LUT5 #(.INIT(32'h96696996)) lut_n12785 (.I0(x4335), .I1(x4336), .I2(x4337), .I3(n12781), .I4(n12782), .O(n12785));
  LUT5 #(.INIT(32'hFF969600)) lut_n12786 (.I0(x4341), .I1(x4342), .I2(x4343), .I3(n12784), .I4(n12785), .O(n12786));
  LUT3 #(.INIT(8'h96)) lut_n12787 (.I0(n12775), .I1(n12778), .I2(n12779), .O(n12787));
  LUT3 #(.INIT(8'hE8)) lut_n12788 (.I0(n12783), .I1(n12786), .I2(n12787), .O(n12788));
  LUT3 #(.INIT(8'h96)) lut_n12789 (.I0(n12762), .I1(n12770), .I2(n12771), .O(n12789));
  LUT3 #(.INIT(8'hE8)) lut_n12790 (.I0(n12780), .I1(n12788), .I2(n12789), .O(n12790));
  LUT3 #(.INIT(8'h96)) lut_n12791 (.I0(n12734), .I1(n12752), .I2(n12753), .O(n12791));
  LUT3 #(.INIT(8'hE8)) lut_n12792 (.I0(n12772), .I1(n12790), .I2(n12791), .O(n12792));
  LUT3 #(.INIT(8'h96)) lut_n12793 (.I0(n12676), .I1(n12714), .I2(n12715), .O(n12793));
  LUT3 #(.INIT(8'hE8)) lut_n12794 (.I0(n12754), .I1(n12792), .I2(n12793), .O(n12794));
  LUT3 #(.INIT(8'h96)) lut_n12795 (.I0(n12556), .I1(n12634), .I2(n12635), .O(n12795));
  LUT3 #(.INIT(8'hE8)) lut_n12796 (.I0(n12716), .I1(n12794), .I2(n12795), .O(n12796));
  LUT3 #(.INIT(8'h96)) lut_n12797 (.I0(x4350), .I1(x4351), .I2(x4352), .O(n12797));
  LUT5 #(.INIT(32'h96696996)) lut_n12798 (.I0(x4341), .I1(x4342), .I2(x4343), .I3(n12784), .I4(n12785), .O(n12798));
  LUT5 #(.INIT(32'hFF969600)) lut_n12799 (.I0(x4347), .I1(x4348), .I2(x4349), .I3(n12797), .I4(n12798), .O(n12799));
  LUT3 #(.INIT(8'h96)) lut_n12800 (.I0(x4356), .I1(x4357), .I2(x4358), .O(n12800));
  LUT5 #(.INIT(32'h96696996)) lut_n12801 (.I0(x4347), .I1(x4348), .I2(x4349), .I3(n12797), .I4(n12798), .O(n12801));
  LUT5 #(.INIT(32'hFF969600)) lut_n12802 (.I0(x4353), .I1(x4354), .I2(x4355), .I3(n12800), .I4(n12801), .O(n12802));
  LUT3 #(.INIT(8'h96)) lut_n12803 (.I0(n12783), .I1(n12786), .I2(n12787), .O(n12803));
  LUT3 #(.INIT(8'hE8)) lut_n12804 (.I0(n12799), .I1(n12802), .I2(n12803), .O(n12804));
  LUT3 #(.INIT(8'h96)) lut_n12805 (.I0(x4362), .I1(x4363), .I2(x4364), .O(n12805));
  LUT5 #(.INIT(32'h96696996)) lut_n12806 (.I0(x4353), .I1(x4354), .I2(x4355), .I3(n12800), .I4(n12801), .O(n12806));
  LUT5 #(.INIT(32'hFF969600)) lut_n12807 (.I0(x4359), .I1(x4360), .I2(x4361), .I3(n12805), .I4(n12806), .O(n12807));
  LUT3 #(.INIT(8'h96)) lut_n12808 (.I0(x4368), .I1(x4369), .I2(x4370), .O(n12808));
  LUT5 #(.INIT(32'h96696996)) lut_n12809 (.I0(x4359), .I1(x4360), .I2(x4361), .I3(n12805), .I4(n12806), .O(n12809));
  LUT5 #(.INIT(32'hFF969600)) lut_n12810 (.I0(x4365), .I1(x4366), .I2(x4367), .I3(n12808), .I4(n12809), .O(n12810));
  LUT3 #(.INIT(8'h96)) lut_n12811 (.I0(n12799), .I1(n12802), .I2(n12803), .O(n12811));
  LUT3 #(.INIT(8'hE8)) lut_n12812 (.I0(n12807), .I1(n12810), .I2(n12811), .O(n12812));
  LUT3 #(.INIT(8'h96)) lut_n12813 (.I0(n12780), .I1(n12788), .I2(n12789), .O(n12813));
  LUT3 #(.INIT(8'hE8)) lut_n12814 (.I0(n12804), .I1(n12812), .I2(n12813), .O(n12814));
  LUT3 #(.INIT(8'h96)) lut_n12815 (.I0(x4374), .I1(x4375), .I2(x4376), .O(n12815));
  LUT5 #(.INIT(32'h96696996)) lut_n12816 (.I0(x4365), .I1(x4366), .I2(x4367), .I3(n12808), .I4(n12809), .O(n12816));
  LUT5 #(.INIT(32'hFF969600)) lut_n12817 (.I0(x4371), .I1(x4372), .I2(x4373), .I3(n12815), .I4(n12816), .O(n12817));
  LUT3 #(.INIT(8'h96)) lut_n12818 (.I0(x4380), .I1(x4381), .I2(x4382), .O(n12818));
  LUT5 #(.INIT(32'h96696996)) lut_n12819 (.I0(x4371), .I1(x4372), .I2(x4373), .I3(n12815), .I4(n12816), .O(n12819));
  LUT5 #(.INIT(32'hFF969600)) lut_n12820 (.I0(x4377), .I1(x4378), .I2(x4379), .I3(n12818), .I4(n12819), .O(n12820));
  LUT3 #(.INIT(8'h96)) lut_n12821 (.I0(n12807), .I1(n12810), .I2(n12811), .O(n12821));
  LUT3 #(.INIT(8'hE8)) lut_n12822 (.I0(n12817), .I1(n12820), .I2(n12821), .O(n12822));
  LUT3 #(.INIT(8'h96)) lut_n12823 (.I0(x4386), .I1(x4387), .I2(x4388), .O(n12823));
  LUT5 #(.INIT(32'h96696996)) lut_n12824 (.I0(x4377), .I1(x4378), .I2(x4379), .I3(n12818), .I4(n12819), .O(n12824));
  LUT5 #(.INIT(32'hFF969600)) lut_n12825 (.I0(x4383), .I1(x4384), .I2(x4385), .I3(n12823), .I4(n12824), .O(n12825));
  LUT3 #(.INIT(8'h96)) lut_n12826 (.I0(x4392), .I1(x4393), .I2(x4394), .O(n12826));
  LUT5 #(.INIT(32'h96696996)) lut_n12827 (.I0(x4383), .I1(x4384), .I2(x4385), .I3(n12823), .I4(n12824), .O(n12827));
  LUT5 #(.INIT(32'hFF969600)) lut_n12828 (.I0(x4389), .I1(x4390), .I2(x4391), .I3(n12826), .I4(n12827), .O(n12828));
  LUT3 #(.INIT(8'h96)) lut_n12829 (.I0(n12817), .I1(n12820), .I2(n12821), .O(n12829));
  LUT3 #(.INIT(8'hE8)) lut_n12830 (.I0(n12825), .I1(n12828), .I2(n12829), .O(n12830));
  LUT3 #(.INIT(8'h96)) lut_n12831 (.I0(n12804), .I1(n12812), .I2(n12813), .O(n12831));
  LUT3 #(.INIT(8'hE8)) lut_n12832 (.I0(n12822), .I1(n12830), .I2(n12831), .O(n12832));
  LUT3 #(.INIT(8'h96)) lut_n12833 (.I0(n12772), .I1(n12790), .I2(n12791), .O(n12833));
  LUT3 #(.INIT(8'hE8)) lut_n12834 (.I0(n12814), .I1(n12832), .I2(n12833), .O(n12834));
  LUT3 #(.INIT(8'h96)) lut_n12835 (.I0(x4398), .I1(x4399), .I2(x4400), .O(n12835));
  LUT5 #(.INIT(32'h96696996)) lut_n12836 (.I0(x4389), .I1(x4390), .I2(x4391), .I3(n12826), .I4(n12827), .O(n12836));
  LUT5 #(.INIT(32'hFF969600)) lut_n12837 (.I0(x4395), .I1(x4396), .I2(x4397), .I3(n12835), .I4(n12836), .O(n12837));
  LUT3 #(.INIT(8'h96)) lut_n12838 (.I0(x4404), .I1(x4405), .I2(x4406), .O(n12838));
  LUT5 #(.INIT(32'h96696996)) lut_n12839 (.I0(x4395), .I1(x4396), .I2(x4397), .I3(n12835), .I4(n12836), .O(n12839));
  LUT5 #(.INIT(32'hFF969600)) lut_n12840 (.I0(x4401), .I1(x4402), .I2(x4403), .I3(n12838), .I4(n12839), .O(n12840));
  LUT3 #(.INIT(8'h96)) lut_n12841 (.I0(n12825), .I1(n12828), .I2(n12829), .O(n12841));
  LUT3 #(.INIT(8'hE8)) lut_n12842 (.I0(n12837), .I1(n12840), .I2(n12841), .O(n12842));
  LUT3 #(.INIT(8'h96)) lut_n12843 (.I0(x4410), .I1(x4411), .I2(x4412), .O(n12843));
  LUT5 #(.INIT(32'h96696996)) lut_n12844 (.I0(x4401), .I1(x4402), .I2(x4403), .I3(n12838), .I4(n12839), .O(n12844));
  LUT5 #(.INIT(32'hFF969600)) lut_n12845 (.I0(x4407), .I1(x4408), .I2(x4409), .I3(n12843), .I4(n12844), .O(n12845));
  LUT3 #(.INIT(8'h96)) lut_n12846 (.I0(x4416), .I1(x4417), .I2(x4418), .O(n12846));
  LUT5 #(.INIT(32'h96696996)) lut_n12847 (.I0(x4407), .I1(x4408), .I2(x4409), .I3(n12843), .I4(n12844), .O(n12847));
  LUT5 #(.INIT(32'hFF969600)) lut_n12848 (.I0(x4413), .I1(x4414), .I2(x4415), .I3(n12846), .I4(n12847), .O(n12848));
  LUT3 #(.INIT(8'h96)) lut_n12849 (.I0(n12837), .I1(n12840), .I2(n12841), .O(n12849));
  LUT3 #(.INIT(8'hE8)) lut_n12850 (.I0(n12845), .I1(n12848), .I2(n12849), .O(n12850));
  LUT3 #(.INIT(8'h96)) lut_n12851 (.I0(n12822), .I1(n12830), .I2(n12831), .O(n12851));
  LUT3 #(.INIT(8'hE8)) lut_n12852 (.I0(n12842), .I1(n12850), .I2(n12851), .O(n12852));
  LUT3 #(.INIT(8'h96)) lut_n12853 (.I0(x4422), .I1(x4423), .I2(x4424), .O(n12853));
  LUT5 #(.INIT(32'h96696996)) lut_n12854 (.I0(x4413), .I1(x4414), .I2(x4415), .I3(n12846), .I4(n12847), .O(n12854));
  LUT5 #(.INIT(32'hFF969600)) lut_n12855 (.I0(x4419), .I1(x4420), .I2(x4421), .I3(n12853), .I4(n12854), .O(n12855));
  LUT3 #(.INIT(8'h96)) lut_n12856 (.I0(x4428), .I1(x4429), .I2(x4430), .O(n12856));
  LUT5 #(.INIT(32'h96696996)) lut_n12857 (.I0(x4419), .I1(x4420), .I2(x4421), .I3(n12853), .I4(n12854), .O(n12857));
  LUT5 #(.INIT(32'hFF969600)) lut_n12858 (.I0(x4425), .I1(x4426), .I2(x4427), .I3(n12856), .I4(n12857), .O(n12858));
  LUT3 #(.INIT(8'h96)) lut_n12859 (.I0(n12845), .I1(n12848), .I2(n12849), .O(n12859));
  LUT3 #(.INIT(8'hE8)) lut_n12860 (.I0(n12855), .I1(n12858), .I2(n12859), .O(n12860));
  LUT3 #(.INIT(8'h96)) lut_n12861 (.I0(x4434), .I1(x4435), .I2(x4436), .O(n12861));
  LUT5 #(.INIT(32'h96696996)) lut_n12862 (.I0(x4425), .I1(x4426), .I2(x4427), .I3(n12856), .I4(n12857), .O(n12862));
  LUT5 #(.INIT(32'hFF969600)) lut_n12863 (.I0(x4431), .I1(x4432), .I2(x4433), .I3(n12861), .I4(n12862), .O(n12863));
  LUT3 #(.INIT(8'h96)) lut_n12864 (.I0(x4440), .I1(x4441), .I2(x4442), .O(n12864));
  LUT5 #(.INIT(32'h96696996)) lut_n12865 (.I0(x4431), .I1(x4432), .I2(x4433), .I3(n12861), .I4(n12862), .O(n12865));
  LUT5 #(.INIT(32'hFF969600)) lut_n12866 (.I0(x4437), .I1(x4438), .I2(x4439), .I3(n12864), .I4(n12865), .O(n12866));
  LUT3 #(.INIT(8'h96)) lut_n12867 (.I0(n12855), .I1(n12858), .I2(n12859), .O(n12867));
  LUT3 #(.INIT(8'hE8)) lut_n12868 (.I0(n12863), .I1(n12866), .I2(n12867), .O(n12868));
  LUT3 #(.INIT(8'h96)) lut_n12869 (.I0(n12842), .I1(n12850), .I2(n12851), .O(n12869));
  LUT3 #(.INIT(8'hE8)) lut_n12870 (.I0(n12860), .I1(n12868), .I2(n12869), .O(n12870));
  LUT3 #(.INIT(8'h96)) lut_n12871 (.I0(n12814), .I1(n12832), .I2(n12833), .O(n12871));
  LUT3 #(.INIT(8'hE8)) lut_n12872 (.I0(n12852), .I1(n12870), .I2(n12871), .O(n12872));
  LUT3 #(.INIT(8'h96)) lut_n12873 (.I0(n12754), .I1(n12792), .I2(n12793), .O(n12873));
  LUT3 #(.INIT(8'hE8)) lut_n12874 (.I0(n12834), .I1(n12872), .I2(n12873), .O(n12874));
  LUT3 #(.INIT(8'h96)) lut_n12875 (.I0(x4446), .I1(x4447), .I2(x4448), .O(n12875));
  LUT5 #(.INIT(32'h96696996)) lut_n12876 (.I0(x4437), .I1(x4438), .I2(x4439), .I3(n12864), .I4(n12865), .O(n12876));
  LUT5 #(.INIT(32'hFF969600)) lut_n12877 (.I0(x4443), .I1(x4444), .I2(x4445), .I3(n12875), .I4(n12876), .O(n12877));
  LUT3 #(.INIT(8'h96)) lut_n12878 (.I0(x4452), .I1(x4453), .I2(x4454), .O(n12878));
  LUT5 #(.INIT(32'h96696996)) lut_n12879 (.I0(x4443), .I1(x4444), .I2(x4445), .I3(n12875), .I4(n12876), .O(n12879));
  LUT5 #(.INIT(32'hFF969600)) lut_n12880 (.I0(x4449), .I1(x4450), .I2(x4451), .I3(n12878), .I4(n12879), .O(n12880));
  LUT3 #(.INIT(8'h96)) lut_n12881 (.I0(n12863), .I1(n12866), .I2(n12867), .O(n12881));
  LUT3 #(.INIT(8'hE8)) lut_n12882 (.I0(n12877), .I1(n12880), .I2(n12881), .O(n12882));
  LUT3 #(.INIT(8'h96)) lut_n12883 (.I0(x4458), .I1(x4459), .I2(x4460), .O(n12883));
  LUT5 #(.INIT(32'h96696996)) lut_n12884 (.I0(x4449), .I1(x4450), .I2(x4451), .I3(n12878), .I4(n12879), .O(n12884));
  LUT5 #(.INIT(32'hFF969600)) lut_n12885 (.I0(x4455), .I1(x4456), .I2(x4457), .I3(n12883), .I4(n12884), .O(n12885));
  LUT3 #(.INIT(8'h96)) lut_n12886 (.I0(x4464), .I1(x4465), .I2(x4466), .O(n12886));
  LUT5 #(.INIT(32'h96696996)) lut_n12887 (.I0(x4455), .I1(x4456), .I2(x4457), .I3(n12883), .I4(n12884), .O(n12887));
  LUT5 #(.INIT(32'hFF969600)) lut_n12888 (.I0(x4461), .I1(x4462), .I2(x4463), .I3(n12886), .I4(n12887), .O(n12888));
  LUT3 #(.INIT(8'h96)) lut_n12889 (.I0(n12877), .I1(n12880), .I2(n12881), .O(n12889));
  LUT3 #(.INIT(8'hE8)) lut_n12890 (.I0(n12885), .I1(n12888), .I2(n12889), .O(n12890));
  LUT3 #(.INIT(8'h96)) lut_n12891 (.I0(n12860), .I1(n12868), .I2(n12869), .O(n12891));
  LUT3 #(.INIT(8'hE8)) lut_n12892 (.I0(n12882), .I1(n12890), .I2(n12891), .O(n12892));
  LUT3 #(.INIT(8'h96)) lut_n12893 (.I0(x4470), .I1(x4471), .I2(x4472), .O(n12893));
  LUT5 #(.INIT(32'h96696996)) lut_n12894 (.I0(x4461), .I1(x4462), .I2(x4463), .I3(n12886), .I4(n12887), .O(n12894));
  LUT5 #(.INIT(32'hFF969600)) lut_n12895 (.I0(x4467), .I1(x4468), .I2(x4469), .I3(n12893), .I4(n12894), .O(n12895));
  LUT3 #(.INIT(8'h96)) lut_n12896 (.I0(x4476), .I1(x4477), .I2(x4478), .O(n12896));
  LUT5 #(.INIT(32'h96696996)) lut_n12897 (.I0(x4467), .I1(x4468), .I2(x4469), .I3(n12893), .I4(n12894), .O(n12897));
  LUT5 #(.INIT(32'hFF969600)) lut_n12898 (.I0(x4473), .I1(x4474), .I2(x4475), .I3(n12896), .I4(n12897), .O(n12898));
  LUT3 #(.INIT(8'h96)) lut_n12899 (.I0(n12885), .I1(n12888), .I2(n12889), .O(n12899));
  LUT3 #(.INIT(8'hE8)) lut_n12900 (.I0(n12895), .I1(n12898), .I2(n12899), .O(n12900));
  LUT3 #(.INIT(8'h96)) lut_n12901 (.I0(x4482), .I1(x4483), .I2(x4484), .O(n12901));
  LUT5 #(.INIT(32'h96696996)) lut_n12902 (.I0(x4473), .I1(x4474), .I2(x4475), .I3(n12896), .I4(n12897), .O(n12902));
  LUT5 #(.INIT(32'hFF969600)) lut_n12903 (.I0(x4479), .I1(x4480), .I2(x4481), .I3(n12901), .I4(n12902), .O(n12903));
  LUT3 #(.INIT(8'h96)) lut_n12904 (.I0(x4488), .I1(x4489), .I2(x4490), .O(n12904));
  LUT5 #(.INIT(32'h96696996)) lut_n12905 (.I0(x4479), .I1(x4480), .I2(x4481), .I3(n12901), .I4(n12902), .O(n12905));
  LUT5 #(.INIT(32'hFF969600)) lut_n12906 (.I0(x4485), .I1(x4486), .I2(x4487), .I3(n12904), .I4(n12905), .O(n12906));
  LUT3 #(.INIT(8'h96)) lut_n12907 (.I0(n12895), .I1(n12898), .I2(n12899), .O(n12907));
  LUT3 #(.INIT(8'hE8)) lut_n12908 (.I0(n12903), .I1(n12906), .I2(n12907), .O(n12908));
  LUT3 #(.INIT(8'h96)) lut_n12909 (.I0(n12882), .I1(n12890), .I2(n12891), .O(n12909));
  LUT3 #(.INIT(8'hE8)) lut_n12910 (.I0(n12900), .I1(n12908), .I2(n12909), .O(n12910));
  LUT3 #(.INIT(8'h96)) lut_n12911 (.I0(n12852), .I1(n12870), .I2(n12871), .O(n12911));
  LUT3 #(.INIT(8'hE8)) lut_n12912 (.I0(n12892), .I1(n12910), .I2(n12911), .O(n12912));
  LUT3 #(.INIT(8'h96)) lut_n12913 (.I0(x4494), .I1(x4495), .I2(x4496), .O(n12913));
  LUT5 #(.INIT(32'h96696996)) lut_n12914 (.I0(x4485), .I1(x4486), .I2(x4487), .I3(n12904), .I4(n12905), .O(n12914));
  LUT5 #(.INIT(32'hFF969600)) lut_n12915 (.I0(x4491), .I1(x4492), .I2(x4493), .I3(n12913), .I4(n12914), .O(n12915));
  LUT3 #(.INIT(8'h96)) lut_n12916 (.I0(x4500), .I1(x4501), .I2(x4502), .O(n12916));
  LUT5 #(.INIT(32'h96696996)) lut_n12917 (.I0(x4491), .I1(x4492), .I2(x4493), .I3(n12913), .I4(n12914), .O(n12917));
  LUT5 #(.INIT(32'hFF969600)) lut_n12918 (.I0(x4497), .I1(x4498), .I2(x4499), .I3(n12916), .I4(n12917), .O(n12918));
  LUT3 #(.INIT(8'h96)) lut_n12919 (.I0(n12903), .I1(n12906), .I2(n12907), .O(n12919));
  LUT3 #(.INIT(8'hE8)) lut_n12920 (.I0(n12915), .I1(n12918), .I2(n12919), .O(n12920));
  LUT3 #(.INIT(8'h96)) lut_n12921 (.I0(x4506), .I1(x4507), .I2(x4508), .O(n12921));
  LUT5 #(.INIT(32'h96696996)) lut_n12922 (.I0(x4497), .I1(x4498), .I2(x4499), .I3(n12916), .I4(n12917), .O(n12922));
  LUT5 #(.INIT(32'hFF969600)) lut_n12923 (.I0(x4503), .I1(x4504), .I2(x4505), .I3(n12921), .I4(n12922), .O(n12923));
  LUT3 #(.INIT(8'h96)) lut_n12924 (.I0(x4512), .I1(x4513), .I2(x4514), .O(n12924));
  LUT5 #(.INIT(32'h96696996)) lut_n12925 (.I0(x4503), .I1(x4504), .I2(x4505), .I3(n12921), .I4(n12922), .O(n12925));
  LUT5 #(.INIT(32'hFF969600)) lut_n12926 (.I0(x4509), .I1(x4510), .I2(x4511), .I3(n12924), .I4(n12925), .O(n12926));
  LUT3 #(.INIT(8'h96)) lut_n12927 (.I0(n12915), .I1(n12918), .I2(n12919), .O(n12927));
  LUT3 #(.INIT(8'hE8)) lut_n12928 (.I0(n12923), .I1(n12926), .I2(n12927), .O(n12928));
  LUT3 #(.INIT(8'h96)) lut_n12929 (.I0(n12900), .I1(n12908), .I2(n12909), .O(n12929));
  LUT3 #(.INIT(8'hE8)) lut_n12930 (.I0(n12920), .I1(n12928), .I2(n12929), .O(n12930));
  LUT3 #(.INIT(8'h96)) lut_n12931 (.I0(x4518), .I1(x4519), .I2(x4520), .O(n12931));
  LUT5 #(.INIT(32'h96696996)) lut_n12932 (.I0(x4509), .I1(x4510), .I2(x4511), .I3(n12924), .I4(n12925), .O(n12932));
  LUT5 #(.INIT(32'hFF969600)) lut_n12933 (.I0(x4515), .I1(x4516), .I2(x4517), .I3(n12931), .I4(n12932), .O(n12933));
  LUT3 #(.INIT(8'h96)) lut_n12934 (.I0(x4524), .I1(x4525), .I2(x4526), .O(n12934));
  LUT5 #(.INIT(32'h96696996)) lut_n12935 (.I0(x4515), .I1(x4516), .I2(x4517), .I3(n12931), .I4(n12932), .O(n12935));
  LUT5 #(.INIT(32'hFF969600)) lut_n12936 (.I0(x4521), .I1(x4522), .I2(x4523), .I3(n12934), .I4(n12935), .O(n12936));
  LUT3 #(.INIT(8'h96)) lut_n12937 (.I0(n12923), .I1(n12926), .I2(n12927), .O(n12937));
  LUT3 #(.INIT(8'hE8)) lut_n12938 (.I0(n12933), .I1(n12936), .I2(n12937), .O(n12938));
  LUT3 #(.INIT(8'h96)) lut_n12939 (.I0(x4530), .I1(x4531), .I2(x4532), .O(n12939));
  LUT5 #(.INIT(32'h96696996)) lut_n12940 (.I0(x4521), .I1(x4522), .I2(x4523), .I3(n12934), .I4(n12935), .O(n12940));
  LUT5 #(.INIT(32'hFF969600)) lut_n12941 (.I0(x4527), .I1(x4528), .I2(x4529), .I3(n12939), .I4(n12940), .O(n12941));
  LUT3 #(.INIT(8'h96)) lut_n12942 (.I0(x4536), .I1(x4537), .I2(x4538), .O(n12942));
  LUT5 #(.INIT(32'h96696996)) lut_n12943 (.I0(x4527), .I1(x4528), .I2(x4529), .I3(n12939), .I4(n12940), .O(n12943));
  LUT5 #(.INIT(32'hFF969600)) lut_n12944 (.I0(x4533), .I1(x4534), .I2(x4535), .I3(n12942), .I4(n12943), .O(n12944));
  LUT3 #(.INIT(8'h96)) lut_n12945 (.I0(n12933), .I1(n12936), .I2(n12937), .O(n12945));
  LUT3 #(.INIT(8'hE8)) lut_n12946 (.I0(n12941), .I1(n12944), .I2(n12945), .O(n12946));
  LUT3 #(.INIT(8'h96)) lut_n12947 (.I0(n12920), .I1(n12928), .I2(n12929), .O(n12947));
  LUT3 #(.INIT(8'hE8)) lut_n12948 (.I0(n12938), .I1(n12946), .I2(n12947), .O(n12948));
  LUT3 #(.INIT(8'h96)) lut_n12949 (.I0(n12892), .I1(n12910), .I2(n12911), .O(n12949));
  LUT3 #(.INIT(8'hE8)) lut_n12950 (.I0(n12930), .I1(n12948), .I2(n12949), .O(n12950));
  LUT3 #(.INIT(8'h96)) lut_n12951 (.I0(n12834), .I1(n12872), .I2(n12873), .O(n12951));
  LUT3 #(.INIT(8'hE8)) lut_n12952 (.I0(n12912), .I1(n12950), .I2(n12951), .O(n12952));
  LUT3 #(.INIT(8'h96)) lut_n12953 (.I0(n12716), .I1(n12794), .I2(n12795), .O(n12953));
  LUT3 #(.INIT(8'hE8)) lut_n12954 (.I0(n12874), .I1(n12952), .I2(n12953), .O(n12954));
  LUT3 #(.INIT(8'h96)) lut_n12955 (.I0(n12478), .I1(n12636), .I2(n12637), .O(n12955));
  LUT3 #(.INIT(8'hE8)) lut_n12956 (.I0(n12796), .I1(n12954), .I2(n12955), .O(n12956));
  LUT3 #(.INIT(8'h96)) lut_n12957 (.I0(n11998), .I1(n12316), .I2(n12317), .O(n12957));
  LUT3 #(.INIT(8'hE8)) lut_n12958 (.I0(n12638), .I1(n12956), .I2(n12957), .O(n12958));
  LUT3 #(.INIT(8'h96)) lut_n12959 (.I0(x4542), .I1(x4543), .I2(x4544), .O(n12959));
  LUT5 #(.INIT(32'h96696996)) lut_n12960 (.I0(x4533), .I1(x4534), .I2(x4535), .I3(n12942), .I4(n12943), .O(n12960));
  LUT5 #(.INIT(32'hFF969600)) lut_n12961 (.I0(x4539), .I1(x4540), .I2(x4541), .I3(n12959), .I4(n12960), .O(n12961));
  LUT3 #(.INIT(8'h96)) lut_n12962 (.I0(x4548), .I1(x4549), .I2(x4550), .O(n12962));
  LUT5 #(.INIT(32'h96696996)) lut_n12963 (.I0(x4539), .I1(x4540), .I2(x4541), .I3(n12959), .I4(n12960), .O(n12963));
  LUT5 #(.INIT(32'hFF969600)) lut_n12964 (.I0(x4545), .I1(x4546), .I2(x4547), .I3(n12962), .I4(n12963), .O(n12964));
  LUT3 #(.INIT(8'h96)) lut_n12965 (.I0(n12941), .I1(n12944), .I2(n12945), .O(n12965));
  LUT3 #(.INIT(8'hE8)) lut_n12966 (.I0(n12961), .I1(n12964), .I2(n12965), .O(n12966));
  LUT3 #(.INIT(8'h96)) lut_n12967 (.I0(x4554), .I1(x4555), .I2(x4556), .O(n12967));
  LUT5 #(.INIT(32'h96696996)) lut_n12968 (.I0(x4545), .I1(x4546), .I2(x4547), .I3(n12962), .I4(n12963), .O(n12968));
  LUT5 #(.INIT(32'hFF969600)) lut_n12969 (.I0(x4551), .I1(x4552), .I2(x4553), .I3(n12967), .I4(n12968), .O(n12969));
  LUT3 #(.INIT(8'h96)) lut_n12970 (.I0(x4560), .I1(x4561), .I2(x4562), .O(n12970));
  LUT5 #(.INIT(32'h96696996)) lut_n12971 (.I0(x4551), .I1(x4552), .I2(x4553), .I3(n12967), .I4(n12968), .O(n12971));
  LUT5 #(.INIT(32'hFF969600)) lut_n12972 (.I0(x4557), .I1(x4558), .I2(x4559), .I3(n12970), .I4(n12971), .O(n12972));
  LUT3 #(.INIT(8'h96)) lut_n12973 (.I0(n12961), .I1(n12964), .I2(n12965), .O(n12973));
  LUT3 #(.INIT(8'hE8)) lut_n12974 (.I0(n12969), .I1(n12972), .I2(n12973), .O(n12974));
  LUT3 #(.INIT(8'h96)) lut_n12975 (.I0(n12938), .I1(n12946), .I2(n12947), .O(n12975));
  LUT3 #(.INIT(8'hE8)) lut_n12976 (.I0(n12966), .I1(n12974), .I2(n12975), .O(n12976));
  LUT3 #(.INIT(8'h96)) lut_n12977 (.I0(x4566), .I1(x4567), .I2(x4568), .O(n12977));
  LUT5 #(.INIT(32'h96696996)) lut_n12978 (.I0(x4557), .I1(x4558), .I2(x4559), .I3(n12970), .I4(n12971), .O(n12978));
  LUT5 #(.INIT(32'hFF969600)) lut_n12979 (.I0(x4563), .I1(x4564), .I2(x4565), .I3(n12977), .I4(n12978), .O(n12979));
  LUT3 #(.INIT(8'h96)) lut_n12980 (.I0(x4572), .I1(x4573), .I2(x4574), .O(n12980));
  LUT5 #(.INIT(32'h96696996)) lut_n12981 (.I0(x4563), .I1(x4564), .I2(x4565), .I3(n12977), .I4(n12978), .O(n12981));
  LUT5 #(.INIT(32'hFF969600)) lut_n12982 (.I0(x4569), .I1(x4570), .I2(x4571), .I3(n12980), .I4(n12981), .O(n12982));
  LUT3 #(.INIT(8'h96)) lut_n12983 (.I0(n12969), .I1(n12972), .I2(n12973), .O(n12983));
  LUT3 #(.INIT(8'hE8)) lut_n12984 (.I0(n12979), .I1(n12982), .I2(n12983), .O(n12984));
  LUT3 #(.INIT(8'h96)) lut_n12985 (.I0(x4578), .I1(x4579), .I2(x4580), .O(n12985));
  LUT5 #(.INIT(32'h96696996)) lut_n12986 (.I0(x4569), .I1(x4570), .I2(x4571), .I3(n12980), .I4(n12981), .O(n12986));
  LUT5 #(.INIT(32'hFF969600)) lut_n12987 (.I0(x4575), .I1(x4576), .I2(x4577), .I3(n12985), .I4(n12986), .O(n12987));
  LUT3 #(.INIT(8'h96)) lut_n12988 (.I0(x4584), .I1(x4585), .I2(x4586), .O(n12988));
  LUT5 #(.INIT(32'h96696996)) lut_n12989 (.I0(x4575), .I1(x4576), .I2(x4577), .I3(n12985), .I4(n12986), .O(n12989));
  LUT5 #(.INIT(32'hFF969600)) lut_n12990 (.I0(x4581), .I1(x4582), .I2(x4583), .I3(n12988), .I4(n12989), .O(n12990));
  LUT3 #(.INIT(8'h96)) lut_n12991 (.I0(n12979), .I1(n12982), .I2(n12983), .O(n12991));
  LUT3 #(.INIT(8'hE8)) lut_n12992 (.I0(n12987), .I1(n12990), .I2(n12991), .O(n12992));
  LUT3 #(.INIT(8'h96)) lut_n12993 (.I0(n12966), .I1(n12974), .I2(n12975), .O(n12993));
  LUT3 #(.INIT(8'hE8)) lut_n12994 (.I0(n12984), .I1(n12992), .I2(n12993), .O(n12994));
  LUT3 #(.INIT(8'h96)) lut_n12995 (.I0(n12930), .I1(n12948), .I2(n12949), .O(n12995));
  LUT3 #(.INIT(8'hE8)) lut_n12996 (.I0(n12976), .I1(n12994), .I2(n12995), .O(n12996));
  LUT3 #(.INIT(8'h96)) lut_n12997 (.I0(x4590), .I1(x4591), .I2(x4592), .O(n12997));
  LUT5 #(.INIT(32'h96696996)) lut_n12998 (.I0(x4581), .I1(x4582), .I2(x4583), .I3(n12988), .I4(n12989), .O(n12998));
  LUT5 #(.INIT(32'hFF969600)) lut_n12999 (.I0(x4587), .I1(x4588), .I2(x4589), .I3(n12997), .I4(n12998), .O(n12999));
  LUT3 #(.INIT(8'h96)) lut_n13000 (.I0(x4596), .I1(x4597), .I2(x4598), .O(n13000));
  LUT5 #(.INIT(32'h96696996)) lut_n13001 (.I0(x4587), .I1(x4588), .I2(x4589), .I3(n12997), .I4(n12998), .O(n13001));
  LUT5 #(.INIT(32'hFF969600)) lut_n13002 (.I0(x4593), .I1(x4594), .I2(x4595), .I3(n13000), .I4(n13001), .O(n13002));
  LUT3 #(.INIT(8'h96)) lut_n13003 (.I0(n12987), .I1(n12990), .I2(n12991), .O(n13003));
  LUT3 #(.INIT(8'hE8)) lut_n13004 (.I0(n12999), .I1(n13002), .I2(n13003), .O(n13004));
  LUT3 #(.INIT(8'h96)) lut_n13005 (.I0(x4602), .I1(x4603), .I2(x4604), .O(n13005));
  LUT5 #(.INIT(32'h96696996)) lut_n13006 (.I0(x4593), .I1(x4594), .I2(x4595), .I3(n13000), .I4(n13001), .O(n13006));
  LUT5 #(.INIT(32'hFF969600)) lut_n13007 (.I0(x4599), .I1(x4600), .I2(x4601), .I3(n13005), .I4(n13006), .O(n13007));
  LUT3 #(.INIT(8'h96)) lut_n13008 (.I0(x4608), .I1(x4609), .I2(x4610), .O(n13008));
  LUT5 #(.INIT(32'h96696996)) lut_n13009 (.I0(x4599), .I1(x4600), .I2(x4601), .I3(n13005), .I4(n13006), .O(n13009));
  LUT5 #(.INIT(32'hFF969600)) lut_n13010 (.I0(x4605), .I1(x4606), .I2(x4607), .I3(n13008), .I4(n13009), .O(n13010));
  LUT3 #(.INIT(8'h96)) lut_n13011 (.I0(n12999), .I1(n13002), .I2(n13003), .O(n13011));
  LUT3 #(.INIT(8'hE8)) lut_n13012 (.I0(n13007), .I1(n13010), .I2(n13011), .O(n13012));
  LUT3 #(.INIT(8'h96)) lut_n13013 (.I0(n12984), .I1(n12992), .I2(n12993), .O(n13013));
  LUT3 #(.INIT(8'hE8)) lut_n13014 (.I0(n13004), .I1(n13012), .I2(n13013), .O(n13014));
  LUT3 #(.INIT(8'h96)) lut_n13015 (.I0(x4614), .I1(x4615), .I2(x4616), .O(n13015));
  LUT5 #(.INIT(32'h96696996)) lut_n13016 (.I0(x4605), .I1(x4606), .I2(x4607), .I3(n13008), .I4(n13009), .O(n13016));
  LUT5 #(.INIT(32'hFF969600)) lut_n13017 (.I0(x4611), .I1(x4612), .I2(x4613), .I3(n13015), .I4(n13016), .O(n13017));
  LUT3 #(.INIT(8'h96)) lut_n13018 (.I0(x4620), .I1(x4621), .I2(x4622), .O(n13018));
  LUT5 #(.INIT(32'h96696996)) lut_n13019 (.I0(x4611), .I1(x4612), .I2(x4613), .I3(n13015), .I4(n13016), .O(n13019));
  LUT5 #(.INIT(32'hFF969600)) lut_n13020 (.I0(x4617), .I1(x4618), .I2(x4619), .I3(n13018), .I4(n13019), .O(n13020));
  LUT3 #(.INIT(8'h96)) lut_n13021 (.I0(n13007), .I1(n13010), .I2(n13011), .O(n13021));
  LUT3 #(.INIT(8'hE8)) lut_n13022 (.I0(n13017), .I1(n13020), .I2(n13021), .O(n13022));
  LUT3 #(.INIT(8'h96)) lut_n13023 (.I0(x4626), .I1(x4627), .I2(x4628), .O(n13023));
  LUT5 #(.INIT(32'h96696996)) lut_n13024 (.I0(x4617), .I1(x4618), .I2(x4619), .I3(n13018), .I4(n13019), .O(n13024));
  LUT5 #(.INIT(32'hFF969600)) lut_n13025 (.I0(x4623), .I1(x4624), .I2(x4625), .I3(n13023), .I4(n13024), .O(n13025));
  LUT3 #(.INIT(8'h96)) lut_n13026 (.I0(x4632), .I1(x4633), .I2(x4634), .O(n13026));
  LUT5 #(.INIT(32'h96696996)) lut_n13027 (.I0(x4623), .I1(x4624), .I2(x4625), .I3(n13023), .I4(n13024), .O(n13027));
  LUT5 #(.INIT(32'hFF969600)) lut_n13028 (.I0(x4629), .I1(x4630), .I2(x4631), .I3(n13026), .I4(n13027), .O(n13028));
  LUT3 #(.INIT(8'h96)) lut_n13029 (.I0(n13017), .I1(n13020), .I2(n13021), .O(n13029));
  LUT3 #(.INIT(8'hE8)) lut_n13030 (.I0(n13025), .I1(n13028), .I2(n13029), .O(n13030));
  LUT3 #(.INIT(8'h96)) lut_n13031 (.I0(n13004), .I1(n13012), .I2(n13013), .O(n13031));
  LUT3 #(.INIT(8'hE8)) lut_n13032 (.I0(n13022), .I1(n13030), .I2(n13031), .O(n13032));
  LUT3 #(.INIT(8'h96)) lut_n13033 (.I0(n12976), .I1(n12994), .I2(n12995), .O(n13033));
  LUT3 #(.INIT(8'hE8)) lut_n13034 (.I0(n13014), .I1(n13032), .I2(n13033), .O(n13034));
  LUT3 #(.INIT(8'h96)) lut_n13035 (.I0(n12912), .I1(n12950), .I2(n12951), .O(n13035));
  LUT3 #(.INIT(8'hE8)) lut_n13036 (.I0(n12996), .I1(n13034), .I2(n13035), .O(n13036));
  LUT3 #(.INIT(8'h96)) lut_n13037 (.I0(x4638), .I1(x4639), .I2(x4640), .O(n13037));
  LUT5 #(.INIT(32'h96696996)) lut_n13038 (.I0(x4629), .I1(x4630), .I2(x4631), .I3(n13026), .I4(n13027), .O(n13038));
  LUT5 #(.INIT(32'hFF969600)) lut_n13039 (.I0(x4635), .I1(x4636), .I2(x4637), .I3(n13037), .I4(n13038), .O(n13039));
  LUT3 #(.INIT(8'h96)) lut_n13040 (.I0(x4644), .I1(x4645), .I2(x4646), .O(n13040));
  LUT5 #(.INIT(32'h96696996)) lut_n13041 (.I0(x4635), .I1(x4636), .I2(x4637), .I3(n13037), .I4(n13038), .O(n13041));
  LUT5 #(.INIT(32'hFF969600)) lut_n13042 (.I0(x4641), .I1(x4642), .I2(x4643), .I3(n13040), .I4(n13041), .O(n13042));
  LUT3 #(.INIT(8'h96)) lut_n13043 (.I0(n13025), .I1(n13028), .I2(n13029), .O(n13043));
  LUT3 #(.INIT(8'hE8)) lut_n13044 (.I0(n13039), .I1(n13042), .I2(n13043), .O(n13044));
  LUT3 #(.INIT(8'h96)) lut_n13045 (.I0(x4650), .I1(x4651), .I2(x4652), .O(n13045));
  LUT5 #(.INIT(32'h96696996)) lut_n13046 (.I0(x4641), .I1(x4642), .I2(x4643), .I3(n13040), .I4(n13041), .O(n13046));
  LUT5 #(.INIT(32'hFF969600)) lut_n13047 (.I0(x4647), .I1(x4648), .I2(x4649), .I3(n13045), .I4(n13046), .O(n13047));
  LUT3 #(.INIT(8'h96)) lut_n13048 (.I0(x4656), .I1(x4657), .I2(x4658), .O(n13048));
  LUT5 #(.INIT(32'h96696996)) lut_n13049 (.I0(x4647), .I1(x4648), .I2(x4649), .I3(n13045), .I4(n13046), .O(n13049));
  LUT5 #(.INIT(32'hFF969600)) lut_n13050 (.I0(x4653), .I1(x4654), .I2(x4655), .I3(n13048), .I4(n13049), .O(n13050));
  LUT3 #(.INIT(8'h96)) lut_n13051 (.I0(n13039), .I1(n13042), .I2(n13043), .O(n13051));
  LUT3 #(.INIT(8'hE8)) lut_n13052 (.I0(n13047), .I1(n13050), .I2(n13051), .O(n13052));
  LUT3 #(.INIT(8'h96)) lut_n13053 (.I0(n13022), .I1(n13030), .I2(n13031), .O(n13053));
  LUT3 #(.INIT(8'hE8)) lut_n13054 (.I0(n13044), .I1(n13052), .I2(n13053), .O(n13054));
  LUT3 #(.INIT(8'h96)) lut_n13055 (.I0(x4662), .I1(x4663), .I2(x4664), .O(n13055));
  LUT5 #(.INIT(32'h96696996)) lut_n13056 (.I0(x4653), .I1(x4654), .I2(x4655), .I3(n13048), .I4(n13049), .O(n13056));
  LUT5 #(.INIT(32'hFF969600)) lut_n13057 (.I0(x4659), .I1(x4660), .I2(x4661), .I3(n13055), .I4(n13056), .O(n13057));
  LUT3 #(.INIT(8'h96)) lut_n13058 (.I0(x4668), .I1(x4669), .I2(x4670), .O(n13058));
  LUT5 #(.INIT(32'h96696996)) lut_n13059 (.I0(x4659), .I1(x4660), .I2(x4661), .I3(n13055), .I4(n13056), .O(n13059));
  LUT5 #(.INIT(32'hFF969600)) lut_n13060 (.I0(x4665), .I1(x4666), .I2(x4667), .I3(n13058), .I4(n13059), .O(n13060));
  LUT3 #(.INIT(8'h96)) lut_n13061 (.I0(n13047), .I1(n13050), .I2(n13051), .O(n13061));
  LUT3 #(.INIT(8'hE8)) lut_n13062 (.I0(n13057), .I1(n13060), .I2(n13061), .O(n13062));
  LUT3 #(.INIT(8'h96)) lut_n13063 (.I0(x4674), .I1(x4675), .I2(x4676), .O(n13063));
  LUT5 #(.INIT(32'h96696996)) lut_n13064 (.I0(x4665), .I1(x4666), .I2(x4667), .I3(n13058), .I4(n13059), .O(n13064));
  LUT5 #(.INIT(32'hFF969600)) lut_n13065 (.I0(x4671), .I1(x4672), .I2(x4673), .I3(n13063), .I4(n13064), .O(n13065));
  LUT3 #(.INIT(8'h96)) lut_n13066 (.I0(x4680), .I1(x4681), .I2(x4682), .O(n13066));
  LUT5 #(.INIT(32'h96696996)) lut_n13067 (.I0(x4671), .I1(x4672), .I2(x4673), .I3(n13063), .I4(n13064), .O(n13067));
  LUT5 #(.INIT(32'hFF969600)) lut_n13068 (.I0(x4677), .I1(x4678), .I2(x4679), .I3(n13066), .I4(n13067), .O(n13068));
  LUT3 #(.INIT(8'h96)) lut_n13069 (.I0(n13057), .I1(n13060), .I2(n13061), .O(n13069));
  LUT3 #(.INIT(8'hE8)) lut_n13070 (.I0(n13065), .I1(n13068), .I2(n13069), .O(n13070));
  LUT3 #(.INIT(8'h96)) lut_n13071 (.I0(n13044), .I1(n13052), .I2(n13053), .O(n13071));
  LUT3 #(.INIT(8'hE8)) lut_n13072 (.I0(n13062), .I1(n13070), .I2(n13071), .O(n13072));
  LUT3 #(.INIT(8'h96)) lut_n13073 (.I0(n13014), .I1(n13032), .I2(n13033), .O(n13073));
  LUT3 #(.INIT(8'hE8)) lut_n13074 (.I0(n13054), .I1(n13072), .I2(n13073), .O(n13074));
  LUT3 #(.INIT(8'h96)) lut_n13075 (.I0(x4686), .I1(x4687), .I2(x4688), .O(n13075));
  LUT5 #(.INIT(32'h96696996)) lut_n13076 (.I0(x4677), .I1(x4678), .I2(x4679), .I3(n13066), .I4(n13067), .O(n13076));
  LUT5 #(.INIT(32'hFF969600)) lut_n13077 (.I0(x4683), .I1(x4684), .I2(x4685), .I3(n13075), .I4(n13076), .O(n13077));
  LUT3 #(.INIT(8'h96)) lut_n13078 (.I0(x4692), .I1(x4693), .I2(x4694), .O(n13078));
  LUT5 #(.INIT(32'h96696996)) lut_n13079 (.I0(x4683), .I1(x4684), .I2(x4685), .I3(n13075), .I4(n13076), .O(n13079));
  LUT5 #(.INIT(32'hFF969600)) lut_n13080 (.I0(x4689), .I1(x4690), .I2(x4691), .I3(n13078), .I4(n13079), .O(n13080));
  LUT3 #(.INIT(8'h96)) lut_n13081 (.I0(n13065), .I1(n13068), .I2(n13069), .O(n13081));
  LUT3 #(.INIT(8'hE8)) lut_n13082 (.I0(n13077), .I1(n13080), .I2(n13081), .O(n13082));
  LUT3 #(.INIT(8'h96)) lut_n13083 (.I0(x4698), .I1(x4699), .I2(x4700), .O(n13083));
  LUT5 #(.INIT(32'h96696996)) lut_n13084 (.I0(x4689), .I1(x4690), .I2(x4691), .I3(n13078), .I4(n13079), .O(n13084));
  LUT5 #(.INIT(32'hFF969600)) lut_n13085 (.I0(x4695), .I1(x4696), .I2(x4697), .I3(n13083), .I4(n13084), .O(n13085));
  LUT3 #(.INIT(8'h96)) lut_n13086 (.I0(x4704), .I1(x4705), .I2(x4706), .O(n13086));
  LUT5 #(.INIT(32'h96696996)) lut_n13087 (.I0(x4695), .I1(x4696), .I2(x4697), .I3(n13083), .I4(n13084), .O(n13087));
  LUT5 #(.INIT(32'hFF969600)) lut_n13088 (.I0(x4701), .I1(x4702), .I2(x4703), .I3(n13086), .I4(n13087), .O(n13088));
  LUT3 #(.INIT(8'h96)) lut_n13089 (.I0(n13077), .I1(n13080), .I2(n13081), .O(n13089));
  LUT3 #(.INIT(8'hE8)) lut_n13090 (.I0(n13085), .I1(n13088), .I2(n13089), .O(n13090));
  LUT3 #(.INIT(8'h96)) lut_n13091 (.I0(n13062), .I1(n13070), .I2(n13071), .O(n13091));
  LUT3 #(.INIT(8'hE8)) lut_n13092 (.I0(n13082), .I1(n13090), .I2(n13091), .O(n13092));
  LUT3 #(.INIT(8'h96)) lut_n13093 (.I0(x4710), .I1(x4711), .I2(x4712), .O(n13093));
  LUT5 #(.INIT(32'h96696996)) lut_n13094 (.I0(x4701), .I1(x4702), .I2(x4703), .I3(n13086), .I4(n13087), .O(n13094));
  LUT5 #(.INIT(32'hFF969600)) lut_n13095 (.I0(x4707), .I1(x4708), .I2(x4709), .I3(n13093), .I4(n13094), .O(n13095));
  LUT3 #(.INIT(8'h96)) lut_n13096 (.I0(x4716), .I1(x4717), .I2(x4718), .O(n13096));
  LUT5 #(.INIT(32'h96696996)) lut_n13097 (.I0(x4707), .I1(x4708), .I2(x4709), .I3(n13093), .I4(n13094), .O(n13097));
  LUT5 #(.INIT(32'hFF969600)) lut_n13098 (.I0(x4713), .I1(x4714), .I2(x4715), .I3(n13096), .I4(n13097), .O(n13098));
  LUT3 #(.INIT(8'h96)) lut_n13099 (.I0(n13085), .I1(n13088), .I2(n13089), .O(n13099));
  LUT3 #(.INIT(8'hE8)) lut_n13100 (.I0(n13095), .I1(n13098), .I2(n13099), .O(n13100));
  LUT3 #(.INIT(8'h96)) lut_n13101 (.I0(x4722), .I1(x4723), .I2(x4724), .O(n13101));
  LUT5 #(.INIT(32'h96696996)) lut_n13102 (.I0(x4713), .I1(x4714), .I2(x4715), .I3(n13096), .I4(n13097), .O(n13102));
  LUT5 #(.INIT(32'hFF969600)) lut_n13103 (.I0(x4719), .I1(x4720), .I2(x4721), .I3(n13101), .I4(n13102), .O(n13103));
  LUT3 #(.INIT(8'h96)) lut_n13104 (.I0(x4728), .I1(x4729), .I2(x4730), .O(n13104));
  LUT5 #(.INIT(32'h96696996)) lut_n13105 (.I0(x4719), .I1(x4720), .I2(x4721), .I3(n13101), .I4(n13102), .O(n13105));
  LUT5 #(.INIT(32'hFF969600)) lut_n13106 (.I0(x4725), .I1(x4726), .I2(x4727), .I3(n13104), .I4(n13105), .O(n13106));
  LUT3 #(.INIT(8'h96)) lut_n13107 (.I0(n13095), .I1(n13098), .I2(n13099), .O(n13107));
  LUT3 #(.INIT(8'hE8)) lut_n13108 (.I0(n13103), .I1(n13106), .I2(n13107), .O(n13108));
  LUT3 #(.INIT(8'h96)) lut_n13109 (.I0(n13082), .I1(n13090), .I2(n13091), .O(n13109));
  LUT3 #(.INIT(8'hE8)) lut_n13110 (.I0(n13100), .I1(n13108), .I2(n13109), .O(n13110));
  LUT3 #(.INIT(8'h96)) lut_n13111 (.I0(n13054), .I1(n13072), .I2(n13073), .O(n13111));
  LUT3 #(.INIT(8'hE8)) lut_n13112 (.I0(n13092), .I1(n13110), .I2(n13111), .O(n13112));
  LUT3 #(.INIT(8'h96)) lut_n13113 (.I0(n12996), .I1(n13034), .I2(n13035), .O(n13113));
  LUT3 #(.INIT(8'hE8)) lut_n13114 (.I0(n13074), .I1(n13112), .I2(n13113), .O(n13114));
  LUT3 #(.INIT(8'h96)) lut_n13115 (.I0(n12874), .I1(n12952), .I2(n12953), .O(n13115));
  LUT3 #(.INIT(8'hE8)) lut_n13116 (.I0(n13036), .I1(n13114), .I2(n13115), .O(n13116));
  LUT3 #(.INIT(8'h96)) lut_n13117 (.I0(x4734), .I1(x4735), .I2(x4736), .O(n13117));
  LUT5 #(.INIT(32'h96696996)) lut_n13118 (.I0(x4725), .I1(x4726), .I2(x4727), .I3(n13104), .I4(n13105), .O(n13118));
  LUT5 #(.INIT(32'hFF969600)) lut_n13119 (.I0(x4731), .I1(x4732), .I2(x4733), .I3(n13117), .I4(n13118), .O(n13119));
  LUT3 #(.INIT(8'h96)) lut_n13120 (.I0(x4740), .I1(x4741), .I2(x4742), .O(n13120));
  LUT5 #(.INIT(32'h96696996)) lut_n13121 (.I0(x4731), .I1(x4732), .I2(x4733), .I3(n13117), .I4(n13118), .O(n13121));
  LUT5 #(.INIT(32'hFF969600)) lut_n13122 (.I0(x4737), .I1(x4738), .I2(x4739), .I3(n13120), .I4(n13121), .O(n13122));
  LUT3 #(.INIT(8'h96)) lut_n13123 (.I0(n13103), .I1(n13106), .I2(n13107), .O(n13123));
  LUT3 #(.INIT(8'hE8)) lut_n13124 (.I0(n13119), .I1(n13122), .I2(n13123), .O(n13124));
  LUT3 #(.INIT(8'h96)) lut_n13125 (.I0(x4746), .I1(x4747), .I2(x4748), .O(n13125));
  LUT5 #(.INIT(32'h96696996)) lut_n13126 (.I0(x4737), .I1(x4738), .I2(x4739), .I3(n13120), .I4(n13121), .O(n13126));
  LUT5 #(.INIT(32'hFF969600)) lut_n13127 (.I0(x4743), .I1(x4744), .I2(x4745), .I3(n13125), .I4(n13126), .O(n13127));
  LUT3 #(.INIT(8'h96)) lut_n13128 (.I0(x4752), .I1(x4753), .I2(x4754), .O(n13128));
  LUT5 #(.INIT(32'h96696996)) lut_n13129 (.I0(x4743), .I1(x4744), .I2(x4745), .I3(n13125), .I4(n13126), .O(n13129));
  LUT5 #(.INIT(32'hFF969600)) lut_n13130 (.I0(x4749), .I1(x4750), .I2(x4751), .I3(n13128), .I4(n13129), .O(n13130));
  LUT3 #(.INIT(8'h96)) lut_n13131 (.I0(n13119), .I1(n13122), .I2(n13123), .O(n13131));
  LUT3 #(.INIT(8'hE8)) lut_n13132 (.I0(n13127), .I1(n13130), .I2(n13131), .O(n13132));
  LUT3 #(.INIT(8'h96)) lut_n13133 (.I0(n13100), .I1(n13108), .I2(n13109), .O(n13133));
  LUT3 #(.INIT(8'hE8)) lut_n13134 (.I0(n13124), .I1(n13132), .I2(n13133), .O(n13134));
  LUT3 #(.INIT(8'h96)) lut_n13135 (.I0(x4758), .I1(x4759), .I2(x4760), .O(n13135));
  LUT5 #(.INIT(32'h96696996)) lut_n13136 (.I0(x4749), .I1(x4750), .I2(x4751), .I3(n13128), .I4(n13129), .O(n13136));
  LUT5 #(.INIT(32'hFF969600)) lut_n13137 (.I0(x4755), .I1(x4756), .I2(x4757), .I3(n13135), .I4(n13136), .O(n13137));
  LUT3 #(.INIT(8'h96)) lut_n13138 (.I0(x4764), .I1(x4765), .I2(x4766), .O(n13138));
  LUT5 #(.INIT(32'h96696996)) lut_n13139 (.I0(x4755), .I1(x4756), .I2(x4757), .I3(n13135), .I4(n13136), .O(n13139));
  LUT5 #(.INIT(32'hFF969600)) lut_n13140 (.I0(x4761), .I1(x4762), .I2(x4763), .I3(n13138), .I4(n13139), .O(n13140));
  LUT3 #(.INIT(8'h96)) lut_n13141 (.I0(n13127), .I1(n13130), .I2(n13131), .O(n13141));
  LUT3 #(.INIT(8'hE8)) lut_n13142 (.I0(n13137), .I1(n13140), .I2(n13141), .O(n13142));
  LUT3 #(.INIT(8'h96)) lut_n13143 (.I0(x4770), .I1(x4771), .I2(x4772), .O(n13143));
  LUT5 #(.INIT(32'h96696996)) lut_n13144 (.I0(x4761), .I1(x4762), .I2(x4763), .I3(n13138), .I4(n13139), .O(n13144));
  LUT5 #(.INIT(32'hFF969600)) lut_n13145 (.I0(x4767), .I1(x4768), .I2(x4769), .I3(n13143), .I4(n13144), .O(n13145));
  LUT3 #(.INIT(8'h96)) lut_n13146 (.I0(x4776), .I1(x4777), .I2(x4778), .O(n13146));
  LUT5 #(.INIT(32'h96696996)) lut_n13147 (.I0(x4767), .I1(x4768), .I2(x4769), .I3(n13143), .I4(n13144), .O(n13147));
  LUT5 #(.INIT(32'hFF969600)) lut_n13148 (.I0(x4773), .I1(x4774), .I2(x4775), .I3(n13146), .I4(n13147), .O(n13148));
  LUT3 #(.INIT(8'h96)) lut_n13149 (.I0(n13137), .I1(n13140), .I2(n13141), .O(n13149));
  LUT3 #(.INIT(8'hE8)) lut_n13150 (.I0(n13145), .I1(n13148), .I2(n13149), .O(n13150));
  LUT3 #(.INIT(8'h96)) lut_n13151 (.I0(n13124), .I1(n13132), .I2(n13133), .O(n13151));
  LUT3 #(.INIT(8'hE8)) lut_n13152 (.I0(n13142), .I1(n13150), .I2(n13151), .O(n13152));
  LUT3 #(.INIT(8'h96)) lut_n13153 (.I0(n13092), .I1(n13110), .I2(n13111), .O(n13153));
  LUT3 #(.INIT(8'hE8)) lut_n13154 (.I0(n13134), .I1(n13152), .I2(n13153), .O(n13154));
  LUT3 #(.INIT(8'h96)) lut_n13155 (.I0(x4782), .I1(x4783), .I2(x4784), .O(n13155));
  LUT5 #(.INIT(32'h96696996)) lut_n13156 (.I0(x4773), .I1(x4774), .I2(x4775), .I3(n13146), .I4(n13147), .O(n13156));
  LUT5 #(.INIT(32'hFF969600)) lut_n13157 (.I0(x4779), .I1(x4780), .I2(x4781), .I3(n13155), .I4(n13156), .O(n13157));
  LUT3 #(.INIT(8'h96)) lut_n13158 (.I0(x4788), .I1(x4789), .I2(x4790), .O(n13158));
  LUT5 #(.INIT(32'h96696996)) lut_n13159 (.I0(x4779), .I1(x4780), .I2(x4781), .I3(n13155), .I4(n13156), .O(n13159));
  LUT5 #(.INIT(32'hFF969600)) lut_n13160 (.I0(x4785), .I1(x4786), .I2(x4787), .I3(n13158), .I4(n13159), .O(n13160));
  LUT3 #(.INIT(8'h96)) lut_n13161 (.I0(n13145), .I1(n13148), .I2(n13149), .O(n13161));
  LUT3 #(.INIT(8'hE8)) lut_n13162 (.I0(n13157), .I1(n13160), .I2(n13161), .O(n13162));
  LUT3 #(.INIT(8'h96)) lut_n13163 (.I0(x4794), .I1(x4795), .I2(x4796), .O(n13163));
  LUT5 #(.INIT(32'h96696996)) lut_n13164 (.I0(x4785), .I1(x4786), .I2(x4787), .I3(n13158), .I4(n13159), .O(n13164));
  LUT5 #(.INIT(32'hFF969600)) lut_n13165 (.I0(x4791), .I1(x4792), .I2(x4793), .I3(n13163), .I4(n13164), .O(n13165));
  LUT3 #(.INIT(8'h96)) lut_n13166 (.I0(x4800), .I1(x4801), .I2(x4802), .O(n13166));
  LUT5 #(.INIT(32'h96696996)) lut_n13167 (.I0(x4791), .I1(x4792), .I2(x4793), .I3(n13163), .I4(n13164), .O(n13167));
  LUT5 #(.INIT(32'hFF969600)) lut_n13168 (.I0(x4797), .I1(x4798), .I2(x4799), .I3(n13166), .I4(n13167), .O(n13168));
  LUT3 #(.INIT(8'h96)) lut_n13169 (.I0(n13157), .I1(n13160), .I2(n13161), .O(n13169));
  LUT3 #(.INIT(8'hE8)) lut_n13170 (.I0(n13165), .I1(n13168), .I2(n13169), .O(n13170));
  LUT3 #(.INIT(8'h96)) lut_n13171 (.I0(n13142), .I1(n13150), .I2(n13151), .O(n13171));
  LUT3 #(.INIT(8'hE8)) lut_n13172 (.I0(n13162), .I1(n13170), .I2(n13171), .O(n13172));
  LUT3 #(.INIT(8'h96)) lut_n13173 (.I0(x4806), .I1(x4807), .I2(x4808), .O(n13173));
  LUT5 #(.INIT(32'h96696996)) lut_n13174 (.I0(x4797), .I1(x4798), .I2(x4799), .I3(n13166), .I4(n13167), .O(n13174));
  LUT5 #(.INIT(32'hFF969600)) lut_n13175 (.I0(x4803), .I1(x4804), .I2(x4805), .I3(n13173), .I4(n13174), .O(n13175));
  LUT3 #(.INIT(8'h96)) lut_n13176 (.I0(x4812), .I1(x4813), .I2(x4814), .O(n13176));
  LUT5 #(.INIT(32'h96696996)) lut_n13177 (.I0(x4803), .I1(x4804), .I2(x4805), .I3(n13173), .I4(n13174), .O(n13177));
  LUT5 #(.INIT(32'hFF969600)) lut_n13178 (.I0(x4809), .I1(x4810), .I2(x4811), .I3(n13176), .I4(n13177), .O(n13178));
  LUT3 #(.INIT(8'h96)) lut_n13179 (.I0(n13165), .I1(n13168), .I2(n13169), .O(n13179));
  LUT3 #(.INIT(8'hE8)) lut_n13180 (.I0(n13175), .I1(n13178), .I2(n13179), .O(n13180));
  LUT3 #(.INIT(8'h96)) lut_n13181 (.I0(x4818), .I1(x4819), .I2(x4820), .O(n13181));
  LUT5 #(.INIT(32'h96696996)) lut_n13182 (.I0(x4809), .I1(x4810), .I2(x4811), .I3(n13176), .I4(n13177), .O(n13182));
  LUT5 #(.INIT(32'hFF969600)) lut_n13183 (.I0(x4815), .I1(x4816), .I2(x4817), .I3(n13181), .I4(n13182), .O(n13183));
  LUT3 #(.INIT(8'h96)) lut_n13184 (.I0(x4824), .I1(x4825), .I2(x4826), .O(n13184));
  LUT5 #(.INIT(32'h96696996)) lut_n13185 (.I0(x4815), .I1(x4816), .I2(x4817), .I3(n13181), .I4(n13182), .O(n13185));
  LUT5 #(.INIT(32'hFF969600)) lut_n13186 (.I0(x4821), .I1(x4822), .I2(x4823), .I3(n13184), .I4(n13185), .O(n13186));
  LUT3 #(.INIT(8'h96)) lut_n13187 (.I0(n13175), .I1(n13178), .I2(n13179), .O(n13187));
  LUT3 #(.INIT(8'hE8)) lut_n13188 (.I0(n13183), .I1(n13186), .I2(n13187), .O(n13188));
  LUT3 #(.INIT(8'h96)) lut_n13189 (.I0(n13162), .I1(n13170), .I2(n13171), .O(n13189));
  LUT3 #(.INIT(8'hE8)) lut_n13190 (.I0(n13180), .I1(n13188), .I2(n13189), .O(n13190));
  LUT3 #(.INIT(8'h96)) lut_n13191 (.I0(n13134), .I1(n13152), .I2(n13153), .O(n13191));
  LUT3 #(.INIT(8'hE8)) lut_n13192 (.I0(n13172), .I1(n13190), .I2(n13191), .O(n13192));
  LUT3 #(.INIT(8'h96)) lut_n13193 (.I0(n13074), .I1(n13112), .I2(n13113), .O(n13193));
  LUT3 #(.INIT(8'hE8)) lut_n13194 (.I0(n13154), .I1(n13192), .I2(n13193), .O(n13194));
  LUT3 #(.INIT(8'h96)) lut_n13195 (.I0(x4830), .I1(x4831), .I2(x4832), .O(n13195));
  LUT5 #(.INIT(32'h96696996)) lut_n13196 (.I0(x4821), .I1(x4822), .I2(x4823), .I3(n13184), .I4(n13185), .O(n13196));
  LUT5 #(.INIT(32'hFF969600)) lut_n13197 (.I0(x4827), .I1(x4828), .I2(x4829), .I3(n13195), .I4(n13196), .O(n13197));
  LUT3 #(.INIT(8'h96)) lut_n13198 (.I0(x4836), .I1(x4837), .I2(x4838), .O(n13198));
  LUT5 #(.INIT(32'h96696996)) lut_n13199 (.I0(x4827), .I1(x4828), .I2(x4829), .I3(n13195), .I4(n13196), .O(n13199));
  LUT5 #(.INIT(32'hFF969600)) lut_n13200 (.I0(x4833), .I1(x4834), .I2(x4835), .I3(n13198), .I4(n13199), .O(n13200));
  LUT3 #(.INIT(8'h96)) lut_n13201 (.I0(n13183), .I1(n13186), .I2(n13187), .O(n13201));
  LUT3 #(.INIT(8'hE8)) lut_n13202 (.I0(n13197), .I1(n13200), .I2(n13201), .O(n13202));
  LUT3 #(.INIT(8'h96)) lut_n13203 (.I0(x4842), .I1(x4843), .I2(x4844), .O(n13203));
  LUT5 #(.INIT(32'h96696996)) lut_n13204 (.I0(x4833), .I1(x4834), .I2(x4835), .I3(n13198), .I4(n13199), .O(n13204));
  LUT5 #(.INIT(32'hFF969600)) lut_n13205 (.I0(x4839), .I1(x4840), .I2(x4841), .I3(n13203), .I4(n13204), .O(n13205));
  LUT3 #(.INIT(8'h96)) lut_n13206 (.I0(x4848), .I1(x4849), .I2(x4850), .O(n13206));
  LUT5 #(.INIT(32'h96696996)) lut_n13207 (.I0(x4839), .I1(x4840), .I2(x4841), .I3(n13203), .I4(n13204), .O(n13207));
  LUT5 #(.INIT(32'hFF969600)) lut_n13208 (.I0(x4845), .I1(x4846), .I2(x4847), .I3(n13206), .I4(n13207), .O(n13208));
  LUT3 #(.INIT(8'h96)) lut_n13209 (.I0(n13197), .I1(n13200), .I2(n13201), .O(n13209));
  LUT3 #(.INIT(8'hE8)) lut_n13210 (.I0(n13205), .I1(n13208), .I2(n13209), .O(n13210));
  LUT3 #(.INIT(8'h96)) lut_n13211 (.I0(n13180), .I1(n13188), .I2(n13189), .O(n13211));
  LUT3 #(.INIT(8'hE8)) lut_n13212 (.I0(n13202), .I1(n13210), .I2(n13211), .O(n13212));
  LUT3 #(.INIT(8'h96)) lut_n13213 (.I0(x4854), .I1(x4855), .I2(x4856), .O(n13213));
  LUT5 #(.INIT(32'h96696996)) lut_n13214 (.I0(x4845), .I1(x4846), .I2(x4847), .I3(n13206), .I4(n13207), .O(n13214));
  LUT5 #(.INIT(32'hFF969600)) lut_n13215 (.I0(x4851), .I1(x4852), .I2(x4853), .I3(n13213), .I4(n13214), .O(n13215));
  LUT3 #(.INIT(8'h96)) lut_n13216 (.I0(x4860), .I1(x4861), .I2(x4862), .O(n13216));
  LUT5 #(.INIT(32'h96696996)) lut_n13217 (.I0(x4851), .I1(x4852), .I2(x4853), .I3(n13213), .I4(n13214), .O(n13217));
  LUT5 #(.INIT(32'hFF969600)) lut_n13218 (.I0(x4857), .I1(x4858), .I2(x4859), .I3(n13216), .I4(n13217), .O(n13218));
  LUT3 #(.INIT(8'h96)) lut_n13219 (.I0(n13205), .I1(n13208), .I2(n13209), .O(n13219));
  LUT3 #(.INIT(8'hE8)) lut_n13220 (.I0(n13215), .I1(n13218), .I2(n13219), .O(n13220));
  LUT3 #(.INIT(8'h96)) lut_n13221 (.I0(x4866), .I1(x4867), .I2(x4868), .O(n13221));
  LUT5 #(.INIT(32'h96696996)) lut_n13222 (.I0(x4857), .I1(x4858), .I2(x4859), .I3(n13216), .I4(n13217), .O(n13222));
  LUT5 #(.INIT(32'hFF969600)) lut_n13223 (.I0(x4863), .I1(x4864), .I2(x4865), .I3(n13221), .I4(n13222), .O(n13223));
  LUT3 #(.INIT(8'h96)) lut_n13224 (.I0(x4872), .I1(x4873), .I2(x4874), .O(n13224));
  LUT5 #(.INIT(32'h96696996)) lut_n13225 (.I0(x4863), .I1(x4864), .I2(x4865), .I3(n13221), .I4(n13222), .O(n13225));
  LUT5 #(.INIT(32'hFF969600)) lut_n13226 (.I0(x4869), .I1(x4870), .I2(x4871), .I3(n13224), .I4(n13225), .O(n13226));
  LUT3 #(.INIT(8'h96)) lut_n13227 (.I0(n13215), .I1(n13218), .I2(n13219), .O(n13227));
  LUT3 #(.INIT(8'hE8)) lut_n13228 (.I0(n13223), .I1(n13226), .I2(n13227), .O(n13228));
  LUT3 #(.INIT(8'h96)) lut_n13229 (.I0(n13202), .I1(n13210), .I2(n13211), .O(n13229));
  LUT3 #(.INIT(8'hE8)) lut_n13230 (.I0(n13220), .I1(n13228), .I2(n13229), .O(n13230));
  LUT3 #(.INIT(8'h96)) lut_n13231 (.I0(n13172), .I1(n13190), .I2(n13191), .O(n13231));
  LUT3 #(.INIT(8'hE8)) lut_n13232 (.I0(n13212), .I1(n13230), .I2(n13231), .O(n13232));
  LUT3 #(.INIT(8'h96)) lut_n13233 (.I0(x4878), .I1(x4879), .I2(x4880), .O(n13233));
  LUT5 #(.INIT(32'h96696996)) lut_n13234 (.I0(x4869), .I1(x4870), .I2(x4871), .I3(n13224), .I4(n13225), .O(n13234));
  LUT5 #(.INIT(32'hFF969600)) lut_n13235 (.I0(x4875), .I1(x4876), .I2(x4877), .I3(n13233), .I4(n13234), .O(n13235));
  LUT3 #(.INIT(8'h96)) lut_n13236 (.I0(x4884), .I1(x4885), .I2(x4886), .O(n13236));
  LUT5 #(.INIT(32'h96696996)) lut_n13237 (.I0(x4875), .I1(x4876), .I2(x4877), .I3(n13233), .I4(n13234), .O(n13237));
  LUT5 #(.INIT(32'hFF969600)) lut_n13238 (.I0(x4881), .I1(x4882), .I2(x4883), .I3(n13236), .I4(n13237), .O(n13238));
  LUT3 #(.INIT(8'h96)) lut_n13239 (.I0(n13223), .I1(n13226), .I2(n13227), .O(n13239));
  LUT3 #(.INIT(8'hE8)) lut_n13240 (.I0(n13235), .I1(n13238), .I2(n13239), .O(n13240));
  LUT3 #(.INIT(8'h96)) lut_n13241 (.I0(x4890), .I1(x4891), .I2(x4892), .O(n13241));
  LUT5 #(.INIT(32'h96696996)) lut_n13242 (.I0(x4881), .I1(x4882), .I2(x4883), .I3(n13236), .I4(n13237), .O(n13242));
  LUT5 #(.INIT(32'hFF969600)) lut_n13243 (.I0(x4887), .I1(x4888), .I2(x4889), .I3(n13241), .I4(n13242), .O(n13243));
  LUT3 #(.INIT(8'h96)) lut_n13244 (.I0(x4896), .I1(x4897), .I2(x4898), .O(n13244));
  LUT5 #(.INIT(32'h96696996)) lut_n13245 (.I0(x4887), .I1(x4888), .I2(x4889), .I3(n13241), .I4(n13242), .O(n13245));
  LUT5 #(.INIT(32'hFF969600)) lut_n13246 (.I0(x4893), .I1(x4894), .I2(x4895), .I3(n13244), .I4(n13245), .O(n13246));
  LUT3 #(.INIT(8'h96)) lut_n13247 (.I0(n13235), .I1(n13238), .I2(n13239), .O(n13247));
  LUT3 #(.INIT(8'hE8)) lut_n13248 (.I0(n13243), .I1(n13246), .I2(n13247), .O(n13248));
  LUT3 #(.INIT(8'h96)) lut_n13249 (.I0(n13220), .I1(n13228), .I2(n13229), .O(n13249));
  LUT3 #(.INIT(8'hE8)) lut_n13250 (.I0(n13240), .I1(n13248), .I2(n13249), .O(n13250));
  LUT3 #(.INIT(8'h96)) lut_n13251 (.I0(x4902), .I1(x4903), .I2(x4904), .O(n13251));
  LUT5 #(.INIT(32'h96696996)) lut_n13252 (.I0(x4893), .I1(x4894), .I2(x4895), .I3(n13244), .I4(n13245), .O(n13252));
  LUT5 #(.INIT(32'hFF969600)) lut_n13253 (.I0(x4899), .I1(x4900), .I2(x4901), .I3(n13251), .I4(n13252), .O(n13253));
  LUT3 #(.INIT(8'h96)) lut_n13254 (.I0(x4908), .I1(x4909), .I2(x4910), .O(n13254));
  LUT5 #(.INIT(32'h96696996)) lut_n13255 (.I0(x4899), .I1(x4900), .I2(x4901), .I3(n13251), .I4(n13252), .O(n13255));
  LUT5 #(.INIT(32'hFF969600)) lut_n13256 (.I0(x4905), .I1(x4906), .I2(x4907), .I3(n13254), .I4(n13255), .O(n13256));
  LUT3 #(.INIT(8'h96)) lut_n13257 (.I0(n13243), .I1(n13246), .I2(n13247), .O(n13257));
  LUT3 #(.INIT(8'hE8)) lut_n13258 (.I0(n13253), .I1(n13256), .I2(n13257), .O(n13258));
  LUT3 #(.INIT(8'h96)) lut_n13259 (.I0(x4914), .I1(x4915), .I2(x4916), .O(n13259));
  LUT5 #(.INIT(32'h96696996)) lut_n13260 (.I0(x4905), .I1(x4906), .I2(x4907), .I3(n13254), .I4(n13255), .O(n13260));
  LUT5 #(.INIT(32'hFF969600)) lut_n13261 (.I0(x4911), .I1(x4912), .I2(x4913), .I3(n13259), .I4(n13260), .O(n13261));
  LUT3 #(.INIT(8'h96)) lut_n13262 (.I0(x4920), .I1(x4921), .I2(x4922), .O(n13262));
  LUT5 #(.INIT(32'h96696996)) lut_n13263 (.I0(x4911), .I1(x4912), .I2(x4913), .I3(n13259), .I4(n13260), .O(n13263));
  LUT5 #(.INIT(32'hFF969600)) lut_n13264 (.I0(x4917), .I1(x4918), .I2(x4919), .I3(n13262), .I4(n13263), .O(n13264));
  LUT3 #(.INIT(8'h96)) lut_n13265 (.I0(n13253), .I1(n13256), .I2(n13257), .O(n13265));
  LUT3 #(.INIT(8'hE8)) lut_n13266 (.I0(n13261), .I1(n13264), .I2(n13265), .O(n13266));
  LUT3 #(.INIT(8'h96)) lut_n13267 (.I0(n13240), .I1(n13248), .I2(n13249), .O(n13267));
  LUT3 #(.INIT(8'hE8)) lut_n13268 (.I0(n13258), .I1(n13266), .I2(n13267), .O(n13268));
  LUT3 #(.INIT(8'h96)) lut_n13269 (.I0(n13212), .I1(n13230), .I2(n13231), .O(n13269));
  LUT3 #(.INIT(8'hE8)) lut_n13270 (.I0(n13250), .I1(n13268), .I2(n13269), .O(n13270));
  LUT3 #(.INIT(8'h96)) lut_n13271 (.I0(n13154), .I1(n13192), .I2(n13193), .O(n13271));
  LUT3 #(.INIT(8'hE8)) lut_n13272 (.I0(n13232), .I1(n13270), .I2(n13271), .O(n13272));
  LUT3 #(.INIT(8'h96)) lut_n13273 (.I0(n13036), .I1(n13114), .I2(n13115), .O(n13273));
  LUT3 #(.INIT(8'hE8)) lut_n13274 (.I0(n13194), .I1(n13272), .I2(n13273), .O(n13274));
  LUT3 #(.INIT(8'h96)) lut_n13275 (.I0(n12796), .I1(n12954), .I2(n12955), .O(n13275));
  LUT3 #(.INIT(8'hE8)) lut_n13276 (.I0(n13116), .I1(n13274), .I2(n13275), .O(n13276));
  LUT3 #(.INIT(8'h96)) lut_n13277 (.I0(x4926), .I1(x4927), .I2(x4928), .O(n13277));
  LUT5 #(.INIT(32'h96696996)) lut_n13278 (.I0(x4917), .I1(x4918), .I2(x4919), .I3(n13262), .I4(n13263), .O(n13278));
  LUT5 #(.INIT(32'hFF969600)) lut_n13279 (.I0(x4923), .I1(x4924), .I2(x4925), .I3(n13277), .I4(n13278), .O(n13279));
  LUT3 #(.INIT(8'h96)) lut_n13280 (.I0(x4932), .I1(x4933), .I2(x4934), .O(n13280));
  LUT5 #(.INIT(32'h96696996)) lut_n13281 (.I0(x4923), .I1(x4924), .I2(x4925), .I3(n13277), .I4(n13278), .O(n13281));
  LUT5 #(.INIT(32'hFF969600)) lut_n13282 (.I0(x4929), .I1(x4930), .I2(x4931), .I3(n13280), .I4(n13281), .O(n13282));
  LUT3 #(.INIT(8'h96)) lut_n13283 (.I0(n13261), .I1(n13264), .I2(n13265), .O(n13283));
  LUT3 #(.INIT(8'hE8)) lut_n13284 (.I0(n13279), .I1(n13282), .I2(n13283), .O(n13284));
  LUT3 #(.INIT(8'h96)) lut_n13285 (.I0(x4938), .I1(x4939), .I2(x4940), .O(n13285));
  LUT5 #(.INIT(32'h96696996)) lut_n13286 (.I0(x4929), .I1(x4930), .I2(x4931), .I3(n13280), .I4(n13281), .O(n13286));
  LUT5 #(.INIT(32'hFF969600)) lut_n13287 (.I0(x4935), .I1(x4936), .I2(x4937), .I3(n13285), .I4(n13286), .O(n13287));
  LUT3 #(.INIT(8'h96)) lut_n13288 (.I0(x4944), .I1(x4945), .I2(x4946), .O(n13288));
  LUT5 #(.INIT(32'h96696996)) lut_n13289 (.I0(x4935), .I1(x4936), .I2(x4937), .I3(n13285), .I4(n13286), .O(n13289));
  LUT5 #(.INIT(32'hFF969600)) lut_n13290 (.I0(x4941), .I1(x4942), .I2(x4943), .I3(n13288), .I4(n13289), .O(n13290));
  LUT3 #(.INIT(8'h96)) lut_n13291 (.I0(n13279), .I1(n13282), .I2(n13283), .O(n13291));
  LUT3 #(.INIT(8'hE8)) lut_n13292 (.I0(n13287), .I1(n13290), .I2(n13291), .O(n13292));
  LUT3 #(.INIT(8'h96)) lut_n13293 (.I0(n13258), .I1(n13266), .I2(n13267), .O(n13293));
  LUT3 #(.INIT(8'hE8)) lut_n13294 (.I0(n13284), .I1(n13292), .I2(n13293), .O(n13294));
  LUT3 #(.INIT(8'h96)) lut_n13295 (.I0(x4950), .I1(x4951), .I2(x4952), .O(n13295));
  LUT5 #(.INIT(32'h96696996)) lut_n13296 (.I0(x4941), .I1(x4942), .I2(x4943), .I3(n13288), .I4(n13289), .O(n13296));
  LUT5 #(.INIT(32'hFF969600)) lut_n13297 (.I0(x4947), .I1(x4948), .I2(x4949), .I3(n13295), .I4(n13296), .O(n13297));
  LUT3 #(.INIT(8'h96)) lut_n13298 (.I0(x4956), .I1(x4957), .I2(x4958), .O(n13298));
  LUT5 #(.INIT(32'h96696996)) lut_n13299 (.I0(x4947), .I1(x4948), .I2(x4949), .I3(n13295), .I4(n13296), .O(n13299));
  LUT5 #(.INIT(32'hFF969600)) lut_n13300 (.I0(x4953), .I1(x4954), .I2(x4955), .I3(n13298), .I4(n13299), .O(n13300));
  LUT3 #(.INIT(8'h96)) lut_n13301 (.I0(n13287), .I1(n13290), .I2(n13291), .O(n13301));
  LUT3 #(.INIT(8'hE8)) lut_n13302 (.I0(n13297), .I1(n13300), .I2(n13301), .O(n13302));
  LUT3 #(.INIT(8'h96)) lut_n13303 (.I0(x4962), .I1(x4963), .I2(x4964), .O(n13303));
  LUT5 #(.INIT(32'h96696996)) lut_n13304 (.I0(x4953), .I1(x4954), .I2(x4955), .I3(n13298), .I4(n13299), .O(n13304));
  LUT5 #(.INIT(32'hFF969600)) lut_n13305 (.I0(x4959), .I1(x4960), .I2(x4961), .I3(n13303), .I4(n13304), .O(n13305));
  LUT3 #(.INIT(8'h96)) lut_n13306 (.I0(x4968), .I1(x4969), .I2(x4970), .O(n13306));
  LUT5 #(.INIT(32'h96696996)) lut_n13307 (.I0(x4959), .I1(x4960), .I2(x4961), .I3(n13303), .I4(n13304), .O(n13307));
  LUT5 #(.INIT(32'hFF969600)) lut_n13308 (.I0(x4965), .I1(x4966), .I2(x4967), .I3(n13306), .I4(n13307), .O(n13308));
  LUT3 #(.INIT(8'h96)) lut_n13309 (.I0(n13297), .I1(n13300), .I2(n13301), .O(n13309));
  LUT3 #(.INIT(8'hE8)) lut_n13310 (.I0(n13305), .I1(n13308), .I2(n13309), .O(n13310));
  LUT3 #(.INIT(8'h96)) lut_n13311 (.I0(n13284), .I1(n13292), .I2(n13293), .O(n13311));
  LUT3 #(.INIT(8'hE8)) lut_n13312 (.I0(n13302), .I1(n13310), .I2(n13311), .O(n13312));
  LUT3 #(.INIT(8'h96)) lut_n13313 (.I0(n13250), .I1(n13268), .I2(n13269), .O(n13313));
  LUT3 #(.INIT(8'hE8)) lut_n13314 (.I0(n13294), .I1(n13312), .I2(n13313), .O(n13314));
  LUT3 #(.INIT(8'h96)) lut_n13315 (.I0(x4974), .I1(x4975), .I2(x4976), .O(n13315));
  LUT5 #(.INIT(32'h96696996)) lut_n13316 (.I0(x4965), .I1(x4966), .I2(x4967), .I3(n13306), .I4(n13307), .O(n13316));
  LUT5 #(.INIT(32'hFF969600)) lut_n13317 (.I0(x4971), .I1(x4972), .I2(x4973), .I3(n13315), .I4(n13316), .O(n13317));
  LUT3 #(.INIT(8'h96)) lut_n13318 (.I0(x4980), .I1(x4981), .I2(x4982), .O(n13318));
  LUT5 #(.INIT(32'h96696996)) lut_n13319 (.I0(x4971), .I1(x4972), .I2(x4973), .I3(n13315), .I4(n13316), .O(n13319));
  LUT5 #(.INIT(32'hFF969600)) lut_n13320 (.I0(x4977), .I1(x4978), .I2(x4979), .I3(n13318), .I4(n13319), .O(n13320));
  LUT3 #(.INIT(8'h96)) lut_n13321 (.I0(n13305), .I1(n13308), .I2(n13309), .O(n13321));
  LUT3 #(.INIT(8'hE8)) lut_n13322 (.I0(n13317), .I1(n13320), .I2(n13321), .O(n13322));
  LUT3 #(.INIT(8'h96)) lut_n13323 (.I0(x4986), .I1(x4987), .I2(x4988), .O(n13323));
  LUT5 #(.INIT(32'h96696996)) lut_n13324 (.I0(x4977), .I1(x4978), .I2(x4979), .I3(n13318), .I4(n13319), .O(n13324));
  LUT5 #(.INIT(32'hFF969600)) lut_n13325 (.I0(x4983), .I1(x4984), .I2(x4985), .I3(n13323), .I4(n13324), .O(n13325));
  LUT3 #(.INIT(8'h96)) lut_n13326 (.I0(x4992), .I1(x4993), .I2(x4994), .O(n13326));
  LUT5 #(.INIT(32'h96696996)) lut_n13327 (.I0(x4983), .I1(x4984), .I2(x4985), .I3(n13323), .I4(n13324), .O(n13327));
  LUT5 #(.INIT(32'hFF969600)) lut_n13328 (.I0(x4989), .I1(x4990), .I2(x4991), .I3(n13326), .I4(n13327), .O(n13328));
  LUT3 #(.INIT(8'h96)) lut_n13329 (.I0(n13317), .I1(n13320), .I2(n13321), .O(n13329));
  LUT3 #(.INIT(8'hE8)) lut_n13330 (.I0(n13325), .I1(n13328), .I2(n13329), .O(n13330));
  LUT3 #(.INIT(8'h96)) lut_n13331 (.I0(n13302), .I1(n13310), .I2(n13311), .O(n13331));
  LUT3 #(.INIT(8'hE8)) lut_n13332 (.I0(n13322), .I1(n13330), .I2(n13331), .O(n13332));
  LUT3 #(.INIT(8'h96)) lut_n13333 (.I0(x4998), .I1(x4999), .I2(x5000), .O(n13333));
  LUT5 #(.INIT(32'h96696996)) lut_n13334 (.I0(x4989), .I1(x4990), .I2(x4991), .I3(n13326), .I4(n13327), .O(n13334));
  LUT5 #(.INIT(32'hFF969600)) lut_n13335 (.I0(x4995), .I1(x4996), .I2(x4997), .I3(n13333), .I4(n13334), .O(n13335));
  LUT3 #(.INIT(8'h96)) lut_n13336 (.I0(x5004), .I1(x5005), .I2(x5006), .O(n13336));
  LUT5 #(.INIT(32'h96696996)) lut_n13337 (.I0(x4995), .I1(x4996), .I2(x4997), .I3(n13333), .I4(n13334), .O(n13337));
  LUT5 #(.INIT(32'hFF969600)) lut_n13338 (.I0(x5001), .I1(x5002), .I2(x5003), .I3(n13336), .I4(n13337), .O(n13338));
  LUT3 #(.INIT(8'h96)) lut_n13339 (.I0(n13325), .I1(n13328), .I2(n13329), .O(n13339));
  LUT3 #(.INIT(8'hE8)) lut_n13340 (.I0(n13335), .I1(n13338), .I2(n13339), .O(n13340));
  LUT3 #(.INIT(8'h96)) lut_n13341 (.I0(x5010), .I1(x5011), .I2(x5012), .O(n13341));
  LUT5 #(.INIT(32'h96696996)) lut_n13342 (.I0(x5001), .I1(x5002), .I2(x5003), .I3(n13336), .I4(n13337), .O(n13342));
  LUT5 #(.INIT(32'hFF969600)) lut_n13343 (.I0(x5007), .I1(x5008), .I2(x5009), .I3(n13341), .I4(n13342), .O(n13343));
  LUT3 #(.INIT(8'h96)) lut_n13344 (.I0(x5016), .I1(x5017), .I2(x5018), .O(n13344));
  LUT5 #(.INIT(32'h96696996)) lut_n13345 (.I0(x5007), .I1(x5008), .I2(x5009), .I3(n13341), .I4(n13342), .O(n13345));
  LUT5 #(.INIT(32'hFF969600)) lut_n13346 (.I0(x5013), .I1(x5014), .I2(x5015), .I3(n13344), .I4(n13345), .O(n13346));
  LUT3 #(.INIT(8'h96)) lut_n13347 (.I0(n13335), .I1(n13338), .I2(n13339), .O(n13347));
  LUT3 #(.INIT(8'hE8)) lut_n13348 (.I0(n13343), .I1(n13346), .I2(n13347), .O(n13348));
  LUT3 #(.INIT(8'h96)) lut_n13349 (.I0(n13322), .I1(n13330), .I2(n13331), .O(n13349));
  LUT3 #(.INIT(8'hE8)) lut_n13350 (.I0(n13340), .I1(n13348), .I2(n13349), .O(n13350));
  LUT3 #(.INIT(8'h96)) lut_n13351 (.I0(n13294), .I1(n13312), .I2(n13313), .O(n13351));
  LUT3 #(.INIT(8'hE8)) lut_n13352 (.I0(n13332), .I1(n13350), .I2(n13351), .O(n13352));
  LUT3 #(.INIT(8'h96)) lut_n13353 (.I0(n13232), .I1(n13270), .I2(n13271), .O(n13353));
  LUT3 #(.INIT(8'hE8)) lut_n13354 (.I0(n13314), .I1(n13352), .I2(n13353), .O(n13354));
  LUT3 #(.INIT(8'h96)) lut_n13355 (.I0(x5019), .I1(x5020), .I2(x5021), .O(n13355));
  LUT5 #(.INIT(32'h96696996)) lut_n13356 (.I0(x5013), .I1(x5014), .I2(x5015), .I3(n13344), .I4(n13345), .O(n13356));
  LUT3 #(.INIT(8'h96)) lut_n13357 (.I0(n13343), .I1(n13346), .I2(n13347), .O(n13357));
  LUT6 #(.INIT(64'hFFFFFF9696000000)) lut_n13358 (.I0(x5022), .I1(x5023), .I2(x5024), .I3(n13355), .I4(n13356), .I5(n13357), .O(n13358));
  LUT6 #(.INIT(64'h9600006969FFFF96)) lut_n13359 (.I0(x5022), .I1(x5023), .I2(x5024), .I3(n13355), .I4(n13356), .I5(n13357), .O(n13359));
  LUT3 #(.INIT(8'h96)) lut_n13360 (.I0(n13340), .I1(n13348), .I2(n13349), .O(n13360));
  LUT3 #(.INIT(8'h96)) lut_n13361 (.I0(n13332), .I1(n13350), .I2(n13351), .O(n13361));
  LUT3 #(.INIT(8'h96)) lut_n13362 (.I0(n13314), .I1(n13352), .I2(n13353), .O(n13362));
  LUT5 #(.INIT(32'hFFFE8000)) lut_n13363 (.I0(n13358), .I1(n13359), .I2(n13360), .I3(n13361), .I4(n13362), .O(n13363));
  LUT3 #(.INIT(8'h96)) lut_n13364 (.I0(n13194), .I1(n13272), .I2(n13273), .O(n13364));
  LUT6 #(.INIT(64'hFF96969696969600)) lut_n13365 (.I0(n13116), .I1(n13274), .I2(n13275), .I3(n13354), .I4(n13363), .I5(n13364), .O(n13365));
  LUT5 #(.INIT(32'hFF969600)) lut_n13366 (.I0(n12638), .I1(n12956), .I2(n12957), .I3(n13276), .I4(n13365), .O(n13366));
  LUT5 #(.INIT(32'hFF969600)) lut_n13367 (.I0(n11680), .I1(n12318), .I2(n12319), .I3(n12958), .I4(n13366), .O(n13367));
  LUT3 #(.INIT(8'h96)) lut_n13368 (.I0(n9761), .I1(n11039), .I2(n11040), .O(n13368));
  LUT6 #(.INIT(64'hFF96969696969600)) lut_n13369 (.I0(n7555), .I1(n8833), .I2(n11041), .I3(n12320), .I4(n13367), .I5(n13368), .O(n13369));
  LUT6 #(.INIT(64'h9669696969696996)) lut_n13370 (.I0(n7555), .I1(n8833), .I2(n11041), .I3(n12320), .I4(n13367), .I5(n13368), .O(n13370));
  LUT3 #(.INIT(8'hE8)) lut_n13371 (.I0(n11042), .I1(n13369), .I2(n13370), .O(n13371));
  assign y0 = n13371;
endmodule
