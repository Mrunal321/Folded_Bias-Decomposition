`timescale 1ns/1ps
`default_nettype none

module tb_top;
  // 127-bit input vector
  reg  [126:0] x = 127'b0;
  wire       y0;
  reg  [63:0] idx;

  // DUT instantiation
  top dut (
    .x0(x[0]), .x1(x[1]), .x2(x[2]), .x3(x[3]), .x4(x[4]), .x5(x[5]), .x6(x[6]), .x7(x[7]), .x8(x[8]), .x9(x[9]), .x10(x[10]), .x11(x[11]), .x12(x[12]), .x13(x[13]), .x14(x[14]), .x15(x[15]), .x16(x[16]), .x17(x[17]), .x18(x[18]), .x19(x[19]), .x20(x[20]), .x21(x[21]), .x22(x[22]), .x23(x[23]), .x24(x[24]), .x25(x[25]), .x26(x[26]), .x27(x[27]), .x28(x[28]), .x29(x[29]), .x30(x[30]), .x31(x[31]), .x32(x[32]), .x33(x[33]), .x34(x[34]), .x35(x[35]), .x36(x[36]), .x37(x[37]), .x38(x[38]), .x39(x[39]), .x40(x[40]), .x41(x[41]), .x42(x[42]), .x43(x[43]), .x44(x[44]), .x45(x[45]), .x46(x[46]), .x47(x[47]), .x48(x[48]), .x49(x[49]), .x50(x[50]), .x51(x[51]), .x52(x[52]), .x53(x[53]), .x54(x[54]), .x55(x[55]), .x56(x[56]), .x57(x[57]), .x58(x[58]), .x59(x[59]), .x60(x[60]), .x61(x[61]), .x62(x[62]), .x63(x[63]), .x64(x[64]), .x65(x[65]), .x66(x[66]), .x67(x[67]), .x68(x[68]), .x69(x[69]), .x70(x[70]), .x71(x[71]), .x72(x[72]), .x73(x[73]), .x74(x[74]), .x75(x[75]), .x76(x[76]), .x77(x[77]), .x78(x[78]), .x79(x[79]), .x80(x[80]), .x81(x[81]), .x82(x[82]), .x83(x[83]), .x84(x[84]), .x85(x[85]), .x86(x[86]), .x87(x[87]), .x88(x[88]), .x89(x[89]), .x90(x[90]), .x91(x[91]), .x92(x[92]), .x93(x[93]), .x94(x[94]), .x95(x[95]), .x96(x[96]), .x97(x[97]), .x98(x[98]), .x99(x[99]), .x100(x[100]), .x101(x[101]), .x102(x[102]), .x103(x[103]), .x104(x[104]), .x105(x[105]), .x106(x[106]), .x107(x[107]), .x108(x[108]), .x109(x[109]), .x110(x[110]), .x111(x[111]), .x112(x[112]), .x113(x[113]), .x114(x[114]), .x115(x[115]), .x116(x[116]), .x117(x[117]), .x118(x[118]), .x119(x[119]), .x120(x[120]), .x121(x[121]), .x122(x[122]), .x123(x[123]), .x124(x[124]), .x125(x[125]), .x126(x[126]),
    .y0(y0)
  );

  // Optional reference function (majority reference for sanity check)
  function [6:0] popcount(input [126:0] v);
    integer i; reg [6:0] c;
    begin
      c = 0;
      for (i = 0; i < 127; i = i + 1)
        c = c + v[i];
      popcount = c;
    end
  endfunction

  // Reference majority: at least 64 ones
  wire y_ref = (popcount(x) >= 64);

  localparam [63:0] TOTAL_VECTORS = 64'd170141183460469231731687303715884105728;

  initial begin
    $display("Time | x126 x125 x124 x123 x122 x121 x120 x119 x118 x117 x116 x115 x114 x113 x112 x111 x110 x109 x108 x107 x106 x105 x104 x103 x102 x101 x100 x99 x98 x97 x96 x95 x94 x93 x92 x91 x90 x89 x88 x87 x86 x85 x84 x83 x82 x81 x80 x79 x78 x77 x76 x75 x74 x73 x72 x71 x70 x69 x68 x67 x66 x65 x64 x63 x62 x61 x60 x59 x58 x57 x56 x55 x54 x53 x52 x51 x50 x49 x48 x47 x46 x45 x44 x43 x42 x41 x40 x39 x38 x37 x36 x35 x34 x33 x32 x31 x30 x29 x28 x27 x26 x25 x24 x23 x22 x21 x20 x19 x18 x17 x16 x15 x14 x13 x12 x11 x10 x9 x8 x7 x6 x5 x4 x3 x2 x1 x0 | y0 (DUT) y_ref (Maj127)");
    $display("-----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------");
    // Loop through all 170141183460469231731687303715884105728 combinations
    for (idx = 0; idx < TOTAL_VECTORS; idx = idx + 1) begin
      x = idx[126:0];
      #10 $display("%4t |  %b  |   %b       %b",
                   $time, x, y0, y_ref);
    end
    #10 $finish;
  end

  // Optional mismatch check
  always #1 if (^x !== 1'bx && y0 !== y_ref)
    $display("Mismatch at t=%0t x=%b HW=%0d y0=%0b ref=%0b",
             $time, x, popcount(x), y0, y_ref);

endmodule

`default_nettype wire
