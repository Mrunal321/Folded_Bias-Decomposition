module top (x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, y0);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42;
  output y0;
  wire n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104;
  LUT3 #(.INIT(8'hE8)) lut_n45 (.I0(x0), .I1(x1), .I2(x2), .O(n45));
  LUT3 #(.INIT(8'hE8)) lut_n46 (.I0(x6), .I1(x7), .I2(x8), .O(n46));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n47 (.I0(x3), .I1(x4), .I2(x5), .I3(n45), .I4(n46), .O(n47));
  LUT3 #(.INIT(8'hE8)) lut_n48 (.I0(x12), .I1(x13), .I2(x14), .O(n48));
  LUT5 #(.INIT(32'hE81717E8)) lut_n49 (.I0(x3), .I1(x4), .I2(x5), .I3(n45), .I4(n46), .O(n49));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n50 (.I0(x9), .I1(x10), .I2(x11), .I3(n48), .I4(n49), .O(n50));
  LUT3 #(.INIT(8'hE8)) lut_n51 (.I0(x18), .I1(x19), .I2(x20), .O(n51));
  LUT5 #(.INIT(32'hE81717E8)) lut_n52 (.I0(x9), .I1(x10), .I2(x11), .I3(n48), .I4(n49), .O(n52));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n53 (.I0(x15), .I1(x16), .I2(x17), .I3(n51), .I4(n52), .O(n53));
  LUT3 #(.INIT(8'hE8)) lut_n54 (.I0(n47), .I1(n50), .I2(n53), .O(n54));
  LUT3 #(.INIT(8'hE8)) lut_n55 (.I0(x24), .I1(x25), .I2(x26), .O(n55));
  LUT5 #(.INIT(32'hE81717E8)) lut_n56 (.I0(x15), .I1(x16), .I2(x17), .I3(n51), .I4(n52), .O(n56));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n57 (.I0(x21), .I1(x22), .I2(x23), .I3(n55), .I4(n56), .O(n57));
  LUT3 #(.INIT(8'hE8)) lut_n58 (.I0(x27), .I1(x28), .I2(x29), .O(n58));
  LUT5 #(.INIT(32'hE81717E8)) lut_n59 (.I0(x21), .I1(x22), .I2(x23), .I3(n55), .I4(n56), .O(n59));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n60 (.I0(x30), .I1(x31), .I2(x32), .I3(n58), .I4(n59), .O(n60));
  LUT3 #(.INIT(8'h96)) lut_n61 (.I0(n47), .I1(n50), .I2(n53), .O(n61));
  LUT3 #(.INIT(8'hE8)) lut_n62 (.I0(n57), .I1(n60), .I2(n61), .O(n62));
  LUT3 #(.INIT(8'hE8)) lut_n63 (.I0(x36), .I1(x37), .I2(x38), .O(n63));
  LUT5 #(.INIT(32'hE81717E8)) lut_n64 (.I0(x30), .I1(x31), .I2(x32), .I3(n58), .I4(n59), .O(n64));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n65 (.I0(x33), .I1(x34), .I2(x35), .I3(n63), .I4(n64), .O(n65));
  LUT5 #(.INIT(32'hE81717E8)) lut_n66 (.I0(x33), .I1(x34), .I2(x35), .I3(n63), .I4(n64), .O(n66));
  LUT4 #(.INIT(16'hFFE8)) lut_n67 (.I0(x39), .I1(x40), .I2(x41), .I3(n66), .O(n67));
  LUT3 #(.INIT(8'h96)) lut_n68 (.I0(n57), .I1(n60), .I2(n61), .O(n68));
  LUT3 #(.INIT(8'hE8)) lut_n69 (.I0(n65), .I1(n67), .I2(n68), .O(n69));
  LUT3 #(.INIT(8'hE8)) lut_n70 (.I0(n54), .I1(n62), .I2(n69), .O(n70));
  LUT4 #(.INIT(16'h17E8)) lut_n71 (.I0(x39), .I1(x40), .I2(x41), .I3(n66), .O(n71));
  LUT3 #(.INIT(8'h96)) lut_n72 (.I0(n65), .I1(n67), .I2(n68), .O(n72));
  LUT2 #(.INIT(4'h2)) lut_n73 (.I0(n71), .I1(n72), .O(n73));
  LUT3 #(.INIT(8'h96)) lut_n74 (.I0(x0), .I1(x1), .I2(x2), .O(n74));
  LUT3 #(.INIT(8'h96)) lut_n75 (.I0(x6), .I1(x7), .I2(x8), .O(n75));
  LUT5 #(.INIT(32'hFF969600)) lut_n76 (.I0(x3), .I1(x4), .I2(x5), .I3(n74), .I4(n75), .O(n76));
  LUT3 #(.INIT(8'h96)) lut_n77 (.I0(x12), .I1(x13), .I2(x14), .O(n77));
  LUT5 #(.INIT(32'h96696996)) lut_n78 (.I0(x3), .I1(x4), .I2(x5), .I3(n74), .I4(n75), .O(n78));
  LUT5 #(.INIT(32'hFF969600)) lut_n79 (.I0(x9), .I1(x10), .I2(x11), .I3(n77), .I4(n78), .O(n79));
  LUT3 #(.INIT(8'hE8)) lut_n80 (.I0(n71), .I1(n76), .I2(n79), .O(n80));
  LUT2 #(.INIT(4'h6)) lut_n81 (.I0(n71), .I1(n72), .O(n81));
  LUT2 #(.INIT(4'h8)) lut_n82 (.I0(n80), .I1(n81), .O(n82));
  LUT3 #(.INIT(8'h96)) lut_n83 (.I0(n54), .I1(n62), .I2(n69), .O(n83));
  LUT3 #(.INIT(8'h96)) lut_n84 (.I0(x18), .I1(x19), .I2(x20), .O(n84));
  LUT5 #(.INIT(32'h96696996)) lut_n85 (.I0(x9), .I1(x10), .I2(x11), .I3(n77), .I4(n78), .O(n85));
  LUT5 #(.INIT(32'hFF969600)) lut_n86 (.I0(x15), .I1(x16), .I2(x17), .I3(n84), .I4(n85), .O(n86));
  LUT3 #(.INIT(8'h96)) lut_n87 (.I0(x24), .I1(x25), .I2(x26), .O(n87));
  LUT5 #(.INIT(32'h96696996)) lut_n88 (.I0(x15), .I1(x16), .I2(x17), .I3(n84), .I4(n85), .O(n88));
  LUT5 #(.INIT(32'hFF969600)) lut_n89 (.I0(x21), .I1(x22), .I2(x23), .I3(n87), .I4(n88), .O(n89));
  LUT3 #(.INIT(8'h96)) lut_n90 (.I0(n71), .I1(n76), .I2(n79), .O(n90));
  LUT3 #(.INIT(8'hE8)) lut_n91 (.I0(n86), .I1(n89), .I2(n90), .O(n91));
  LUT3 #(.INIT(8'h96)) lut_n92 (.I0(x27), .I1(x28), .I2(x29), .O(n92));
  LUT5 #(.INIT(32'h96696996)) lut_n93 (.I0(x21), .I1(x22), .I2(x23), .I3(n87), .I4(n88), .O(n93));
  LUT5 #(.INIT(32'hFF969600)) lut_n94 (.I0(x30), .I1(x31), .I2(x32), .I3(n92), .I4(n93), .O(n94));
  LUT3 #(.INIT(8'h96)) lut_n95 (.I0(x36), .I1(x37), .I2(x38), .O(n95));
  LUT5 #(.INIT(32'h96696996)) lut_n96 (.I0(x30), .I1(x31), .I2(x32), .I3(n92), .I4(n93), .O(n96));
  LUT5 #(.INIT(32'hFF969600)) lut_n97 (.I0(x33), .I1(x34), .I2(x35), .I3(n95), .I4(n96), .O(n97));
  LUT3 #(.INIT(8'h96)) lut_n98 (.I0(n86), .I1(n89), .I2(n90), .O(n98));
  LUT2 #(.INIT(4'h6)) lut_n99 (.I0(n80), .I1(n81), .O(n99));
  LUT5 #(.INIT(32'hFEEAA880)) lut_n100 (.I0(n91), .I1(n94), .I2(n97), .I3(n98), .I4(n99), .O(n100));
  LUT5 #(.INIT(32'h96696996)) lut_n101 (.I0(x33), .I1(x34), .I2(x35), .I3(n95), .I4(n96), .O(n101));
  LUT5 #(.INIT(32'hFF969600)) lut_n102 (.I0(x39), .I1(x40), .I2(x41), .I3(x42), .I4(n101), .O(n102));
  LUT6 #(.INIT(64'hA995566A81144228)) lut_n103 (.I0(n91), .I1(n94), .I2(n97), .I3(n98), .I4(n99), .I5(n102), .O(n103));
  LUT6 #(.INIT(64'hFBBABAA2BAA2A220)) lut_n104 (.I0(n70), .I1(n73), .I2(n82), .I3(n83), .I4(n100), .I5(n103), .O(n104));
  assign y0 = n104;
endmodule
