module top (x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255, x256, x257, x258, x259, x260, x261, x262, x263, x264, x265, x266, x267, x268, x269, x270, x271, x272, x273, x274, x275, x276, x277, x278, x279, x280, x281, x282, x283, x284, x285, x286, x287, x288, x289, x290, x291, x292, x293, x294, x295, x296, x297, x298, x299, x300, x301, x302, x303, x304, x305, x306, x307, x308, x309, x310, x311, x312, x313, x314, x315, x316, x317, x318, x319, x320, x321, x322, x323, x324, x325, x326, x327, x328, x329, x330, x331, x332, x333, x334, x335, x336, x337, x338, x339, x340, x341, x342, x343, x344, x345, x346, x347, x348, x349, x350, x351, x352, x353, x354, x355, x356, x357, x358, x359, x360, x361, x362, x363, x364, x365, x366, x367, x368, x369, x370, x371, x372, x373, x374, x375, x376, x377, x378, x379, x380, x381, x382, x383, x384, x385, x386, x387, x388, x389, x390, x391, x392, x393, x394, x395, x396, x397, x398, x399, x400, x401, x402, x403, x404, x405, x406, x407, x408, x409, x410, x411, x412, x413, x414, x415, x416, x417, x418, x419, x420, x421, x422, x423, x424, x425, x426, x427, x428, x429, x430, x431, x432, x433, x434, x435, x436, x437, x438, x439, x440, x441, x442, x443, x444, x445, x446, x447, x448, x449, x450, x451, x452, x453, x454, x455, x456, x457, x458, x459, x460, x461, x462, x463, x464, x465, x466, x467, x468, x469, x470, x471, x472, x473, x474, x475, x476, x477, x478, x479, x480, x481, x482, x483, x484, x485, x486, x487, x488, x489, x490, x491, x492, x493, x494, x495, x496, x497, x498, x499, x500, x501, x502, x503, x504, x505, x506, x507, x508, x509, x510, y0);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255, x256, x257, x258, x259, x260, x261, x262, x263, x264, x265, x266, x267, x268, x269, x270, x271, x272, x273, x274, x275, x276, x277, x278, x279, x280, x281, x282, x283, x284, x285, x286, x287, x288, x289, x290, x291, x292, x293, x294, x295, x296, x297, x298, x299, x300, x301, x302, x303, x304, x305, x306, x307, x308, x309, x310, x311, x312, x313, x314, x315, x316, x317, x318, x319, x320, x321, x322, x323, x324, x325, x326, x327, x328, x329, x330, x331, x332, x333, x334, x335, x336, x337, x338, x339, x340, x341, x342, x343, x344, x345, x346, x347, x348, x349, x350, x351, x352, x353, x354, x355, x356, x357, x358, x359, x360, x361, x362, x363, x364, x365, x366, x367, x368, x369, x370, x371, x372, x373, x374, x375, x376, x377, x378, x379, x380, x381, x382, x383, x384, x385, x386, x387, x388, x389, x390, x391, x392, x393, x394, x395, x396, x397, x398, x399, x400, x401, x402, x403, x404, x405, x406, x407, x408, x409, x410, x411, x412, x413, x414, x415, x416, x417, x418, x419, x420, x421, x422, x423, x424, x425, x426, x427, x428, x429, x430, x431, x432, x433, x434, x435, x436, x437, x438, x439, x440, x441, x442, x443, x444, x445, x446, x447, x448, x449, x450, x451, x452, x453, x454, x455, x456, x457, x458, x459, x460, x461, x462, x463, x464, x465, x466, x467, x468, x469, x470, x471, x472, x473, x474, x475, x476, x477, x478, x479, x480, x481, x482, x483, x484, x485, x486, x487, x488, x489, x490, x491, x492, x493, x494, x495, x496, x497, x498, x499, x500, x501, x502, x503, x504, x505, x506, x507, x508, x509, x510;
  output y0;
  wire n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328;
  LUT3 #(.INIT(8'hE8)) lut_n513 (.I0(x0), .I1(x1), .I2(x2), .O(n513));
  LUT3 #(.INIT(8'hE8)) lut_n514 (.I0(x6), .I1(x7), .I2(x8), .O(n514));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n515 (.I0(x3), .I1(x4), .I2(x5), .I3(n513), .I4(n514), .O(n515));
  LUT3 #(.INIT(8'hE8)) lut_n516 (.I0(x12), .I1(x13), .I2(x14), .O(n516));
  LUT5 #(.INIT(32'hE81717E8)) lut_n517 (.I0(x3), .I1(x4), .I2(x5), .I3(n513), .I4(n514), .O(n517));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n518 (.I0(x9), .I1(x10), .I2(x11), .I3(n516), .I4(n517), .O(n518));
  LUT3 #(.INIT(8'hE8)) lut_n519 (.I0(x18), .I1(x19), .I2(x20), .O(n519));
  LUT5 #(.INIT(32'hE81717E8)) lut_n520 (.I0(x9), .I1(x10), .I2(x11), .I3(n516), .I4(n517), .O(n520));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n521 (.I0(x15), .I1(x16), .I2(x17), .I3(n519), .I4(n520), .O(n521));
  LUT3 #(.INIT(8'hE8)) lut_n522 (.I0(n515), .I1(n518), .I2(n521), .O(n522));
  LUT3 #(.INIT(8'hE8)) lut_n523 (.I0(x24), .I1(x25), .I2(x26), .O(n523));
  LUT5 #(.INIT(32'hE81717E8)) lut_n524 (.I0(x15), .I1(x16), .I2(x17), .I3(n519), .I4(n520), .O(n524));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n525 (.I0(x21), .I1(x22), .I2(x23), .I3(n523), .I4(n524), .O(n525));
  LUT3 #(.INIT(8'hE8)) lut_n526 (.I0(x27), .I1(x28), .I2(x29), .O(n526));
  LUT5 #(.INIT(32'hE81717E8)) lut_n527 (.I0(x21), .I1(x22), .I2(x23), .I3(n523), .I4(n524), .O(n527));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n528 (.I0(x30), .I1(x31), .I2(x32), .I3(n526), .I4(n527), .O(n528));
  LUT3 #(.INIT(8'h96)) lut_n529 (.I0(n515), .I1(n518), .I2(n521), .O(n529));
  LUT3 #(.INIT(8'hE8)) lut_n530 (.I0(n525), .I1(n528), .I2(n529), .O(n530));
  LUT3 #(.INIT(8'hE8)) lut_n531 (.I0(x36), .I1(x37), .I2(x38), .O(n531));
  LUT5 #(.INIT(32'hE81717E8)) lut_n532 (.I0(x30), .I1(x31), .I2(x32), .I3(n526), .I4(n527), .O(n532));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n533 (.I0(x33), .I1(x34), .I2(x35), .I3(n531), .I4(n532), .O(n533));
  LUT3 #(.INIT(8'hE8)) lut_n534 (.I0(x42), .I1(x43), .I2(x44), .O(n534));
  LUT5 #(.INIT(32'hE81717E8)) lut_n535 (.I0(x33), .I1(x34), .I2(x35), .I3(n531), .I4(n532), .O(n535));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n536 (.I0(x39), .I1(x40), .I2(x41), .I3(n534), .I4(n535), .O(n536));
  LUT3 #(.INIT(8'h96)) lut_n537 (.I0(n525), .I1(n528), .I2(n529), .O(n537));
  LUT3 #(.INIT(8'hE8)) lut_n538 (.I0(n533), .I1(n536), .I2(n537), .O(n538));
  LUT3 #(.INIT(8'hE8)) lut_n539 (.I0(n522), .I1(n530), .I2(n538), .O(n539));
  LUT3 #(.INIT(8'hE8)) lut_n540 (.I0(x48), .I1(x49), .I2(x50), .O(n540));
  LUT5 #(.INIT(32'hE81717E8)) lut_n541 (.I0(x39), .I1(x40), .I2(x41), .I3(n534), .I4(n535), .O(n541));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n542 (.I0(x45), .I1(x46), .I2(x47), .I3(n540), .I4(n541), .O(n542));
  LUT3 #(.INIT(8'hE8)) lut_n543 (.I0(x54), .I1(x55), .I2(x56), .O(n543));
  LUT5 #(.INIT(32'hE81717E8)) lut_n544 (.I0(x45), .I1(x46), .I2(x47), .I3(n540), .I4(n541), .O(n544));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n545 (.I0(x51), .I1(x52), .I2(x53), .I3(n543), .I4(n544), .O(n545));
  LUT3 #(.INIT(8'h96)) lut_n546 (.I0(n533), .I1(n536), .I2(n537), .O(n546));
  LUT3 #(.INIT(8'hE8)) lut_n547 (.I0(n542), .I1(n545), .I2(n546), .O(n547));
  LUT3 #(.INIT(8'hE8)) lut_n548 (.I0(x60), .I1(x61), .I2(x62), .O(n548));
  LUT5 #(.INIT(32'hE81717E8)) lut_n549 (.I0(x51), .I1(x52), .I2(x53), .I3(n543), .I4(n544), .O(n549));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n550 (.I0(x57), .I1(x58), .I2(x59), .I3(n548), .I4(n549), .O(n550));
  LUT3 #(.INIT(8'hE8)) lut_n551 (.I0(x66), .I1(x67), .I2(x68), .O(n551));
  LUT5 #(.INIT(32'hE81717E8)) lut_n552 (.I0(x57), .I1(x58), .I2(x59), .I3(n548), .I4(n549), .O(n552));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n553 (.I0(x63), .I1(x64), .I2(x65), .I3(n551), .I4(n552), .O(n553));
  LUT3 #(.INIT(8'h96)) lut_n554 (.I0(n542), .I1(n545), .I2(n546), .O(n554));
  LUT3 #(.INIT(8'hE8)) lut_n555 (.I0(n550), .I1(n553), .I2(n554), .O(n555));
  LUT3 #(.INIT(8'h96)) lut_n556 (.I0(n522), .I1(n530), .I2(n538), .O(n556));
  LUT3 #(.INIT(8'hE8)) lut_n557 (.I0(n547), .I1(n555), .I2(n556), .O(n557));
  LUT3 #(.INIT(8'hE8)) lut_n558 (.I0(x72), .I1(x73), .I2(x74), .O(n558));
  LUT5 #(.INIT(32'hE81717E8)) lut_n559 (.I0(x63), .I1(x64), .I2(x65), .I3(n551), .I4(n552), .O(n559));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n560 (.I0(x69), .I1(x70), .I2(x71), .I3(n558), .I4(n559), .O(n560));
  LUT3 #(.INIT(8'hE8)) lut_n561 (.I0(x78), .I1(x79), .I2(x80), .O(n561));
  LUT5 #(.INIT(32'hE81717E8)) lut_n562 (.I0(x69), .I1(x70), .I2(x71), .I3(n558), .I4(n559), .O(n562));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n563 (.I0(x75), .I1(x76), .I2(x77), .I3(n561), .I4(n562), .O(n563));
  LUT3 #(.INIT(8'h96)) lut_n564 (.I0(n550), .I1(n553), .I2(n554), .O(n564));
  LUT3 #(.INIT(8'hE8)) lut_n565 (.I0(n560), .I1(n563), .I2(n564), .O(n565));
  LUT3 #(.INIT(8'hE8)) lut_n566 (.I0(x84), .I1(x85), .I2(x86), .O(n566));
  LUT5 #(.INIT(32'hE81717E8)) lut_n567 (.I0(x75), .I1(x76), .I2(x77), .I3(n561), .I4(n562), .O(n567));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n568 (.I0(x81), .I1(x82), .I2(x83), .I3(n566), .I4(n567), .O(n568));
  LUT3 #(.INIT(8'hE8)) lut_n569 (.I0(x90), .I1(x91), .I2(x92), .O(n569));
  LUT5 #(.INIT(32'hE81717E8)) lut_n570 (.I0(x81), .I1(x82), .I2(x83), .I3(n566), .I4(n567), .O(n570));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n571 (.I0(x87), .I1(x88), .I2(x89), .I3(n569), .I4(n570), .O(n571));
  LUT3 #(.INIT(8'h96)) lut_n572 (.I0(n560), .I1(n563), .I2(n564), .O(n572));
  LUT3 #(.INIT(8'hE8)) lut_n573 (.I0(n568), .I1(n571), .I2(n572), .O(n573));
  LUT3 #(.INIT(8'h96)) lut_n574 (.I0(n547), .I1(n555), .I2(n556), .O(n574));
  LUT3 #(.INIT(8'hE8)) lut_n575 (.I0(n565), .I1(n573), .I2(n574), .O(n575));
  LUT3 #(.INIT(8'hE8)) lut_n576 (.I0(n539), .I1(n557), .I2(n575), .O(n576));
  LUT3 #(.INIT(8'hE8)) lut_n577 (.I0(x96), .I1(x97), .I2(x98), .O(n577));
  LUT5 #(.INIT(32'hE81717E8)) lut_n578 (.I0(x87), .I1(x88), .I2(x89), .I3(n569), .I4(n570), .O(n578));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n579 (.I0(x93), .I1(x94), .I2(x95), .I3(n577), .I4(n578), .O(n579));
  LUT3 #(.INIT(8'hE8)) lut_n580 (.I0(x102), .I1(x103), .I2(x104), .O(n580));
  LUT5 #(.INIT(32'hE81717E8)) lut_n581 (.I0(x93), .I1(x94), .I2(x95), .I3(n577), .I4(n578), .O(n581));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n582 (.I0(x99), .I1(x100), .I2(x101), .I3(n580), .I4(n581), .O(n582));
  LUT3 #(.INIT(8'h96)) lut_n583 (.I0(n568), .I1(n571), .I2(n572), .O(n583));
  LUT3 #(.INIT(8'hE8)) lut_n584 (.I0(n579), .I1(n582), .I2(n583), .O(n584));
  LUT3 #(.INIT(8'hE8)) lut_n585 (.I0(x108), .I1(x109), .I2(x110), .O(n585));
  LUT5 #(.INIT(32'hE81717E8)) lut_n586 (.I0(x99), .I1(x100), .I2(x101), .I3(n580), .I4(n581), .O(n586));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n587 (.I0(x105), .I1(x106), .I2(x107), .I3(n585), .I4(n586), .O(n587));
  LUT3 #(.INIT(8'hE8)) lut_n588 (.I0(x114), .I1(x115), .I2(x116), .O(n588));
  LUT5 #(.INIT(32'hE81717E8)) lut_n589 (.I0(x105), .I1(x106), .I2(x107), .I3(n585), .I4(n586), .O(n589));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n590 (.I0(x111), .I1(x112), .I2(x113), .I3(n588), .I4(n589), .O(n590));
  LUT3 #(.INIT(8'h96)) lut_n591 (.I0(n579), .I1(n582), .I2(n583), .O(n591));
  LUT3 #(.INIT(8'hE8)) lut_n592 (.I0(n587), .I1(n590), .I2(n591), .O(n592));
  LUT3 #(.INIT(8'h96)) lut_n593 (.I0(n565), .I1(n573), .I2(n574), .O(n593));
  LUT3 #(.INIT(8'hE8)) lut_n594 (.I0(n584), .I1(n592), .I2(n593), .O(n594));
  LUT3 #(.INIT(8'hE8)) lut_n595 (.I0(x120), .I1(x121), .I2(x122), .O(n595));
  LUT5 #(.INIT(32'hE81717E8)) lut_n596 (.I0(x111), .I1(x112), .I2(x113), .I3(n588), .I4(n589), .O(n596));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n597 (.I0(x117), .I1(x118), .I2(x119), .I3(n595), .I4(n596), .O(n597));
  LUT3 #(.INIT(8'hE8)) lut_n598 (.I0(x126), .I1(x127), .I2(x128), .O(n598));
  LUT5 #(.INIT(32'hE81717E8)) lut_n599 (.I0(x117), .I1(x118), .I2(x119), .I3(n595), .I4(n596), .O(n599));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n600 (.I0(x123), .I1(x124), .I2(x125), .I3(n598), .I4(n599), .O(n600));
  LUT3 #(.INIT(8'h96)) lut_n601 (.I0(n587), .I1(n590), .I2(n591), .O(n601));
  LUT3 #(.INIT(8'hE8)) lut_n602 (.I0(n597), .I1(n600), .I2(n601), .O(n602));
  LUT3 #(.INIT(8'hE8)) lut_n603 (.I0(x132), .I1(x133), .I2(x134), .O(n603));
  LUT5 #(.INIT(32'hE81717E8)) lut_n604 (.I0(x123), .I1(x124), .I2(x125), .I3(n598), .I4(n599), .O(n604));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n605 (.I0(x129), .I1(x130), .I2(x131), .I3(n603), .I4(n604), .O(n605));
  LUT3 #(.INIT(8'hE8)) lut_n606 (.I0(x138), .I1(x139), .I2(x140), .O(n606));
  LUT5 #(.INIT(32'hE81717E8)) lut_n607 (.I0(x129), .I1(x130), .I2(x131), .I3(n603), .I4(n604), .O(n607));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n608 (.I0(x135), .I1(x136), .I2(x137), .I3(n606), .I4(n607), .O(n608));
  LUT3 #(.INIT(8'h96)) lut_n609 (.I0(n597), .I1(n600), .I2(n601), .O(n609));
  LUT3 #(.INIT(8'hE8)) lut_n610 (.I0(n605), .I1(n608), .I2(n609), .O(n610));
  LUT3 #(.INIT(8'h96)) lut_n611 (.I0(n584), .I1(n592), .I2(n593), .O(n611));
  LUT3 #(.INIT(8'hE8)) lut_n612 (.I0(n602), .I1(n610), .I2(n611), .O(n612));
  LUT3 #(.INIT(8'h96)) lut_n613 (.I0(n539), .I1(n557), .I2(n575), .O(n613));
  LUT3 #(.INIT(8'hE8)) lut_n614 (.I0(n594), .I1(n612), .I2(n613), .O(n614));
  LUT3 #(.INIT(8'hE8)) lut_n615 (.I0(x144), .I1(x145), .I2(x146), .O(n615));
  LUT5 #(.INIT(32'hE81717E8)) lut_n616 (.I0(x135), .I1(x136), .I2(x137), .I3(n606), .I4(n607), .O(n616));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n617 (.I0(x141), .I1(x142), .I2(x143), .I3(n615), .I4(n616), .O(n617));
  LUT3 #(.INIT(8'hE8)) lut_n618 (.I0(x150), .I1(x151), .I2(x152), .O(n618));
  LUT5 #(.INIT(32'hE81717E8)) lut_n619 (.I0(x141), .I1(x142), .I2(x143), .I3(n615), .I4(n616), .O(n619));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n620 (.I0(x147), .I1(x148), .I2(x149), .I3(n618), .I4(n619), .O(n620));
  LUT3 #(.INIT(8'h96)) lut_n621 (.I0(n605), .I1(n608), .I2(n609), .O(n621));
  LUT3 #(.INIT(8'hE8)) lut_n622 (.I0(n617), .I1(n620), .I2(n621), .O(n622));
  LUT3 #(.INIT(8'hE8)) lut_n623 (.I0(x156), .I1(x157), .I2(x158), .O(n623));
  LUT5 #(.INIT(32'hE81717E8)) lut_n624 (.I0(x147), .I1(x148), .I2(x149), .I3(n618), .I4(n619), .O(n624));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n625 (.I0(x153), .I1(x154), .I2(x155), .I3(n623), .I4(n624), .O(n625));
  LUT3 #(.INIT(8'hE8)) lut_n626 (.I0(x162), .I1(x163), .I2(x164), .O(n626));
  LUT5 #(.INIT(32'hE81717E8)) lut_n627 (.I0(x153), .I1(x154), .I2(x155), .I3(n623), .I4(n624), .O(n627));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n628 (.I0(x159), .I1(x160), .I2(x161), .I3(n626), .I4(n627), .O(n628));
  LUT3 #(.INIT(8'h96)) lut_n629 (.I0(n617), .I1(n620), .I2(n621), .O(n629));
  LUT3 #(.INIT(8'hE8)) lut_n630 (.I0(n625), .I1(n628), .I2(n629), .O(n630));
  LUT3 #(.INIT(8'h96)) lut_n631 (.I0(n602), .I1(n610), .I2(n611), .O(n631));
  LUT3 #(.INIT(8'hE8)) lut_n632 (.I0(n622), .I1(n630), .I2(n631), .O(n632));
  LUT3 #(.INIT(8'hE8)) lut_n633 (.I0(x168), .I1(x169), .I2(x170), .O(n633));
  LUT5 #(.INIT(32'hE81717E8)) lut_n634 (.I0(x159), .I1(x160), .I2(x161), .I3(n626), .I4(n627), .O(n634));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n635 (.I0(x165), .I1(x166), .I2(x167), .I3(n633), .I4(n634), .O(n635));
  LUT3 #(.INIT(8'hE8)) lut_n636 (.I0(x174), .I1(x175), .I2(x176), .O(n636));
  LUT5 #(.INIT(32'hE81717E8)) lut_n637 (.I0(x165), .I1(x166), .I2(x167), .I3(n633), .I4(n634), .O(n637));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n638 (.I0(x171), .I1(x172), .I2(x173), .I3(n636), .I4(n637), .O(n638));
  LUT3 #(.INIT(8'h96)) lut_n639 (.I0(n625), .I1(n628), .I2(n629), .O(n639));
  LUT3 #(.INIT(8'hE8)) lut_n640 (.I0(n635), .I1(n638), .I2(n639), .O(n640));
  LUT3 #(.INIT(8'hE8)) lut_n641 (.I0(x180), .I1(x181), .I2(x182), .O(n641));
  LUT5 #(.INIT(32'hE81717E8)) lut_n642 (.I0(x171), .I1(x172), .I2(x173), .I3(n636), .I4(n637), .O(n642));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n643 (.I0(x177), .I1(x178), .I2(x179), .I3(n641), .I4(n642), .O(n643));
  LUT3 #(.INIT(8'hE8)) lut_n644 (.I0(x186), .I1(x187), .I2(x188), .O(n644));
  LUT5 #(.INIT(32'hE81717E8)) lut_n645 (.I0(x177), .I1(x178), .I2(x179), .I3(n641), .I4(n642), .O(n645));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n646 (.I0(x183), .I1(x184), .I2(x185), .I3(n644), .I4(n645), .O(n646));
  LUT3 #(.INIT(8'h96)) lut_n647 (.I0(n635), .I1(n638), .I2(n639), .O(n647));
  LUT3 #(.INIT(8'hE8)) lut_n648 (.I0(n643), .I1(n646), .I2(n647), .O(n648));
  LUT3 #(.INIT(8'h96)) lut_n649 (.I0(n622), .I1(n630), .I2(n631), .O(n649));
  LUT3 #(.INIT(8'hE8)) lut_n650 (.I0(n640), .I1(n648), .I2(n649), .O(n650));
  LUT3 #(.INIT(8'h96)) lut_n651 (.I0(n594), .I1(n612), .I2(n613), .O(n651));
  LUT3 #(.INIT(8'hE8)) lut_n652 (.I0(n632), .I1(n650), .I2(n651), .O(n652));
  LUT3 #(.INIT(8'hE8)) lut_n653 (.I0(n576), .I1(n614), .I2(n652), .O(n653));
  LUT3 #(.INIT(8'hE8)) lut_n654 (.I0(x192), .I1(x193), .I2(x194), .O(n654));
  LUT5 #(.INIT(32'hE81717E8)) lut_n655 (.I0(x183), .I1(x184), .I2(x185), .I3(n644), .I4(n645), .O(n655));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n656 (.I0(x189), .I1(x190), .I2(x191), .I3(n654), .I4(n655), .O(n656));
  LUT3 #(.INIT(8'hE8)) lut_n657 (.I0(x198), .I1(x199), .I2(x200), .O(n657));
  LUT5 #(.INIT(32'hE81717E8)) lut_n658 (.I0(x189), .I1(x190), .I2(x191), .I3(n654), .I4(n655), .O(n658));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n659 (.I0(x195), .I1(x196), .I2(x197), .I3(n657), .I4(n658), .O(n659));
  LUT3 #(.INIT(8'h96)) lut_n660 (.I0(n643), .I1(n646), .I2(n647), .O(n660));
  LUT3 #(.INIT(8'hE8)) lut_n661 (.I0(n656), .I1(n659), .I2(n660), .O(n661));
  LUT3 #(.INIT(8'hE8)) lut_n662 (.I0(x204), .I1(x205), .I2(x206), .O(n662));
  LUT5 #(.INIT(32'hE81717E8)) lut_n663 (.I0(x195), .I1(x196), .I2(x197), .I3(n657), .I4(n658), .O(n663));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n664 (.I0(x201), .I1(x202), .I2(x203), .I3(n662), .I4(n663), .O(n664));
  LUT3 #(.INIT(8'hE8)) lut_n665 (.I0(x210), .I1(x211), .I2(x212), .O(n665));
  LUT5 #(.INIT(32'hE81717E8)) lut_n666 (.I0(x201), .I1(x202), .I2(x203), .I3(n662), .I4(n663), .O(n666));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n667 (.I0(x207), .I1(x208), .I2(x209), .I3(n665), .I4(n666), .O(n667));
  LUT3 #(.INIT(8'h96)) lut_n668 (.I0(n656), .I1(n659), .I2(n660), .O(n668));
  LUT3 #(.INIT(8'hE8)) lut_n669 (.I0(n664), .I1(n667), .I2(n668), .O(n669));
  LUT3 #(.INIT(8'h96)) lut_n670 (.I0(n640), .I1(n648), .I2(n649), .O(n670));
  LUT3 #(.INIT(8'hE8)) lut_n671 (.I0(n661), .I1(n669), .I2(n670), .O(n671));
  LUT3 #(.INIT(8'hE8)) lut_n672 (.I0(x216), .I1(x217), .I2(x218), .O(n672));
  LUT5 #(.INIT(32'hE81717E8)) lut_n673 (.I0(x207), .I1(x208), .I2(x209), .I3(n665), .I4(n666), .O(n673));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n674 (.I0(x213), .I1(x214), .I2(x215), .I3(n672), .I4(n673), .O(n674));
  LUT3 #(.INIT(8'hE8)) lut_n675 (.I0(x222), .I1(x223), .I2(x224), .O(n675));
  LUT5 #(.INIT(32'hE81717E8)) lut_n676 (.I0(x213), .I1(x214), .I2(x215), .I3(n672), .I4(n673), .O(n676));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n677 (.I0(x219), .I1(x220), .I2(x221), .I3(n675), .I4(n676), .O(n677));
  LUT3 #(.INIT(8'h96)) lut_n678 (.I0(n664), .I1(n667), .I2(n668), .O(n678));
  LUT3 #(.INIT(8'hE8)) lut_n679 (.I0(n674), .I1(n677), .I2(n678), .O(n679));
  LUT3 #(.INIT(8'hE8)) lut_n680 (.I0(x228), .I1(x229), .I2(x230), .O(n680));
  LUT5 #(.INIT(32'hE81717E8)) lut_n681 (.I0(x219), .I1(x220), .I2(x221), .I3(n675), .I4(n676), .O(n681));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n682 (.I0(x225), .I1(x226), .I2(x227), .I3(n680), .I4(n681), .O(n682));
  LUT3 #(.INIT(8'hE8)) lut_n683 (.I0(x234), .I1(x235), .I2(x236), .O(n683));
  LUT5 #(.INIT(32'hE81717E8)) lut_n684 (.I0(x225), .I1(x226), .I2(x227), .I3(n680), .I4(n681), .O(n684));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n685 (.I0(x231), .I1(x232), .I2(x233), .I3(n683), .I4(n684), .O(n685));
  LUT3 #(.INIT(8'h96)) lut_n686 (.I0(n674), .I1(n677), .I2(n678), .O(n686));
  LUT3 #(.INIT(8'hE8)) lut_n687 (.I0(n682), .I1(n685), .I2(n686), .O(n687));
  LUT3 #(.INIT(8'h96)) lut_n688 (.I0(n661), .I1(n669), .I2(n670), .O(n688));
  LUT3 #(.INIT(8'hE8)) lut_n689 (.I0(n679), .I1(n687), .I2(n688), .O(n689));
  LUT3 #(.INIT(8'h96)) lut_n690 (.I0(n632), .I1(n650), .I2(n651), .O(n690));
  LUT3 #(.INIT(8'hE8)) lut_n691 (.I0(n671), .I1(n689), .I2(n690), .O(n691));
  LUT3 #(.INIT(8'hE8)) lut_n692 (.I0(x240), .I1(x241), .I2(x242), .O(n692));
  LUT5 #(.INIT(32'hE81717E8)) lut_n693 (.I0(x231), .I1(x232), .I2(x233), .I3(n683), .I4(n684), .O(n693));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n694 (.I0(x237), .I1(x238), .I2(x239), .I3(n692), .I4(n693), .O(n694));
  LUT3 #(.INIT(8'hE8)) lut_n695 (.I0(x246), .I1(x247), .I2(x248), .O(n695));
  LUT5 #(.INIT(32'hE81717E8)) lut_n696 (.I0(x237), .I1(x238), .I2(x239), .I3(n692), .I4(n693), .O(n696));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n697 (.I0(x243), .I1(x244), .I2(x245), .I3(n695), .I4(n696), .O(n697));
  LUT3 #(.INIT(8'h96)) lut_n698 (.I0(n682), .I1(n685), .I2(n686), .O(n698));
  LUT3 #(.INIT(8'hE8)) lut_n699 (.I0(n694), .I1(n697), .I2(n698), .O(n699));
  LUT3 #(.INIT(8'hE8)) lut_n700 (.I0(x252), .I1(x253), .I2(x254), .O(n700));
  LUT5 #(.INIT(32'hE81717E8)) lut_n701 (.I0(x243), .I1(x244), .I2(x245), .I3(n695), .I4(n696), .O(n701));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n702 (.I0(x249), .I1(x250), .I2(x251), .I3(n700), .I4(n701), .O(n702));
  LUT3 #(.INIT(8'hE8)) lut_n703 (.I0(x258), .I1(x259), .I2(x260), .O(n703));
  LUT5 #(.INIT(32'hE81717E8)) lut_n704 (.I0(x249), .I1(x250), .I2(x251), .I3(n700), .I4(n701), .O(n704));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n705 (.I0(x255), .I1(x256), .I2(x257), .I3(n703), .I4(n704), .O(n705));
  LUT3 #(.INIT(8'h96)) lut_n706 (.I0(n694), .I1(n697), .I2(n698), .O(n706));
  LUT3 #(.INIT(8'hE8)) lut_n707 (.I0(n702), .I1(n705), .I2(n706), .O(n707));
  LUT3 #(.INIT(8'h96)) lut_n708 (.I0(n679), .I1(n687), .I2(n688), .O(n708));
  LUT3 #(.INIT(8'hE8)) lut_n709 (.I0(n699), .I1(n707), .I2(n708), .O(n709));
  LUT3 #(.INIT(8'hE8)) lut_n710 (.I0(x264), .I1(x265), .I2(x266), .O(n710));
  LUT5 #(.INIT(32'hE81717E8)) lut_n711 (.I0(x255), .I1(x256), .I2(x257), .I3(n703), .I4(n704), .O(n711));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n712 (.I0(x261), .I1(x262), .I2(x263), .I3(n710), .I4(n711), .O(n712));
  LUT3 #(.INIT(8'hE8)) lut_n713 (.I0(x270), .I1(x271), .I2(x272), .O(n713));
  LUT5 #(.INIT(32'hE81717E8)) lut_n714 (.I0(x261), .I1(x262), .I2(x263), .I3(n710), .I4(n711), .O(n714));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n715 (.I0(x267), .I1(x268), .I2(x269), .I3(n713), .I4(n714), .O(n715));
  LUT3 #(.INIT(8'h96)) lut_n716 (.I0(n702), .I1(n705), .I2(n706), .O(n716));
  LUT3 #(.INIT(8'hE8)) lut_n717 (.I0(n712), .I1(n715), .I2(n716), .O(n717));
  LUT3 #(.INIT(8'hE8)) lut_n718 (.I0(x276), .I1(x277), .I2(x278), .O(n718));
  LUT5 #(.INIT(32'hE81717E8)) lut_n719 (.I0(x267), .I1(x268), .I2(x269), .I3(n713), .I4(n714), .O(n719));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n720 (.I0(x273), .I1(x274), .I2(x275), .I3(n718), .I4(n719), .O(n720));
  LUT3 #(.INIT(8'hE8)) lut_n721 (.I0(x282), .I1(x283), .I2(x284), .O(n721));
  LUT5 #(.INIT(32'hE81717E8)) lut_n722 (.I0(x273), .I1(x274), .I2(x275), .I3(n718), .I4(n719), .O(n722));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n723 (.I0(x279), .I1(x280), .I2(x281), .I3(n721), .I4(n722), .O(n723));
  LUT3 #(.INIT(8'h96)) lut_n724 (.I0(n712), .I1(n715), .I2(n716), .O(n724));
  LUT3 #(.INIT(8'hE8)) lut_n725 (.I0(n720), .I1(n723), .I2(n724), .O(n725));
  LUT3 #(.INIT(8'h96)) lut_n726 (.I0(n699), .I1(n707), .I2(n708), .O(n726));
  LUT3 #(.INIT(8'hE8)) lut_n727 (.I0(n717), .I1(n725), .I2(n726), .O(n727));
  LUT3 #(.INIT(8'h96)) lut_n728 (.I0(n671), .I1(n689), .I2(n690), .O(n728));
  LUT3 #(.INIT(8'hE8)) lut_n729 (.I0(n709), .I1(n727), .I2(n728), .O(n729));
  LUT3 #(.INIT(8'h96)) lut_n730 (.I0(n576), .I1(n614), .I2(n652), .O(n730));
  LUT3 #(.INIT(8'hE8)) lut_n731 (.I0(n691), .I1(n729), .I2(n730), .O(n731));
  LUT3 #(.INIT(8'hE8)) lut_n732 (.I0(x288), .I1(x289), .I2(x290), .O(n732));
  LUT5 #(.INIT(32'hE81717E8)) lut_n733 (.I0(x279), .I1(x280), .I2(x281), .I3(n721), .I4(n722), .O(n733));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n734 (.I0(x285), .I1(x286), .I2(x287), .I3(n732), .I4(n733), .O(n734));
  LUT3 #(.INIT(8'hE8)) lut_n735 (.I0(x294), .I1(x295), .I2(x296), .O(n735));
  LUT5 #(.INIT(32'hE81717E8)) lut_n736 (.I0(x285), .I1(x286), .I2(x287), .I3(n732), .I4(n733), .O(n736));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n737 (.I0(x291), .I1(x292), .I2(x293), .I3(n735), .I4(n736), .O(n737));
  LUT3 #(.INIT(8'h96)) lut_n738 (.I0(n720), .I1(n723), .I2(n724), .O(n738));
  LUT3 #(.INIT(8'hE8)) lut_n739 (.I0(n734), .I1(n737), .I2(n738), .O(n739));
  LUT3 #(.INIT(8'hE8)) lut_n740 (.I0(x297), .I1(x298), .I2(x299), .O(n740));
  LUT5 #(.INIT(32'hE81717E8)) lut_n741 (.I0(x291), .I1(x292), .I2(x293), .I3(n735), .I4(n736), .O(n741));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n742 (.I0(x300), .I1(x301), .I2(x302), .I3(n740), .I4(n741), .O(n742));
  LUT3 #(.INIT(8'hE8)) lut_n743 (.I0(x306), .I1(x307), .I2(x308), .O(n743));
  LUT5 #(.INIT(32'hE81717E8)) lut_n744 (.I0(x300), .I1(x301), .I2(x302), .I3(n740), .I4(n741), .O(n744));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n745 (.I0(x303), .I1(x304), .I2(x305), .I3(n743), .I4(n744), .O(n745));
  LUT3 #(.INIT(8'h96)) lut_n746 (.I0(n734), .I1(n737), .I2(n738), .O(n746));
  LUT3 #(.INIT(8'hE8)) lut_n747 (.I0(n742), .I1(n745), .I2(n746), .O(n747));
  LUT3 #(.INIT(8'h96)) lut_n748 (.I0(n717), .I1(n725), .I2(n726), .O(n748));
  LUT3 #(.INIT(8'hE8)) lut_n749 (.I0(n739), .I1(n747), .I2(n748), .O(n749));
  LUT3 #(.INIT(8'hE8)) lut_n750 (.I0(x312), .I1(x313), .I2(x314), .O(n750));
  LUT5 #(.INIT(32'hE81717E8)) lut_n751 (.I0(x303), .I1(x304), .I2(x305), .I3(n743), .I4(n744), .O(n751));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n752 (.I0(x309), .I1(x310), .I2(x311), .I3(n750), .I4(n751), .O(n752));
  LUT3 #(.INIT(8'hE8)) lut_n753 (.I0(x318), .I1(x319), .I2(x320), .O(n753));
  LUT5 #(.INIT(32'hE81717E8)) lut_n754 (.I0(x309), .I1(x310), .I2(x311), .I3(n750), .I4(n751), .O(n754));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n755 (.I0(x315), .I1(x316), .I2(x317), .I3(n753), .I4(n754), .O(n755));
  LUT3 #(.INIT(8'h96)) lut_n756 (.I0(n742), .I1(n745), .I2(n746), .O(n756));
  LUT3 #(.INIT(8'hE8)) lut_n757 (.I0(n752), .I1(n755), .I2(n756), .O(n757));
  LUT3 #(.INIT(8'hE8)) lut_n758 (.I0(x324), .I1(x325), .I2(x326), .O(n758));
  LUT5 #(.INIT(32'hE81717E8)) lut_n759 (.I0(x315), .I1(x316), .I2(x317), .I3(n753), .I4(n754), .O(n759));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n760 (.I0(x321), .I1(x322), .I2(x323), .I3(n758), .I4(n759), .O(n760));
  LUT3 #(.INIT(8'hE8)) lut_n761 (.I0(x330), .I1(x331), .I2(x332), .O(n761));
  LUT5 #(.INIT(32'hE81717E8)) lut_n762 (.I0(x321), .I1(x322), .I2(x323), .I3(n758), .I4(n759), .O(n762));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n763 (.I0(x327), .I1(x328), .I2(x329), .I3(n761), .I4(n762), .O(n763));
  LUT3 #(.INIT(8'h96)) lut_n764 (.I0(n752), .I1(n755), .I2(n756), .O(n764));
  LUT3 #(.INIT(8'hE8)) lut_n765 (.I0(n760), .I1(n763), .I2(n764), .O(n765));
  LUT3 #(.INIT(8'h96)) lut_n766 (.I0(n739), .I1(n747), .I2(n748), .O(n766));
  LUT3 #(.INIT(8'hE8)) lut_n767 (.I0(n757), .I1(n765), .I2(n766), .O(n767));
  LUT3 #(.INIT(8'h96)) lut_n768 (.I0(n709), .I1(n727), .I2(n728), .O(n768));
  LUT3 #(.INIT(8'hE8)) lut_n769 (.I0(n749), .I1(n767), .I2(n768), .O(n769));
  LUT3 #(.INIT(8'hE8)) lut_n770 (.I0(x336), .I1(x337), .I2(x338), .O(n770));
  LUT5 #(.INIT(32'hE81717E8)) lut_n771 (.I0(x327), .I1(x328), .I2(x329), .I3(n761), .I4(n762), .O(n771));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n772 (.I0(x333), .I1(x334), .I2(x335), .I3(n770), .I4(n771), .O(n772));
  LUT3 #(.INIT(8'hE8)) lut_n773 (.I0(x342), .I1(x343), .I2(x344), .O(n773));
  LUT5 #(.INIT(32'hE81717E8)) lut_n774 (.I0(x333), .I1(x334), .I2(x335), .I3(n770), .I4(n771), .O(n774));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n775 (.I0(x339), .I1(x340), .I2(x341), .I3(n773), .I4(n774), .O(n775));
  LUT3 #(.INIT(8'h96)) lut_n776 (.I0(n760), .I1(n763), .I2(n764), .O(n776));
  LUT3 #(.INIT(8'hE8)) lut_n777 (.I0(n772), .I1(n775), .I2(n776), .O(n777));
  LUT3 #(.INIT(8'hE8)) lut_n778 (.I0(x348), .I1(x349), .I2(x350), .O(n778));
  LUT5 #(.INIT(32'hE81717E8)) lut_n779 (.I0(x339), .I1(x340), .I2(x341), .I3(n773), .I4(n774), .O(n779));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n780 (.I0(x345), .I1(x346), .I2(x347), .I3(n778), .I4(n779), .O(n780));
  LUT3 #(.INIT(8'hE8)) lut_n781 (.I0(x354), .I1(x355), .I2(x356), .O(n781));
  LUT5 #(.INIT(32'hE81717E8)) lut_n782 (.I0(x345), .I1(x346), .I2(x347), .I3(n778), .I4(n779), .O(n782));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n783 (.I0(x351), .I1(x352), .I2(x353), .I3(n781), .I4(n782), .O(n783));
  LUT3 #(.INIT(8'h96)) lut_n784 (.I0(n772), .I1(n775), .I2(n776), .O(n784));
  LUT3 #(.INIT(8'hE8)) lut_n785 (.I0(n780), .I1(n783), .I2(n784), .O(n785));
  LUT3 #(.INIT(8'h96)) lut_n786 (.I0(n757), .I1(n765), .I2(n766), .O(n786));
  LUT3 #(.INIT(8'hE8)) lut_n787 (.I0(n777), .I1(n785), .I2(n786), .O(n787));
  LUT3 #(.INIT(8'hE8)) lut_n788 (.I0(x360), .I1(x361), .I2(x362), .O(n788));
  LUT5 #(.INIT(32'hE81717E8)) lut_n789 (.I0(x351), .I1(x352), .I2(x353), .I3(n781), .I4(n782), .O(n789));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n790 (.I0(x357), .I1(x358), .I2(x359), .I3(n788), .I4(n789), .O(n790));
  LUT3 #(.INIT(8'hE8)) lut_n791 (.I0(x366), .I1(x367), .I2(x368), .O(n791));
  LUT5 #(.INIT(32'hE81717E8)) lut_n792 (.I0(x357), .I1(x358), .I2(x359), .I3(n788), .I4(n789), .O(n792));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n793 (.I0(x363), .I1(x364), .I2(x365), .I3(n791), .I4(n792), .O(n793));
  LUT3 #(.INIT(8'h96)) lut_n794 (.I0(n780), .I1(n783), .I2(n784), .O(n794));
  LUT3 #(.INIT(8'hE8)) lut_n795 (.I0(n790), .I1(n793), .I2(n794), .O(n795));
  LUT3 #(.INIT(8'hE8)) lut_n796 (.I0(x372), .I1(x373), .I2(x374), .O(n796));
  LUT5 #(.INIT(32'hE81717E8)) lut_n797 (.I0(x363), .I1(x364), .I2(x365), .I3(n791), .I4(n792), .O(n797));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n798 (.I0(x369), .I1(x370), .I2(x371), .I3(n796), .I4(n797), .O(n798));
  LUT3 #(.INIT(8'hE8)) lut_n799 (.I0(x378), .I1(x379), .I2(x380), .O(n799));
  LUT5 #(.INIT(32'hE81717E8)) lut_n800 (.I0(x369), .I1(x370), .I2(x371), .I3(n796), .I4(n797), .O(n800));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n801 (.I0(x375), .I1(x376), .I2(x377), .I3(n799), .I4(n800), .O(n801));
  LUT3 #(.INIT(8'h96)) lut_n802 (.I0(n790), .I1(n793), .I2(n794), .O(n802));
  LUT3 #(.INIT(8'hE8)) lut_n803 (.I0(n798), .I1(n801), .I2(n802), .O(n803));
  LUT3 #(.INIT(8'h96)) lut_n804 (.I0(n777), .I1(n785), .I2(n786), .O(n804));
  LUT3 #(.INIT(8'hE8)) lut_n805 (.I0(n795), .I1(n803), .I2(n804), .O(n805));
  LUT3 #(.INIT(8'h96)) lut_n806 (.I0(n749), .I1(n767), .I2(n768), .O(n806));
  LUT3 #(.INIT(8'hE8)) lut_n807 (.I0(n787), .I1(n805), .I2(n806), .O(n807));
  LUT3 #(.INIT(8'h96)) lut_n808 (.I0(n691), .I1(n729), .I2(n730), .O(n808));
  LUT3 #(.INIT(8'hE8)) lut_n809 (.I0(n769), .I1(n807), .I2(n808), .O(n809));
  LUT3 #(.INIT(8'hE8)) lut_n810 (.I0(n653), .I1(n731), .I2(n809), .O(n810));
  LUT3 #(.INIT(8'hE8)) lut_n811 (.I0(x384), .I1(x385), .I2(x386), .O(n811));
  LUT5 #(.INIT(32'hE81717E8)) lut_n812 (.I0(x375), .I1(x376), .I2(x377), .I3(n799), .I4(n800), .O(n812));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n813 (.I0(x381), .I1(x382), .I2(x383), .I3(n811), .I4(n812), .O(n813));
  LUT3 #(.INIT(8'hE8)) lut_n814 (.I0(x390), .I1(x391), .I2(x392), .O(n814));
  LUT5 #(.INIT(32'hE81717E8)) lut_n815 (.I0(x381), .I1(x382), .I2(x383), .I3(n811), .I4(n812), .O(n815));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n816 (.I0(x387), .I1(x388), .I2(x389), .I3(n814), .I4(n815), .O(n816));
  LUT3 #(.INIT(8'h96)) lut_n817 (.I0(n798), .I1(n801), .I2(n802), .O(n817));
  LUT3 #(.INIT(8'hE8)) lut_n818 (.I0(n813), .I1(n816), .I2(n817), .O(n818));
  LUT3 #(.INIT(8'hE8)) lut_n819 (.I0(x396), .I1(x397), .I2(x398), .O(n819));
  LUT5 #(.INIT(32'hE81717E8)) lut_n820 (.I0(x387), .I1(x388), .I2(x389), .I3(n814), .I4(n815), .O(n820));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n821 (.I0(x393), .I1(x394), .I2(x395), .I3(n819), .I4(n820), .O(n821));
  LUT3 #(.INIT(8'hE8)) lut_n822 (.I0(x402), .I1(x403), .I2(x404), .O(n822));
  LUT5 #(.INIT(32'hE81717E8)) lut_n823 (.I0(x393), .I1(x394), .I2(x395), .I3(n819), .I4(n820), .O(n823));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n824 (.I0(x399), .I1(x400), .I2(x401), .I3(n822), .I4(n823), .O(n824));
  LUT3 #(.INIT(8'h96)) lut_n825 (.I0(n813), .I1(n816), .I2(n817), .O(n825));
  LUT3 #(.INIT(8'hE8)) lut_n826 (.I0(n821), .I1(n824), .I2(n825), .O(n826));
  LUT3 #(.INIT(8'h96)) lut_n827 (.I0(n795), .I1(n803), .I2(n804), .O(n827));
  LUT3 #(.INIT(8'hE8)) lut_n828 (.I0(n818), .I1(n826), .I2(n827), .O(n828));
  LUT3 #(.INIT(8'hE8)) lut_n829 (.I0(x408), .I1(x409), .I2(x410), .O(n829));
  LUT5 #(.INIT(32'hE81717E8)) lut_n830 (.I0(x399), .I1(x400), .I2(x401), .I3(n822), .I4(n823), .O(n830));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n831 (.I0(x405), .I1(x406), .I2(x407), .I3(n829), .I4(n830), .O(n831));
  LUT3 #(.INIT(8'hE8)) lut_n832 (.I0(x414), .I1(x415), .I2(x416), .O(n832));
  LUT5 #(.INIT(32'hE81717E8)) lut_n833 (.I0(x405), .I1(x406), .I2(x407), .I3(n829), .I4(n830), .O(n833));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n834 (.I0(x411), .I1(x412), .I2(x413), .I3(n832), .I4(n833), .O(n834));
  LUT3 #(.INIT(8'h96)) lut_n835 (.I0(n821), .I1(n824), .I2(n825), .O(n835));
  LUT3 #(.INIT(8'hE8)) lut_n836 (.I0(n831), .I1(n834), .I2(n835), .O(n836));
  LUT3 #(.INIT(8'hE8)) lut_n837 (.I0(x420), .I1(x421), .I2(x422), .O(n837));
  LUT5 #(.INIT(32'hE81717E8)) lut_n838 (.I0(x411), .I1(x412), .I2(x413), .I3(n832), .I4(n833), .O(n838));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n839 (.I0(x417), .I1(x418), .I2(x419), .I3(n837), .I4(n838), .O(n839));
  LUT3 #(.INIT(8'hE8)) lut_n840 (.I0(x426), .I1(x427), .I2(x428), .O(n840));
  LUT5 #(.INIT(32'hE81717E8)) lut_n841 (.I0(x417), .I1(x418), .I2(x419), .I3(n837), .I4(n838), .O(n841));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n842 (.I0(x423), .I1(x424), .I2(x425), .I3(n840), .I4(n841), .O(n842));
  LUT3 #(.INIT(8'h96)) lut_n843 (.I0(n831), .I1(n834), .I2(n835), .O(n843));
  LUT3 #(.INIT(8'hE8)) lut_n844 (.I0(n839), .I1(n842), .I2(n843), .O(n844));
  LUT3 #(.INIT(8'h96)) lut_n845 (.I0(n818), .I1(n826), .I2(n827), .O(n845));
  LUT3 #(.INIT(8'hE8)) lut_n846 (.I0(n836), .I1(n844), .I2(n845), .O(n846));
  LUT3 #(.INIT(8'h96)) lut_n847 (.I0(n787), .I1(n805), .I2(n806), .O(n847));
  LUT3 #(.INIT(8'hE8)) lut_n848 (.I0(n828), .I1(n846), .I2(n847), .O(n848));
  LUT3 #(.INIT(8'hE8)) lut_n849 (.I0(x432), .I1(x433), .I2(x434), .O(n849));
  LUT5 #(.INIT(32'hE81717E8)) lut_n850 (.I0(x423), .I1(x424), .I2(x425), .I3(n840), .I4(n841), .O(n850));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n851 (.I0(x429), .I1(x430), .I2(x431), .I3(n849), .I4(n850), .O(n851));
  LUT3 #(.INIT(8'hE8)) lut_n852 (.I0(x438), .I1(x439), .I2(x440), .O(n852));
  LUT5 #(.INIT(32'hE81717E8)) lut_n853 (.I0(x429), .I1(x430), .I2(x431), .I3(n849), .I4(n850), .O(n853));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n854 (.I0(x435), .I1(x436), .I2(x437), .I3(n852), .I4(n853), .O(n854));
  LUT3 #(.INIT(8'h96)) lut_n855 (.I0(n839), .I1(n842), .I2(n843), .O(n855));
  LUT3 #(.INIT(8'hE8)) lut_n856 (.I0(n851), .I1(n854), .I2(n855), .O(n856));
  LUT3 #(.INIT(8'hE8)) lut_n857 (.I0(x444), .I1(x445), .I2(x446), .O(n857));
  LUT5 #(.INIT(32'hE81717E8)) lut_n858 (.I0(x435), .I1(x436), .I2(x437), .I3(n852), .I4(n853), .O(n858));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n859 (.I0(x441), .I1(x442), .I2(x443), .I3(n857), .I4(n858), .O(n859));
  LUT3 #(.INIT(8'hE8)) lut_n860 (.I0(x450), .I1(x451), .I2(x452), .O(n860));
  LUT5 #(.INIT(32'hE81717E8)) lut_n861 (.I0(x441), .I1(x442), .I2(x443), .I3(n857), .I4(n858), .O(n861));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n862 (.I0(x447), .I1(x448), .I2(x449), .I3(n860), .I4(n861), .O(n862));
  LUT3 #(.INIT(8'h96)) lut_n863 (.I0(n851), .I1(n854), .I2(n855), .O(n863));
  LUT3 #(.INIT(8'hE8)) lut_n864 (.I0(n859), .I1(n862), .I2(n863), .O(n864));
  LUT3 #(.INIT(8'h96)) lut_n865 (.I0(n836), .I1(n844), .I2(n845), .O(n865));
  LUT3 #(.INIT(8'hE8)) lut_n866 (.I0(n856), .I1(n864), .I2(n865), .O(n866));
  LUT3 #(.INIT(8'hE8)) lut_n867 (.I0(x456), .I1(x457), .I2(x458), .O(n867));
  LUT5 #(.INIT(32'hE81717E8)) lut_n868 (.I0(x447), .I1(x448), .I2(x449), .I3(n860), .I4(n861), .O(n868));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n869 (.I0(x453), .I1(x454), .I2(x455), .I3(n867), .I4(n868), .O(n869));
  LUT3 #(.INIT(8'hE8)) lut_n870 (.I0(x462), .I1(x463), .I2(x464), .O(n870));
  LUT5 #(.INIT(32'hE81717E8)) lut_n871 (.I0(x453), .I1(x454), .I2(x455), .I3(n867), .I4(n868), .O(n871));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n872 (.I0(x459), .I1(x460), .I2(x461), .I3(n870), .I4(n871), .O(n872));
  LUT3 #(.INIT(8'h96)) lut_n873 (.I0(n859), .I1(n862), .I2(n863), .O(n873));
  LUT3 #(.INIT(8'hE8)) lut_n874 (.I0(n869), .I1(n872), .I2(n873), .O(n874));
  LUT3 #(.INIT(8'hE8)) lut_n875 (.I0(x468), .I1(x469), .I2(x470), .O(n875));
  LUT5 #(.INIT(32'hE81717E8)) lut_n876 (.I0(x459), .I1(x460), .I2(x461), .I3(n870), .I4(n871), .O(n876));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n877 (.I0(x465), .I1(x466), .I2(x467), .I3(n875), .I4(n876), .O(n877));
  LUT3 #(.INIT(8'hE8)) lut_n878 (.I0(x474), .I1(x475), .I2(x476), .O(n878));
  LUT5 #(.INIT(32'hE81717E8)) lut_n879 (.I0(x465), .I1(x466), .I2(x467), .I3(n875), .I4(n876), .O(n879));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n880 (.I0(x471), .I1(x472), .I2(x473), .I3(n878), .I4(n879), .O(n880));
  LUT3 #(.INIT(8'h96)) lut_n881 (.I0(n869), .I1(n872), .I2(n873), .O(n881));
  LUT3 #(.INIT(8'hE8)) lut_n882 (.I0(n877), .I1(n880), .I2(n881), .O(n882));
  LUT3 #(.INIT(8'h96)) lut_n883 (.I0(n856), .I1(n864), .I2(n865), .O(n883));
  LUT3 #(.INIT(8'hE8)) lut_n884 (.I0(n874), .I1(n882), .I2(n883), .O(n884));
  LUT3 #(.INIT(8'h96)) lut_n885 (.I0(n828), .I1(n846), .I2(n847), .O(n885));
  LUT3 #(.INIT(8'hE8)) lut_n886 (.I0(n866), .I1(n884), .I2(n885), .O(n886));
  LUT3 #(.INIT(8'h96)) lut_n887 (.I0(n769), .I1(n807), .I2(n808), .O(n887));
  LUT3 #(.INIT(8'hE8)) lut_n888 (.I0(n848), .I1(n886), .I2(n887), .O(n888));
  LUT3 #(.INIT(8'hE8)) lut_n889 (.I0(x480), .I1(x481), .I2(x482), .O(n889));
  LUT5 #(.INIT(32'hE81717E8)) lut_n890 (.I0(x471), .I1(x472), .I2(x473), .I3(n878), .I4(n879), .O(n890));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n891 (.I0(x477), .I1(x478), .I2(x479), .I3(n889), .I4(n890), .O(n891));
  LUT3 #(.INIT(8'hE8)) lut_n892 (.I0(x486), .I1(x487), .I2(x488), .O(n892));
  LUT5 #(.INIT(32'hE81717E8)) lut_n893 (.I0(x477), .I1(x478), .I2(x479), .I3(n889), .I4(n890), .O(n893));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n894 (.I0(x483), .I1(x484), .I2(x485), .I3(n892), .I4(n893), .O(n894));
  LUT3 #(.INIT(8'h96)) lut_n895 (.I0(n877), .I1(n880), .I2(n881), .O(n895));
  LUT3 #(.INIT(8'hE8)) lut_n896 (.I0(n891), .I1(n894), .I2(n895), .O(n896));
  LUT3 #(.INIT(8'hE8)) lut_n897 (.I0(x492), .I1(x493), .I2(x494), .O(n897));
  LUT5 #(.INIT(32'hE81717E8)) lut_n898 (.I0(x483), .I1(x484), .I2(x485), .I3(n892), .I4(n893), .O(n898));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n899 (.I0(x489), .I1(x490), .I2(x491), .I3(n897), .I4(n898), .O(n899));
  LUT3 #(.INIT(8'hE8)) lut_n900 (.I0(x498), .I1(x499), .I2(x500), .O(n900));
  LUT5 #(.INIT(32'hE81717E8)) lut_n901 (.I0(x489), .I1(x490), .I2(x491), .I3(n897), .I4(n898), .O(n901));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n902 (.I0(x495), .I1(x496), .I2(x497), .I3(n900), .I4(n901), .O(n902));
  LUT3 #(.INIT(8'h96)) lut_n903 (.I0(n891), .I1(n894), .I2(n895), .O(n903));
  LUT3 #(.INIT(8'hE8)) lut_n904 (.I0(n899), .I1(n902), .I2(n903), .O(n904));
  LUT3 #(.INIT(8'h96)) lut_n905 (.I0(n874), .I1(n882), .I2(n883), .O(n905));
  LUT3 #(.INIT(8'hE8)) lut_n906 (.I0(n896), .I1(n904), .I2(n905), .O(n906));
  LUT3 #(.INIT(8'hE8)) lut_n907 (.I0(x504), .I1(x505), .I2(x506), .O(n907));
  LUT5 #(.INIT(32'hE81717E8)) lut_n908 (.I0(x495), .I1(x496), .I2(x497), .I3(n900), .I4(n901), .O(n908));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n909 (.I0(x501), .I1(x502), .I2(x503), .I3(n907), .I4(n908), .O(n909));
  LUT3 #(.INIT(8'h96)) lut_n910 (.I0(x0), .I1(x1), .I2(x2), .O(n910));
  LUT3 #(.INIT(8'h96)) lut_n911 (.I0(x6), .I1(x7), .I2(x8), .O(n911));
  LUT5 #(.INIT(32'hFF969600)) lut_n912 (.I0(x3), .I1(x4), .I2(x5), .I3(n910), .I4(n911), .O(n912));
  LUT5 #(.INIT(32'hE81717E8)) lut_n913 (.I0(x501), .I1(x502), .I2(x503), .I3(n907), .I4(n908), .O(n913));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n914 (.I0(x507), .I1(x508), .I2(x509), .I3(n912), .I4(n913), .O(n914));
  LUT3 #(.INIT(8'h96)) lut_n915 (.I0(n899), .I1(n902), .I2(n903), .O(n915));
  LUT3 #(.INIT(8'hE8)) lut_n916 (.I0(n909), .I1(n914), .I2(n915), .O(n916));
  LUT3 #(.INIT(8'h96)) lut_n917 (.I0(x12), .I1(x13), .I2(x14), .O(n917));
  LUT5 #(.INIT(32'h96696996)) lut_n918 (.I0(x3), .I1(x4), .I2(x5), .I3(n910), .I4(n911), .O(n918));
  LUT5 #(.INIT(32'hFF969600)) lut_n919 (.I0(x9), .I1(x10), .I2(x11), .I3(n917), .I4(n918), .O(n919));
  LUT3 #(.INIT(8'h96)) lut_n920 (.I0(x18), .I1(x19), .I2(x20), .O(n920));
  LUT5 #(.INIT(32'h96696996)) lut_n921 (.I0(x9), .I1(x10), .I2(x11), .I3(n917), .I4(n918), .O(n921));
  LUT5 #(.INIT(32'hFF969600)) lut_n922 (.I0(x15), .I1(x16), .I2(x17), .I3(n920), .I4(n921), .O(n922));
  LUT5 #(.INIT(32'hE81717E8)) lut_n923 (.I0(x507), .I1(x508), .I2(x509), .I3(n912), .I4(n913), .O(n923));
  LUT3 #(.INIT(8'hE8)) lut_n924 (.I0(n919), .I1(n922), .I2(n923), .O(n924));
  LUT3 #(.INIT(8'h96)) lut_n925 (.I0(x24), .I1(x25), .I2(x26), .O(n925));
  LUT5 #(.INIT(32'h96696996)) lut_n926 (.I0(x15), .I1(x16), .I2(x17), .I3(n920), .I4(n921), .O(n926));
  LUT5 #(.INIT(32'hFF969600)) lut_n927 (.I0(x21), .I1(x22), .I2(x23), .I3(n925), .I4(n926), .O(n927));
  LUT3 #(.INIT(8'h96)) lut_n928 (.I0(x27), .I1(x28), .I2(x29), .O(n928));
  LUT5 #(.INIT(32'h96696996)) lut_n929 (.I0(x21), .I1(x22), .I2(x23), .I3(n925), .I4(n926), .O(n929));
  LUT5 #(.INIT(32'hFF969600)) lut_n930 (.I0(x30), .I1(x31), .I2(x32), .I3(n928), .I4(n929), .O(n930));
  LUT3 #(.INIT(8'h96)) lut_n931 (.I0(n919), .I1(n922), .I2(n923), .O(n931));
  LUT3 #(.INIT(8'hE8)) lut_n932 (.I0(n927), .I1(n930), .I2(n931), .O(n932));
  LUT3 #(.INIT(8'h96)) lut_n933 (.I0(n909), .I1(n914), .I2(n915), .O(n933));
  LUT3 #(.INIT(8'hE8)) lut_n934 (.I0(n924), .I1(n932), .I2(n933), .O(n934));
  LUT3 #(.INIT(8'h96)) lut_n935 (.I0(n896), .I1(n904), .I2(n905), .O(n935));
  LUT3 #(.INIT(8'hE8)) lut_n936 (.I0(n916), .I1(n934), .I2(n935), .O(n936));
  LUT3 #(.INIT(8'h96)) lut_n937 (.I0(n866), .I1(n884), .I2(n885), .O(n937));
  LUT3 #(.INIT(8'hE8)) lut_n938 (.I0(n906), .I1(n936), .I2(n937), .O(n938));
  LUT3 #(.INIT(8'h96)) lut_n939 (.I0(x36), .I1(x37), .I2(x38), .O(n939));
  LUT5 #(.INIT(32'h96696996)) lut_n940 (.I0(x30), .I1(x31), .I2(x32), .I3(n928), .I4(n929), .O(n940));
  LUT5 #(.INIT(32'hFF969600)) lut_n941 (.I0(x33), .I1(x34), .I2(x35), .I3(n939), .I4(n940), .O(n941));
  LUT3 #(.INIT(8'h96)) lut_n942 (.I0(x42), .I1(x43), .I2(x44), .O(n942));
  LUT5 #(.INIT(32'h96696996)) lut_n943 (.I0(x33), .I1(x34), .I2(x35), .I3(n939), .I4(n940), .O(n943));
  LUT5 #(.INIT(32'hFF969600)) lut_n944 (.I0(x39), .I1(x40), .I2(x41), .I3(n942), .I4(n943), .O(n944));
  LUT3 #(.INIT(8'h96)) lut_n945 (.I0(n927), .I1(n930), .I2(n931), .O(n945));
  LUT3 #(.INIT(8'hE8)) lut_n946 (.I0(n941), .I1(n944), .I2(n945), .O(n946));
  LUT3 #(.INIT(8'h96)) lut_n947 (.I0(x48), .I1(x49), .I2(x50), .O(n947));
  LUT5 #(.INIT(32'h96696996)) lut_n948 (.I0(x39), .I1(x40), .I2(x41), .I3(n942), .I4(n943), .O(n948));
  LUT5 #(.INIT(32'hFF969600)) lut_n949 (.I0(x45), .I1(x46), .I2(x47), .I3(n947), .I4(n948), .O(n949));
  LUT3 #(.INIT(8'h96)) lut_n950 (.I0(x54), .I1(x55), .I2(x56), .O(n950));
  LUT5 #(.INIT(32'h96696996)) lut_n951 (.I0(x45), .I1(x46), .I2(x47), .I3(n947), .I4(n948), .O(n951));
  LUT5 #(.INIT(32'hFF969600)) lut_n952 (.I0(x51), .I1(x52), .I2(x53), .I3(n950), .I4(n951), .O(n952));
  LUT3 #(.INIT(8'h96)) lut_n953 (.I0(n941), .I1(n944), .I2(n945), .O(n953));
  LUT3 #(.INIT(8'hE8)) lut_n954 (.I0(n949), .I1(n952), .I2(n953), .O(n954));
  LUT3 #(.INIT(8'h96)) lut_n955 (.I0(n924), .I1(n932), .I2(n933), .O(n955));
  LUT3 #(.INIT(8'hE8)) lut_n956 (.I0(n946), .I1(n954), .I2(n955), .O(n956));
  LUT3 #(.INIT(8'h96)) lut_n957 (.I0(x60), .I1(x61), .I2(x62), .O(n957));
  LUT5 #(.INIT(32'h96696996)) lut_n958 (.I0(x51), .I1(x52), .I2(x53), .I3(n950), .I4(n951), .O(n958));
  LUT5 #(.INIT(32'hFF969600)) lut_n959 (.I0(x57), .I1(x58), .I2(x59), .I3(n957), .I4(n958), .O(n959));
  LUT3 #(.INIT(8'h96)) lut_n960 (.I0(x66), .I1(x67), .I2(x68), .O(n960));
  LUT5 #(.INIT(32'h96696996)) lut_n961 (.I0(x57), .I1(x58), .I2(x59), .I3(n957), .I4(n958), .O(n961));
  LUT5 #(.INIT(32'hFF969600)) lut_n962 (.I0(x63), .I1(x64), .I2(x65), .I3(n960), .I4(n961), .O(n962));
  LUT3 #(.INIT(8'h96)) lut_n963 (.I0(n949), .I1(n952), .I2(n953), .O(n963));
  LUT3 #(.INIT(8'hE8)) lut_n964 (.I0(n959), .I1(n962), .I2(n963), .O(n964));
  LUT3 #(.INIT(8'h96)) lut_n965 (.I0(x72), .I1(x73), .I2(x74), .O(n965));
  LUT5 #(.INIT(32'h96696996)) lut_n966 (.I0(x63), .I1(x64), .I2(x65), .I3(n960), .I4(n961), .O(n966));
  LUT5 #(.INIT(32'hFF969600)) lut_n967 (.I0(x69), .I1(x70), .I2(x71), .I3(n965), .I4(n966), .O(n967));
  LUT3 #(.INIT(8'h96)) lut_n968 (.I0(x78), .I1(x79), .I2(x80), .O(n968));
  LUT5 #(.INIT(32'h96696996)) lut_n969 (.I0(x69), .I1(x70), .I2(x71), .I3(n965), .I4(n966), .O(n969));
  LUT5 #(.INIT(32'hFF969600)) lut_n970 (.I0(x75), .I1(x76), .I2(x77), .I3(n968), .I4(n969), .O(n970));
  LUT3 #(.INIT(8'h96)) lut_n971 (.I0(n959), .I1(n962), .I2(n963), .O(n971));
  LUT3 #(.INIT(8'hE8)) lut_n972 (.I0(n967), .I1(n970), .I2(n971), .O(n972));
  LUT3 #(.INIT(8'h96)) lut_n973 (.I0(n946), .I1(n954), .I2(n955), .O(n973));
  LUT3 #(.INIT(8'hE8)) lut_n974 (.I0(n964), .I1(n972), .I2(n973), .O(n974));
  LUT3 #(.INIT(8'h96)) lut_n975 (.I0(n916), .I1(n934), .I2(n935), .O(n975));
  LUT3 #(.INIT(8'hE8)) lut_n976 (.I0(n956), .I1(n974), .I2(n975), .O(n976));
  LUT3 #(.INIT(8'h96)) lut_n977 (.I0(x84), .I1(x85), .I2(x86), .O(n977));
  LUT5 #(.INIT(32'h96696996)) lut_n978 (.I0(x75), .I1(x76), .I2(x77), .I3(n968), .I4(n969), .O(n978));
  LUT5 #(.INIT(32'hFF969600)) lut_n979 (.I0(x81), .I1(x82), .I2(x83), .I3(n977), .I4(n978), .O(n979));
  LUT3 #(.INIT(8'h96)) lut_n980 (.I0(x90), .I1(x91), .I2(x92), .O(n980));
  LUT5 #(.INIT(32'h96696996)) lut_n981 (.I0(x81), .I1(x82), .I2(x83), .I3(n977), .I4(n978), .O(n981));
  LUT5 #(.INIT(32'hFF969600)) lut_n982 (.I0(x87), .I1(x88), .I2(x89), .I3(n980), .I4(n981), .O(n982));
  LUT3 #(.INIT(8'h96)) lut_n983 (.I0(n967), .I1(n970), .I2(n971), .O(n983));
  LUT3 #(.INIT(8'hE8)) lut_n984 (.I0(n979), .I1(n982), .I2(n983), .O(n984));
  LUT3 #(.INIT(8'h96)) lut_n985 (.I0(x96), .I1(x97), .I2(x98), .O(n985));
  LUT5 #(.INIT(32'h96696996)) lut_n986 (.I0(x87), .I1(x88), .I2(x89), .I3(n980), .I4(n981), .O(n986));
  LUT5 #(.INIT(32'hFF969600)) lut_n987 (.I0(x93), .I1(x94), .I2(x95), .I3(n985), .I4(n986), .O(n987));
  LUT3 #(.INIT(8'h96)) lut_n988 (.I0(x102), .I1(x103), .I2(x104), .O(n988));
  LUT5 #(.INIT(32'h96696996)) lut_n989 (.I0(x93), .I1(x94), .I2(x95), .I3(n985), .I4(n986), .O(n989));
  LUT5 #(.INIT(32'hFF969600)) lut_n990 (.I0(x99), .I1(x100), .I2(x101), .I3(n988), .I4(n989), .O(n990));
  LUT3 #(.INIT(8'h96)) lut_n991 (.I0(n979), .I1(n982), .I2(n983), .O(n991));
  LUT3 #(.INIT(8'hE8)) lut_n992 (.I0(n987), .I1(n990), .I2(n991), .O(n992));
  LUT3 #(.INIT(8'h96)) lut_n993 (.I0(n964), .I1(n972), .I2(n973), .O(n993));
  LUT3 #(.INIT(8'hE8)) lut_n994 (.I0(n984), .I1(n992), .I2(n993), .O(n994));
  LUT3 #(.INIT(8'h96)) lut_n995 (.I0(x108), .I1(x109), .I2(x110), .O(n995));
  LUT5 #(.INIT(32'h96696996)) lut_n996 (.I0(x99), .I1(x100), .I2(x101), .I3(n988), .I4(n989), .O(n996));
  LUT5 #(.INIT(32'hFF969600)) lut_n997 (.I0(x105), .I1(x106), .I2(x107), .I3(n995), .I4(n996), .O(n997));
  LUT3 #(.INIT(8'h96)) lut_n998 (.I0(x114), .I1(x115), .I2(x116), .O(n998));
  LUT5 #(.INIT(32'h96696996)) lut_n999 (.I0(x105), .I1(x106), .I2(x107), .I3(n995), .I4(n996), .O(n999));
  LUT5 #(.INIT(32'hFF969600)) lut_n1000 (.I0(x111), .I1(x112), .I2(x113), .I3(n998), .I4(n999), .O(n1000));
  LUT3 #(.INIT(8'h96)) lut_n1001 (.I0(n987), .I1(n990), .I2(n991), .O(n1001));
  LUT3 #(.INIT(8'hE8)) lut_n1002 (.I0(n997), .I1(n1000), .I2(n1001), .O(n1002));
  LUT3 #(.INIT(8'h96)) lut_n1003 (.I0(x120), .I1(x121), .I2(x122), .O(n1003));
  LUT5 #(.INIT(32'h96696996)) lut_n1004 (.I0(x111), .I1(x112), .I2(x113), .I3(n998), .I4(n999), .O(n1004));
  LUT5 #(.INIT(32'hFF969600)) lut_n1005 (.I0(x117), .I1(x118), .I2(x119), .I3(n1003), .I4(n1004), .O(n1005));
  LUT3 #(.INIT(8'h96)) lut_n1006 (.I0(x126), .I1(x127), .I2(x128), .O(n1006));
  LUT5 #(.INIT(32'h96696996)) lut_n1007 (.I0(x117), .I1(x118), .I2(x119), .I3(n1003), .I4(n1004), .O(n1007));
  LUT5 #(.INIT(32'hFF969600)) lut_n1008 (.I0(x123), .I1(x124), .I2(x125), .I3(n1006), .I4(n1007), .O(n1008));
  LUT3 #(.INIT(8'h96)) lut_n1009 (.I0(n997), .I1(n1000), .I2(n1001), .O(n1009));
  LUT3 #(.INIT(8'hE8)) lut_n1010 (.I0(n1005), .I1(n1008), .I2(n1009), .O(n1010));
  LUT3 #(.INIT(8'h96)) lut_n1011 (.I0(n984), .I1(n992), .I2(n993), .O(n1011));
  LUT3 #(.INIT(8'hE8)) lut_n1012 (.I0(n1002), .I1(n1010), .I2(n1011), .O(n1012));
  LUT3 #(.INIT(8'h96)) lut_n1013 (.I0(n956), .I1(n974), .I2(n975), .O(n1013));
  LUT3 #(.INIT(8'hE8)) lut_n1014 (.I0(n994), .I1(n1012), .I2(n1013), .O(n1014));
  LUT3 #(.INIT(8'h96)) lut_n1015 (.I0(n906), .I1(n936), .I2(n937), .O(n1015));
  LUT3 #(.INIT(8'hE8)) lut_n1016 (.I0(n976), .I1(n1014), .I2(n1015), .O(n1016));
  LUT3 #(.INIT(8'h96)) lut_n1017 (.I0(n848), .I1(n886), .I2(n887), .O(n1017));
  LUT3 #(.INIT(8'hE8)) lut_n1018 (.I0(n938), .I1(n1016), .I2(n1017), .O(n1018));
  LUT3 #(.INIT(8'h96)) lut_n1019 (.I0(n653), .I1(n731), .I2(n809), .O(n1019));
  LUT3 #(.INIT(8'h96)) lut_n1020 (.I0(x132), .I1(x133), .I2(x134), .O(n1020));
  LUT5 #(.INIT(32'h96696996)) lut_n1021 (.I0(x123), .I1(x124), .I2(x125), .I3(n1006), .I4(n1007), .O(n1021));
  LUT5 #(.INIT(32'hFF969600)) lut_n1022 (.I0(x129), .I1(x130), .I2(x131), .I3(n1020), .I4(n1021), .O(n1022));
  LUT3 #(.INIT(8'h96)) lut_n1023 (.I0(x138), .I1(x139), .I2(x140), .O(n1023));
  LUT5 #(.INIT(32'h96696996)) lut_n1024 (.I0(x129), .I1(x130), .I2(x131), .I3(n1020), .I4(n1021), .O(n1024));
  LUT5 #(.INIT(32'hFF969600)) lut_n1025 (.I0(x135), .I1(x136), .I2(x137), .I3(n1023), .I4(n1024), .O(n1025));
  LUT3 #(.INIT(8'h96)) lut_n1026 (.I0(n1005), .I1(n1008), .I2(n1009), .O(n1026));
  LUT3 #(.INIT(8'hE8)) lut_n1027 (.I0(n1022), .I1(n1025), .I2(n1026), .O(n1027));
  LUT3 #(.INIT(8'h96)) lut_n1028 (.I0(x144), .I1(x145), .I2(x146), .O(n1028));
  LUT5 #(.INIT(32'h96696996)) lut_n1029 (.I0(x135), .I1(x136), .I2(x137), .I3(n1023), .I4(n1024), .O(n1029));
  LUT5 #(.INIT(32'hFF969600)) lut_n1030 (.I0(x141), .I1(x142), .I2(x143), .I3(n1028), .I4(n1029), .O(n1030));
  LUT3 #(.INIT(8'h96)) lut_n1031 (.I0(x150), .I1(x151), .I2(x152), .O(n1031));
  LUT5 #(.INIT(32'h96696996)) lut_n1032 (.I0(x141), .I1(x142), .I2(x143), .I3(n1028), .I4(n1029), .O(n1032));
  LUT5 #(.INIT(32'hFF969600)) lut_n1033 (.I0(x147), .I1(x148), .I2(x149), .I3(n1031), .I4(n1032), .O(n1033));
  LUT3 #(.INIT(8'h96)) lut_n1034 (.I0(n1022), .I1(n1025), .I2(n1026), .O(n1034));
  LUT3 #(.INIT(8'hE8)) lut_n1035 (.I0(n1030), .I1(n1033), .I2(n1034), .O(n1035));
  LUT3 #(.INIT(8'h96)) lut_n1036 (.I0(n1002), .I1(n1010), .I2(n1011), .O(n1036));
  LUT3 #(.INIT(8'hE8)) lut_n1037 (.I0(n1027), .I1(n1035), .I2(n1036), .O(n1037));
  LUT3 #(.INIT(8'h96)) lut_n1038 (.I0(x156), .I1(x157), .I2(x158), .O(n1038));
  LUT5 #(.INIT(32'h96696996)) lut_n1039 (.I0(x147), .I1(x148), .I2(x149), .I3(n1031), .I4(n1032), .O(n1039));
  LUT5 #(.INIT(32'hFF969600)) lut_n1040 (.I0(x153), .I1(x154), .I2(x155), .I3(n1038), .I4(n1039), .O(n1040));
  LUT3 #(.INIT(8'h96)) lut_n1041 (.I0(x162), .I1(x163), .I2(x164), .O(n1041));
  LUT5 #(.INIT(32'h96696996)) lut_n1042 (.I0(x153), .I1(x154), .I2(x155), .I3(n1038), .I4(n1039), .O(n1042));
  LUT5 #(.INIT(32'hFF969600)) lut_n1043 (.I0(x159), .I1(x160), .I2(x161), .I3(n1041), .I4(n1042), .O(n1043));
  LUT3 #(.INIT(8'h96)) lut_n1044 (.I0(n1030), .I1(n1033), .I2(n1034), .O(n1044));
  LUT3 #(.INIT(8'hE8)) lut_n1045 (.I0(n1040), .I1(n1043), .I2(n1044), .O(n1045));
  LUT3 #(.INIT(8'h96)) lut_n1046 (.I0(x168), .I1(x169), .I2(x170), .O(n1046));
  LUT5 #(.INIT(32'h96696996)) lut_n1047 (.I0(x159), .I1(x160), .I2(x161), .I3(n1041), .I4(n1042), .O(n1047));
  LUT5 #(.INIT(32'hFF969600)) lut_n1048 (.I0(x165), .I1(x166), .I2(x167), .I3(n1046), .I4(n1047), .O(n1048));
  LUT3 #(.INIT(8'h96)) lut_n1049 (.I0(x174), .I1(x175), .I2(x176), .O(n1049));
  LUT5 #(.INIT(32'h96696996)) lut_n1050 (.I0(x165), .I1(x166), .I2(x167), .I3(n1046), .I4(n1047), .O(n1050));
  LUT5 #(.INIT(32'hFF969600)) lut_n1051 (.I0(x171), .I1(x172), .I2(x173), .I3(n1049), .I4(n1050), .O(n1051));
  LUT3 #(.INIT(8'h96)) lut_n1052 (.I0(n1040), .I1(n1043), .I2(n1044), .O(n1052));
  LUT3 #(.INIT(8'hE8)) lut_n1053 (.I0(n1048), .I1(n1051), .I2(n1052), .O(n1053));
  LUT3 #(.INIT(8'h96)) lut_n1054 (.I0(n1027), .I1(n1035), .I2(n1036), .O(n1054));
  LUT3 #(.INIT(8'hE8)) lut_n1055 (.I0(n1045), .I1(n1053), .I2(n1054), .O(n1055));
  LUT3 #(.INIT(8'h96)) lut_n1056 (.I0(n994), .I1(n1012), .I2(n1013), .O(n1056));
  LUT3 #(.INIT(8'hE8)) lut_n1057 (.I0(n1037), .I1(n1055), .I2(n1056), .O(n1057));
  LUT3 #(.INIT(8'h96)) lut_n1058 (.I0(x180), .I1(x181), .I2(x182), .O(n1058));
  LUT5 #(.INIT(32'h96696996)) lut_n1059 (.I0(x171), .I1(x172), .I2(x173), .I3(n1049), .I4(n1050), .O(n1059));
  LUT5 #(.INIT(32'hFF969600)) lut_n1060 (.I0(x177), .I1(x178), .I2(x179), .I3(n1058), .I4(n1059), .O(n1060));
  LUT3 #(.INIT(8'h96)) lut_n1061 (.I0(x186), .I1(x187), .I2(x188), .O(n1061));
  LUT5 #(.INIT(32'h96696996)) lut_n1062 (.I0(x177), .I1(x178), .I2(x179), .I3(n1058), .I4(n1059), .O(n1062));
  LUT5 #(.INIT(32'hFF969600)) lut_n1063 (.I0(x183), .I1(x184), .I2(x185), .I3(n1061), .I4(n1062), .O(n1063));
  LUT3 #(.INIT(8'h96)) lut_n1064 (.I0(n1048), .I1(n1051), .I2(n1052), .O(n1064));
  LUT3 #(.INIT(8'hE8)) lut_n1065 (.I0(n1060), .I1(n1063), .I2(n1064), .O(n1065));
  LUT3 #(.INIT(8'h96)) lut_n1066 (.I0(x192), .I1(x193), .I2(x194), .O(n1066));
  LUT5 #(.INIT(32'h96696996)) lut_n1067 (.I0(x183), .I1(x184), .I2(x185), .I3(n1061), .I4(n1062), .O(n1067));
  LUT5 #(.INIT(32'hFF969600)) lut_n1068 (.I0(x189), .I1(x190), .I2(x191), .I3(n1066), .I4(n1067), .O(n1068));
  LUT3 #(.INIT(8'h96)) lut_n1069 (.I0(x198), .I1(x199), .I2(x200), .O(n1069));
  LUT5 #(.INIT(32'h96696996)) lut_n1070 (.I0(x189), .I1(x190), .I2(x191), .I3(n1066), .I4(n1067), .O(n1070));
  LUT5 #(.INIT(32'hFF969600)) lut_n1071 (.I0(x195), .I1(x196), .I2(x197), .I3(n1069), .I4(n1070), .O(n1071));
  LUT3 #(.INIT(8'h96)) lut_n1072 (.I0(n1060), .I1(n1063), .I2(n1064), .O(n1072));
  LUT3 #(.INIT(8'hE8)) lut_n1073 (.I0(n1068), .I1(n1071), .I2(n1072), .O(n1073));
  LUT3 #(.INIT(8'h96)) lut_n1074 (.I0(n1045), .I1(n1053), .I2(n1054), .O(n1074));
  LUT3 #(.INIT(8'hE8)) lut_n1075 (.I0(n1065), .I1(n1073), .I2(n1074), .O(n1075));
  LUT3 #(.INIT(8'h96)) lut_n1076 (.I0(x204), .I1(x205), .I2(x206), .O(n1076));
  LUT5 #(.INIT(32'h96696996)) lut_n1077 (.I0(x195), .I1(x196), .I2(x197), .I3(n1069), .I4(n1070), .O(n1077));
  LUT5 #(.INIT(32'hFF969600)) lut_n1078 (.I0(x201), .I1(x202), .I2(x203), .I3(n1076), .I4(n1077), .O(n1078));
  LUT3 #(.INIT(8'h96)) lut_n1079 (.I0(x210), .I1(x211), .I2(x212), .O(n1079));
  LUT5 #(.INIT(32'h96696996)) lut_n1080 (.I0(x201), .I1(x202), .I2(x203), .I3(n1076), .I4(n1077), .O(n1080));
  LUT5 #(.INIT(32'hFF969600)) lut_n1081 (.I0(x207), .I1(x208), .I2(x209), .I3(n1079), .I4(n1080), .O(n1081));
  LUT3 #(.INIT(8'h96)) lut_n1082 (.I0(n1068), .I1(n1071), .I2(n1072), .O(n1082));
  LUT3 #(.INIT(8'hE8)) lut_n1083 (.I0(n1078), .I1(n1081), .I2(n1082), .O(n1083));
  LUT3 #(.INIT(8'h96)) lut_n1084 (.I0(x216), .I1(x217), .I2(x218), .O(n1084));
  LUT5 #(.INIT(32'h96696996)) lut_n1085 (.I0(x207), .I1(x208), .I2(x209), .I3(n1079), .I4(n1080), .O(n1085));
  LUT5 #(.INIT(32'hFF969600)) lut_n1086 (.I0(x213), .I1(x214), .I2(x215), .I3(n1084), .I4(n1085), .O(n1086));
  LUT3 #(.INIT(8'h96)) lut_n1087 (.I0(x222), .I1(x223), .I2(x224), .O(n1087));
  LUT5 #(.INIT(32'h96696996)) lut_n1088 (.I0(x213), .I1(x214), .I2(x215), .I3(n1084), .I4(n1085), .O(n1088));
  LUT5 #(.INIT(32'hFF969600)) lut_n1089 (.I0(x219), .I1(x220), .I2(x221), .I3(n1087), .I4(n1088), .O(n1089));
  LUT3 #(.INIT(8'h96)) lut_n1090 (.I0(n1078), .I1(n1081), .I2(n1082), .O(n1090));
  LUT3 #(.INIT(8'hE8)) lut_n1091 (.I0(n1086), .I1(n1089), .I2(n1090), .O(n1091));
  LUT3 #(.INIT(8'h96)) lut_n1092 (.I0(n1065), .I1(n1073), .I2(n1074), .O(n1092));
  LUT3 #(.INIT(8'hE8)) lut_n1093 (.I0(n1083), .I1(n1091), .I2(n1092), .O(n1093));
  LUT3 #(.INIT(8'h96)) lut_n1094 (.I0(n1037), .I1(n1055), .I2(n1056), .O(n1094));
  LUT3 #(.INIT(8'hE8)) lut_n1095 (.I0(n1075), .I1(n1093), .I2(n1094), .O(n1095));
  LUT3 #(.INIT(8'h96)) lut_n1096 (.I0(n976), .I1(n1014), .I2(n1015), .O(n1096));
  LUT3 #(.INIT(8'hE8)) lut_n1097 (.I0(n1057), .I1(n1095), .I2(n1096), .O(n1097));
  LUT3 #(.INIT(8'h96)) lut_n1098 (.I0(x228), .I1(x229), .I2(x230), .O(n1098));
  LUT5 #(.INIT(32'h96696996)) lut_n1099 (.I0(x219), .I1(x220), .I2(x221), .I3(n1087), .I4(n1088), .O(n1099));
  LUT5 #(.INIT(32'hFF969600)) lut_n1100 (.I0(x225), .I1(x226), .I2(x227), .I3(n1098), .I4(n1099), .O(n1100));
  LUT3 #(.INIT(8'h96)) lut_n1101 (.I0(x234), .I1(x235), .I2(x236), .O(n1101));
  LUT5 #(.INIT(32'h96696996)) lut_n1102 (.I0(x225), .I1(x226), .I2(x227), .I3(n1098), .I4(n1099), .O(n1102));
  LUT5 #(.INIT(32'hFF969600)) lut_n1103 (.I0(x231), .I1(x232), .I2(x233), .I3(n1101), .I4(n1102), .O(n1103));
  LUT3 #(.INIT(8'h96)) lut_n1104 (.I0(n1086), .I1(n1089), .I2(n1090), .O(n1104));
  LUT3 #(.INIT(8'hE8)) lut_n1105 (.I0(n1100), .I1(n1103), .I2(n1104), .O(n1105));
  LUT3 #(.INIT(8'h96)) lut_n1106 (.I0(x240), .I1(x241), .I2(x242), .O(n1106));
  LUT5 #(.INIT(32'h96696996)) lut_n1107 (.I0(x231), .I1(x232), .I2(x233), .I3(n1101), .I4(n1102), .O(n1107));
  LUT5 #(.INIT(32'hFF969600)) lut_n1108 (.I0(x237), .I1(x238), .I2(x239), .I3(n1106), .I4(n1107), .O(n1108));
  LUT3 #(.INIT(8'h96)) lut_n1109 (.I0(x246), .I1(x247), .I2(x248), .O(n1109));
  LUT5 #(.INIT(32'h96696996)) lut_n1110 (.I0(x237), .I1(x238), .I2(x239), .I3(n1106), .I4(n1107), .O(n1110));
  LUT5 #(.INIT(32'hFF969600)) lut_n1111 (.I0(x243), .I1(x244), .I2(x245), .I3(n1109), .I4(n1110), .O(n1111));
  LUT3 #(.INIT(8'h96)) lut_n1112 (.I0(n1100), .I1(n1103), .I2(n1104), .O(n1112));
  LUT3 #(.INIT(8'hE8)) lut_n1113 (.I0(n1108), .I1(n1111), .I2(n1112), .O(n1113));
  LUT3 #(.INIT(8'h96)) lut_n1114 (.I0(n1083), .I1(n1091), .I2(n1092), .O(n1114));
  LUT3 #(.INIT(8'hE8)) lut_n1115 (.I0(n1105), .I1(n1113), .I2(n1114), .O(n1115));
  LUT3 #(.INIT(8'h96)) lut_n1116 (.I0(x252), .I1(x253), .I2(x254), .O(n1116));
  LUT5 #(.INIT(32'h96696996)) lut_n1117 (.I0(x243), .I1(x244), .I2(x245), .I3(n1109), .I4(n1110), .O(n1117));
  LUT5 #(.INIT(32'hFF969600)) lut_n1118 (.I0(x249), .I1(x250), .I2(x251), .I3(n1116), .I4(n1117), .O(n1118));
  LUT3 #(.INIT(8'h96)) lut_n1119 (.I0(x258), .I1(x259), .I2(x260), .O(n1119));
  LUT5 #(.INIT(32'h96696996)) lut_n1120 (.I0(x249), .I1(x250), .I2(x251), .I3(n1116), .I4(n1117), .O(n1120));
  LUT5 #(.INIT(32'hFF969600)) lut_n1121 (.I0(x255), .I1(x256), .I2(x257), .I3(n1119), .I4(n1120), .O(n1121));
  LUT3 #(.INIT(8'h96)) lut_n1122 (.I0(n1108), .I1(n1111), .I2(n1112), .O(n1122));
  LUT3 #(.INIT(8'hE8)) lut_n1123 (.I0(n1118), .I1(n1121), .I2(n1122), .O(n1123));
  LUT3 #(.INIT(8'h96)) lut_n1124 (.I0(x264), .I1(x265), .I2(x266), .O(n1124));
  LUT5 #(.INIT(32'h96696996)) lut_n1125 (.I0(x255), .I1(x256), .I2(x257), .I3(n1119), .I4(n1120), .O(n1125));
  LUT5 #(.INIT(32'hFF969600)) lut_n1126 (.I0(x261), .I1(x262), .I2(x263), .I3(n1124), .I4(n1125), .O(n1126));
  LUT3 #(.INIT(8'h96)) lut_n1127 (.I0(x270), .I1(x271), .I2(x272), .O(n1127));
  LUT5 #(.INIT(32'h96696996)) lut_n1128 (.I0(x261), .I1(x262), .I2(x263), .I3(n1124), .I4(n1125), .O(n1128));
  LUT5 #(.INIT(32'hFF969600)) lut_n1129 (.I0(x267), .I1(x268), .I2(x269), .I3(n1127), .I4(n1128), .O(n1129));
  LUT3 #(.INIT(8'h96)) lut_n1130 (.I0(n1118), .I1(n1121), .I2(n1122), .O(n1130));
  LUT3 #(.INIT(8'hE8)) lut_n1131 (.I0(n1126), .I1(n1129), .I2(n1130), .O(n1131));
  LUT3 #(.INIT(8'h96)) lut_n1132 (.I0(n1105), .I1(n1113), .I2(n1114), .O(n1132));
  LUT3 #(.INIT(8'hE8)) lut_n1133 (.I0(n1123), .I1(n1131), .I2(n1132), .O(n1133));
  LUT3 #(.INIT(8'h96)) lut_n1134 (.I0(n1075), .I1(n1093), .I2(n1094), .O(n1134));
  LUT3 #(.INIT(8'hE8)) lut_n1135 (.I0(n1115), .I1(n1133), .I2(n1134), .O(n1135));
  LUT3 #(.INIT(8'h96)) lut_n1136 (.I0(x276), .I1(x277), .I2(x278), .O(n1136));
  LUT5 #(.INIT(32'h96696996)) lut_n1137 (.I0(x267), .I1(x268), .I2(x269), .I3(n1127), .I4(n1128), .O(n1137));
  LUT5 #(.INIT(32'hFF969600)) lut_n1138 (.I0(x273), .I1(x274), .I2(x275), .I3(n1136), .I4(n1137), .O(n1138));
  LUT3 #(.INIT(8'h96)) lut_n1139 (.I0(x282), .I1(x283), .I2(x284), .O(n1139));
  LUT5 #(.INIT(32'h96696996)) lut_n1140 (.I0(x273), .I1(x274), .I2(x275), .I3(n1136), .I4(n1137), .O(n1140));
  LUT5 #(.INIT(32'hFF969600)) lut_n1141 (.I0(x279), .I1(x280), .I2(x281), .I3(n1139), .I4(n1140), .O(n1141));
  LUT3 #(.INIT(8'h96)) lut_n1142 (.I0(n1126), .I1(n1129), .I2(n1130), .O(n1142));
  LUT3 #(.INIT(8'hE8)) lut_n1143 (.I0(n1138), .I1(n1141), .I2(n1142), .O(n1143));
  LUT3 #(.INIT(8'h96)) lut_n1144 (.I0(x288), .I1(x289), .I2(x290), .O(n1144));
  LUT5 #(.INIT(32'h96696996)) lut_n1145 (.I0(x279), .I1(x280), .I2(x281), .I3(n1139), .I4(n1140), .O(n1145));
  LUT5 #(.INIT(32'hFF969600)) lut_n1146 (.I0(x285), .I1(x286), .I2(x287), .I3(n1144), .I4(n1145), .O(n1146));
  LUT3 #(.INIT(8'h96)) lut_n1147 (.I0(x294), .I1(x295), .I2(x296), .O(n1147));
  LUT5 #(.INIT(32'h96696996)) lut_n1148 (.I0(x285), .I1(x286), .I2(x287), .I3(n1144), .I4(n1145), .O(n1148));
  LUT5 #(.INIT(32'hFF969600)) lut_n1149 (.I0(x291), .I1(x292), .I2(x293), .I3(n1147), .I4(n1148), .O(n1149));
  LUT3 #(.INIT(8'h96)) lut_n1150 (.I0(n1138), .I1(n1141), .I2(n1142), .O(n1150));
  LUT3 #(.INIT(8'hE8)) lut_n1151 (.I0(n1146), .I1(n1149), .I2(n1150), .O(n1151));
  LUT3 #(.INIT(8'h96)) lut_n1152 (.I0(n1123), .I1(n1131), .I2(n1132), .O(n1152));
  LUT3 #(.INIT(8'hE8)) lut_n1153 (.I0(n1143), .I1(n1151), .I2(n1152), .O(n1153));
  LUT3 #(.INIT(8'h96)) lut_n1154 (.I0(x297), .I1(x298), .I2(x299), .O(n1154));
  LUT5 #(.INIT(32'h96696996)) lut_n1155 (.I0(x291), .I1(x292), .I2(x293), .I3(n1147), .I4(n1148), .O(n1155));
  LUT5 #(.INIT(32'hFF969600)) lut_n1156 (.I0(x300), .I1(x301), .I2(x302), .I3(n1154), .I4(n1155), .O(n1156));
  LUT3 #(.INIT(8'h96)) lut_n1157 (.I0(x306), .I1(x307), .I2(x308), .O(n1157));
  LUT5 #(.INIT(32'h96696996)) lut_n1158 (.I0(x300), .I1(x301), .I2(x302), .I3(n1154), .I4(n1155), .O(n1158));
  LUT5 #(.INIT(32'hFF969600)) lut_n1159 (.I0(x303), .I1(x304), .I2(x305), .I3(n1157), .I4(n1158), .O(n1159));
  LUT3 #(.INIT(8'h96)) lut_n1160 (.I0(n1146), .I1(n1149), .I2(n1150), .O(n1160));
  LUT3 #(.INIT(8'hE8)) lut_n1161 (.I0(n1156), .I1(n1159), .I2(n1160), .O(n1161));
  LUT3 #(.INIT(8'h96)) lut_n1162 (.I0(x312), .I1(x313), .I2(x314), .O(n1162));
  LUT5 #(.INIT(32'h96696996)) lut_n1163 (.I0(x303), .I1(x304), .I2(x305), .I3(n1157), .I4(n1158), .O(n1163));
  LUT5 #(.INIT(32'hFF969600)) lut_n1164 (.I0(x309), .I1(x310), .I2(x311), .I3(n1162), .I4(n1163), .O(n1164));
  LUT3 #(.INIT(8'h96)) lut_n1165 (.I0(x318), .I1(x319), .I2(x320), .O(n1165));
  LUT5 #(.INIT(32'h96696996)) lut_n1166 (.I0(x309), .I1(x310), .I2(x311), .I3(n1162), .I4(n1163), .O(n1166));
  LUT5 #(.INIT(32'hFF969600)) lut_n1167 (.I0(x315), .I1(x316), .I2(x317), .I3(n1165), .I4(n1166), .O(n1167));
  LUT3 #(.INIT(8'h96)) lut_n1168 (.I0(n1156), .I1(n1159), .I2(n1160), .O(n1168));
  LUT3 #(.INIT(8'hE8)) lut_n1169 (.I0(n1164), .I1(n1167), .I2(n1168), .O(n1169));
  LUT3 #(.INIT(8'h96)) lut_n1170 (.I0(n1143), .I1(n1151), .I2(n1152), .O(n1170));
  LUT3 #(.INIT(8'hE8)) lut_n1171 (.I0(n1161), .I1(n1169), .I2(n1170), .O(n1171));
  LUT3 #(.INIT(8'h96)) lut_n1172 (.I0(n1115), .I1(n1133), .I2(n1134), .O(n1172));
  LUT3 #(.INIT(8'hE8)) lut_n1173 (.I0(n1153), .I1(n1171), .I2(n1172), .O(n1173));
  LUT3 #(.INIT(8'h96)) lut_n1174 (.I0(n1057), .I1(n1095), .I2(n1096), .O(n1174));
  LUT3 #(.INIT(8'hE8)) lut_n1175 (.I0(n1135), .I1(n1173), .I2(n1174), .O(n1175));
  LUT3 #(.INIT(8'h96)) lut_n1176 (.I0(n938), .I1(n1016), .I2(n1017), .O(n1176));
  LUT3 #(.INIT(8'hE8)) lut_n1177 (.I0(n1097), .I1(n1175), .I2(n1176), .O(n1177));
  LUT3 #(.INIT(8'h96)) lut_n1178 (.I0(x324), .I1(x325), .I2(x326), .O(n1178));
  LUT5 #(.INIT(32'h96696996)) lut_n1179 (.I0(x315), .I1(x316), .I2(x317), .I3(n1165), .I4(n1166), .O(n1179));
  LUT5 #(.INIT(32'hFF969600)) lut_n1180 (.I0(x321), .I1(x322), .I2(x323), .I3(n1178), .I4(n1179), .O(n1180));
  LUT3 #(.INIT(8'h96)) lut_n1181 (.I0(x330), .I1(x331), .I2(x332), .O(n1181));
  LUT5 #(.INIT(32'h96696996)) lut_n1182 (.I0(x321), .I1(x322), .I2(x323), .I3(n1178), .I4(n1179), .O(n1182));
  LUT5 #(.INIT(32'hFF969600)) lut_n1183 (.I0(x327), .I1(x328), .I2(x329), .I3(n1181), .I4(n1182), .O(n1183));
  LUT3 #(.INIT(8'h96)) lut_n1184 (.I0(n1164), .I1(n1167), .I2(n1168), .O(n1184));
  LUT3 #(.INIT(8'hE8)) lut_n1185 (.I0(n1180), .I1(n1183), .I2(n1184), .O(n1185));
  LUT3 #(.INIT(8'h96)) lut_n1186 (.I0(x336), .I1(x337), .I2(x338), .O(n1186));
  LUT5 #(.INIT(32'h96696996)) lut_n1187 (.I0(x327), .I1(x328), .I2(x329), .I3(n1181), .I4(n1182), .O(n1187));
  LUT5 #(.INIT(32'hFF969600)) lut_n1188 (.I0(x333), .I1(x334), .I2(x335), .I3(n1186), .I4(n1187), .O(n1188));
  LUT3 #(.INIT(8'h96)) lut_n1189 (.I0(x342), .I1(x343), .I2(x344), .O(n1189));
  LUT5 #(.INIT(32'h96696996)) lut_n1190 (.I0(x333), .I1(x334), .I2(x335), .I3(n1186), .I4(n1187), .O(n1190));
  LUT5 #(.INIT(32'hFF969600)) lut_n1191 (.I0(x339), .I1(x340), .I2(x341), .I3(n1189), .I4(n1190), .O(n1191));
  LUT3 #(.INIT(8'h96)) lut_n1192 (.I0(n1180), .I1(n1183), .I2(n1184), .O(n1192));
  LUT3 #(.INIT(8'hE8)) lut_n1193 (.I0(n1188), .I1(n1191), .I2(n1192), .O(n1193));
  LUT3 #(.INIT(8'h96)) lut_n1194 (.I0(n1161), .I1(n1169), .I2(n1170), .O(n1194));
  LUT3 #(.INIT(8'hE8)) lut_n1195 (.I0(n1185), .I1(n1193), .I2(n1194), .O(n1195));
  LUT3 #(.INIT(8'h96)) lut_n1196 (.I0(x348), .I1(x349), .I2(x350), .O(n1196));
  LUT5 #(.INIT(32'h96696996)) lut_n1197 (.I0(x339), .I1(x340), .I2(x341), .I3(n1189), .I4(n1190), .O(n1197));
  LUT5 #(.INIT(32'hFF969600)) lut_n1198 (.I0(x345), .I1(x346), .I2(x347), .I3(n1196), .I4(n1197), .O(n1198));
  LUT3 #(.INIT(8'h96)) lut_n1199 (.I0(x354), .I1(x355), .I2(x356), .O(n1199));
  LUT5 #(.INIT(32'h96696996)) lut_n1200 (.I0(x345), .I1(x346), .I2(x347), .I3(n1196), .I4(n1197), .O(n1200));
  LUT5 #(.INIT(32'hFF969600)) lut_n1201 (.I0(x351), .I1(x352), .I2(x353), .I3(n1199), .I4(n1200), .O(n1201));
  LUT3 #(.INIT(8'h96)) lut_n1202 (.I0(n1188), .I1(n1191), .I2(n1192), .O(n1202));
  LUT3 #(.INIT(8'hE8)) lut_n1203 (.I0(n1198), .I1(n1201), .I2(n1202), .O(n1203));
  LUT3 #(.INIT(8'h96)) lut_n1204 (.I0(x360), .I1(x361), .I2(x362), .O(n1204));
  LUT5 #(.INIT(32'h96696996)) lut_n1205 (.I0(x351), .I1(x352), .I2(x353), .I3(n1199), .I4(n1200), .O(n1205));
  LUT5 #(.INIT(32'hFF969600)) lut_n1206 (.I0(x357), .I1(x358), .I2(x359), .I3(n1204), .I4(n1205), .O(n1206));
  LUT3 #(.INIT(8'h96)) lut_n1207 (.I0(x366), .I1(x367), .I2(x368), .O(n1207));
  LUT5 #(.INIT(32'h96696996)) lut_n1208 (.I0(x357), .I1(x358), .I2(x359), .I3(n1204), .I4(n1205), .O(n1208));
  LUT5 #(.INIT(32'hFF969600)) lut_n1209 (.I0(x363), .I1(x364), .I2(x365), .I3(n1207), .I4(n1208), .O(n1209));
  LUT3 #(.INIT(8'h96)) lut_n1210 (.I0(n1198), .I1(n1201), .I2(n1202), .O(n1210));
  LUT3 #(.INIT(8'hE8)) lut_n1211 (.I0(n1206), .I1(n1209), .I2(n1210), .O(n1211));
  LUT3 #(.INIT(8'h96)) lut_n1212 (.I0(n1185), .I1(n1193), .I2(n1194), .O(n1212));
  LUT3 #(.INIT(8'hE8)) lut_n1213 (.I0(n1203), .I1(n1211), .I2(n1212), .O(n1213));
  LUT3 #(.INIT(8'h96)) lut_n1214 (.I0(n1153), .I1(n1171), .I2(n1172), .O(n1214));
  LUT3 #(.INIT(8'hE8)) lut_n1215 (.I0(n1195), .I1(n1213), .I2(n1214), .O(n1215));
  LUT3 #(.INIT(8'h96)) lut_n1216 (.I0(x372), .I1(x373), .I2(x374), .O(n1216));
  LUT5 #(.INIT(32'h96696996)) lut_n1217 (.I0(x363), .I1(x364), .I2(x365), .I3(n1207), .I4(n1208), .O(n1217));
  LUT5 #(.INIT(32'hFF969600)) lut_n1218 (.I0(x369), .I1(x370), .I2(x371), .I3(n1216), .I4(n1217), .O(n1218));
  LUT3 #(.INIT(8'h96)) lut_n1219 (.I0(x378), .I1(x379), .I2(x380), .O(n1219));
  LUT5 #(.INIT(32'h96696996)) lut_n1220 (.I0(x369), .I1(x370), .I2(x371), .I3(n1216), .I4(n1217), .O(n1220));
  LUT5 #(.INIT(32'hFF969600)) lut_n1221 (.I0(x375), .I1(x376), .I2(x377), .I3(n1219), .I4(n1220), .O(n1221));
  LUT3 #(.INIT(8'h96)) lut_n1222 (.I0(n1206), .I1(n1209), .I2(n1210), .O(n1222));
  LUT3 #(.INIT(8'hE8)) lut_n1223 (.I0(n1218), .I1(n1221), .I2(n1222), .O(n1223));
  LUT3 #(.INIT(8'h96)) lut_n1224 (.I0(x384), .I1(x385), .I2(x386), .O(n1224));
  LUT5 #(.INIT(32'h96696996)) lut_n1225 (.I0(x375), .I1(x376), .I2(x377), .I3(n1219), .I4(n1220), .O(n1225));
  LUT5 #(.INIT(32'hFF969600)) lut_n1226 (.I0(x381), .I1(x382), .I2(x383), .I3(n1224), .I4(n1225), .O(n1226));
  LUT3 #(.INIT(8'h96)) lut_n1227 (.I0(x390), .I1(x391), .I2(x392), .O(n1227));
  LUT5 #(.INIT(32'h96696996)) lut_n1228 (.I0(x381), .I1(x382), .I2(x383), .I3(n1224), .I4(n1225), .O(n1228));
  LUT5 #(.INIT(32'hFF969600)) lut_n1229 (.I0(x387), .I1(x388), .I2(x389), .I3(n1227), .I4(n1228), .O(n1229));
  LUT3 #(.INIT(8'h96)) lut_n1230 (.I0(n1218), .I1(n1221), .I2(n1222), .O(n1230));
  LUT3 #(.INIT(8'hE8)) lut_n1231 (.I0(n1226), .I1(n1229), .I2(n1230), .O(n1231));
  LUT3 #(.INIT(8'h96)) lut_n1232 (.I0(n1203), .I1(n1211), .I2(n1212), .O(n1232));
  LUT3 #(.INIT(8'hE8)) lut_n1233 (.I0(n1223), .I1(n1231), .I2(n1232), .O(n1233));
  LUT3 #(.INIT(8'h96)) lut_n1234 (.I0(x396), .I1(x397), .I2(x398), .O(n1234));
  LUT5 #(.INIT(32'h96696996)) lut_n1235 (.I0(x387), .I1(x388), .I2(x389), .I3(n1227), .I4(n1228), .O(n1235));
  LUT5 #(.INIT(32'hFF969600)) lut_n1236 (.I0(x393), .I1(x394), .I2(x395), .I3(n1234), .I4(n1235), .O(n1236));
  LUT3 #(.INIT(8'h96)) lut_n1237 (.I0(x402), .I1(x403), .I2(x404), .O(n1237));
  LUT5 #(.INIT(32'h96696996)) lut_n1238 (.I0(x393), .I1(x394), .I2(x395), .I3(n1234), .I4(n1235), .O(n1238));
  LUT5 #(.INIT(32'hFF969600)) lut_n1239 (.I0(x399), .I1(x400), .I2(x401), .I3(n1237), .I4(n1238), .O(n1239));
  LUT3 #(.INIT(8'h96)) lut_n1240 (.I0(n1226), .I1(n1229), .I2(n1230), .O(n1240));
  LUT3 #(.INIT(8'hE8)) lut_n1241 (.I0(n1236), .I1(n1239), .I2(n1240), .O(n1241));
  LUT3 #(.INIT(8'h96)) lut_n1242 (.I0(x408), .I1(x409), .I2(x410), .O(n1242));
  LUT5 #(.INIT(32'h96696996)) lut_n1243 (.I0(x399), .I1(x400), .I2(x401), .I3(n1237), .I4(n1238), .O(n1243));
  LUT5 #(.INIT(32'hFF969600)) lut_n1244 (.I0(x405), .I1(x406), .I2(x407), .I3(n1242), .I4(n1243), .O(n1244));
  LUT3 #(.INIT(8'h96)) lut_n1245 (.I0(x414), .I1(x415), .I2(x416), .O(n1245));
  LUT5 #(.INIT(32'h96696996)) lut_n1246 (.I0(x405), .I1(x406), .I2(x407), .I3(n1242), .I4(n1243), .O(n1246));
  LUT5 #(.INIT(32'hFF969600)) lut_n1247 (.I0(x411), .I1(x412), .I2(x413), .I3(n1245), .I4(n1246), .O(n1247));
  LUT3 #(.INIT(8'h96)) lut_n1248 (.I0(n1236), .I1(n1239), .I2(n1240), .O(n1248));
  LUT3 #(.INIT(8'hE8)) lut_n1249 (.I0(n1244), .I1(n1247), .I2(n1248), .O(n1249));
  LUT3 #(.INIT(8'h96)) lut_n1250 (.I0(n1223), .I1(n1231), .I2(n1232), .O(n1250));
  LUT3 #(.INIT(8'hE8)) lut_n1251 (.I0(n1241), .I1(n1249), .I2(n1250), .O(n1251));
  LUT3 #(.INIT(8'h96)) lut_n1252 (.I0(n1195), .I1(n1213), .I2(n1214), .O(n1252));
  LUT3 #(.INIT(8'hE8)) lut_n1253 (.I0(n1233), .I1(n1251), .I2(n1252), .O(n1253));
  LUT3 #(.INIT(8'h96)) lut_n1254 (.I0(n1135), .I1(n1173), .I2(n1174), .O(n1254));
  LUT3 #(.INIT(8'h96)) lut_n1255 (.I0(x420), .I1(x421), .I2(x422), .O(n1255));
  LUT5 #(.INIT(32'h96696996)) lut_n1256 (.I0(x411), .I1(x412), .I2(x413), .I3(n1245), .I4(n1246), .O(n1256));
  LUT5 #(.INIT(32'hFF969600)) lut_n1257 (.I0(x417), .I1(x418), .I2(x419), .I3(n1255), .I4(n1256), .O(n1257));
  LUT3 #(.INIT(8'h96)) lut_n1258 (.I0(x426), .I1(x427), .I2(x428), .O(n1258));
  LUT5 #(.INIT(32'h96696996)) lut_n1259 (.I0(x417), .I1(x418), .I2(x419), .I3(n1255), .I4(n1256), .O(n1259));
  LUT5 #(.INIT(32'hFF969600)) lut_n1260 (.I0(x423), .I1(x424), .I2(x425), .I3(n1258), .I4(n1259), .O(n1260));
  LUT3 #(.INIT(8'h96)) lut_n1261 (.I0(n1244), .I1(n1247), .I2(n1248), .O(n1261));
  LUT3 #(.INIT(8'hE8)) lut_n1262 (.I0(n1257), .I1(n1260), .I2(n1261), .O(n1262));
  LUT3 #(.INIT(8'h96)) lut_n1263 (.I0(x432), .I1(x433), .I2(x434), .O(n1263));
  LUT5 #(.INIT(32'h96696996)) lut_n1264 (.I0(x423), .I1(x424), .I2(x425), .I3(n1258), .I4(n1259), .O(n1264));
  LUT5 #(.INIT(32'hFF969600)) lut_n1265 (.I0(x429), .I1(x430), .I2(x431), .I3(n1263), .I4(n1264), .O(n1265));
  LUT3 #(.INIT(8'h96)) lut_n1266 (.I0(x438), .I1(x439), .I2(x440), .O(n1266));
  LUT5 #(.INIT(32'h96696996)) lut_n1267 (.I0(x429), .I1(x430), .I2(x431), .I3(n1263), .I4(n1264), .O(n1267));
  LUT5 #(.INIT(32'hFF969600)) lut_n1268 (.I0(x435), .I1(x436), .I2(x437), .I3(n1266), .I4(n1267), .O(n1268));
  LUT3 #(.INIT(8'h96)) lut_n1269 (.I0(n1257), .I1(n1260), .I2(n1261), .O(n1269));
  LUT3 #(.INIT(8'hE8)) lut_n1270 (.I0(n1265), .I1(n1268), .I2(n1269), .O(n1270));
  LUT3 #(.INIT(8'h96)) lut_n1271 (.I0(n1241), .I1(n1249), .I2(n1250), .O(n1271));
  LUT3 #(.INIT(8'hE8)) lut_n1272 (.I0(n1262), .I1(n1270), .I2(n1271), .O(n1272));
  LUT3 #(.INIT(8'h96)) lut_n1273 (.I0(x444), .I1(x445), .I2(x446), .O(n1273));
  LUT5 #(.INIT(32'h96696996)) lut_n1274 (.I0(x435), .I1(x436), .I2(x437), .I3(n1266), .I4(n1267), .O(n1274));
  LUT5 #(.INIT(32'hFF969600)) lut_n1275 (.I0(x441), .I1(x442), .I2(x443), .I3(n1273), .I4(n1274), .O(n1275));
  LUT3 #(.INIT(8'h96)) lut_n1276 (.I0(x450), .I1(x451), .I2(x452), .O(n1276));
  LUT5 #(.INIT(32'h96696996)) lut_n1277 (.I0(x441), .I1(x442), .I2(x443), .I3(n1273), .I4(n1274), .O(n1277));
  LUT5 #(.INIT(32'hFF969600)) lut_n1278 (.I0(x447), .I1(x448), .I2(x449), .I3(n1276), .I4(n1277), .O(n1278));
  LUT3 #(.INIT(8'h96)) lut_n1279 (.I0(n1265), .I1(n1268), .I2(n1269), .O(n1279));
  LUT3 #(.INIT(8'hE8)) lut_n1280 (.I0(n1275), .I1(n1278), .I2(n1279), .O(n1280));
  LUT3 #(.INIT(8'h96)) lut_n1281 (.I0(x456), .I1(x457), .I2(x458), .O(n1281));
  LUT5 #(.INIT(32'h96696996)) lut_n1282 (.I0(x447), .I1(x448), .I2(x449), .I3(n1276), .I4(n1277), .O(n1282));
  LUT5 #(.INIT(32'hFF969600)) lut_n1283 (.I0(x453), .I1(x454), .I2(x455), .I3(n1281), .I4(n1282), .O(n1283));
  LUT3 #(.INIT(8'h96)) lut_n1284 (.I0(x462), .I1(x463), .I2(x464), .O(n1284));
  LUT5 #(.INIT(32'h96696996)) lut_n1285 (.I0(x453), .I1(x454), .I2(x455), .I3(n1281), .I4(n1282), .O(n1285));
  LUT5 #(.INIT(32'hFF969600)) lut_n1286 (.I0(x459), .I1(x460), .I2(x461), .I3(n1284), .I4(n1285), .O(n1286));
  LUT3 #(.INIT(8'h96)) lut_n1287 (.I0(n1275), .I1(n1278), .I2(n1279), .O(n1287));
  LUT3 #(.INIT(8'hE8)) lut_n1288 (.I0(n1283), .I1(n1286), .I2(n1287), .O(n1288));
  LUT3 #(.INIT(8'h96)) lut_n1289 (.I0(n1262), .I1(n1270), .I2(n1271), .O(n1289));
  LUT3 #(.INIT(8'hE8)) lut_n1290 (.I0(n1280), .I1(n1288), .I2(n1289), .O(n1290));
  LUT3 #(.INIT(8'h96)) lut_n1291 (.I0(n1233), .I1(n1251), .I2(n1252), .O(n1291));
  LUT3 #(.INIT(8'hE8)) lut_n1292 (.I0(n1272), .I1(n1290), .I2(n1291), .O(n1292));
  LUT3 #(.INIT(8'h96)) lut_n1293 (.I0(x468), .I1(x469), .I2(x470), .O(n1293));
  LUT5 #(.INIT(32'h96696996)) lut_n1294 (.I0(x459), .I1(x460), .I2(x461), .I3(n1284), .I4(n1285), .O(n1294));
  LUT5 #(.INIT(32'hFF969600)) lut_n1295 (.I0(x465), .I1(x466), .I2(x467), .I3(n1293), .I4(n1294), .O(n1295));
  LUT3 #(.INIT(8'h96)) lut_n1296 (.I0(x474), .I1(x475), .I2(x476), .O(n1296));
  LUT5 #(.INIT(32'h96696996)) lut_n1297 (.I0(x465), .I1(x466), .I2(x467), .I3(n1293), .I4(n1294), .O(n1297));
  LUT5 #(.INIT(32'hFF969600)) lut_n1298 (.I0(x471), .I1(x472), .I2(x473), .I3(n1296), .I4(n1297), .O(n1298));
  LUT3 #(.INIT(8'h96)) lut_n1299 (.I0(n1283), .I1(n1286), .I2(n1287), .O(n1299));
  LUT3 #(.INIT(8'hE8)) lut_n1300 (.I0(n1295), .I1(n1298), .I2(n1299), .O(n1300));
  LUT3 #(.INIT(8'h96)) lut_n1301 (.I0(x480), .I1(x481), .I2(x482), .O(n1301));
  LUT5 #(.INIT(32'h96696996)) lut_n1302 (.I0(x471), .I1(x472), .I2(x473), .I3(n1296), .I4(n1297), .O(n1302));
  LUT5 #(.INIT(32'hFF969600)) lut_n1303 (.I0(x477), .I1(x478), .I2(x479), .I3(n1301), .I4(n1302), .O(n1303));
  LUT3 #(.INIT(8'h96)) lut_n1304 (.I0(x486), .I1(x487), .I2(x488), .O(n1304));
  LUT5 #(.INIT(32'h96696996)) lut_n1305 (.I0(x477), .I1(x478), .I2(x479), .I3(n1301), .I4(n1302), .O(n1305));
  LUT5 #(.INIT(32'hFF969600)) lut_n1306 (.I0(x483), .I1(x484), .I2(x485), .I3(n1304), .I4(n1305), .O(n1306));
  LUT3 #(.INIT(8'h96)) lut_n1307 (.I0(n1295), .I1(n1298), .I2(n1299), .O(n1307));
  LUT3 #(.INIT(8'hE8)) lut_n1308 (.I0(n1303), .I1(n1306), .I2(n1307), .O(n1308));
  LUT3 #(.INIT(8'h96)) lut_n1309 (.I0(n1280), .I1(n1288), .I2(n1289), .O(n1309));
  LUT3 #(.INIT(8'h96)) lut_n1310 (.I0(x492), .I1(x493), .I2(x494), .O(n1310));
  LUT5 #(.INIT(32'h96696996)) lut_n1311 (.I0(x483), .I1(x484), .I2(x485), .I3(n1304), .I4(n1305), .O(n1311));
  LUT5 #(.INIT(32'hFF969600)) lut_n1312 (.I0(x489), .I1(x490), .I2(x491), .I3(n1310), .I4(n1311), .O(n1312));
  LUT3 #(.INIT(8'h96)) lut_n1313 (.I0(x498), .I1(x499), .I2(x500), .O(n1313));
  LUT5 #(.INIT(32'h96696996)) lut_n1314 (.I0(x489), .I1(x490), .I2(x491), .I3(n1310), .I4(n1311), .O(n1314));
  LUT5 #(.INIT(32'hFF969600)) lut_n1315 (.I0(x495), .I1(x496), .I2(x497), .I3(n1313), .I4(n1314), .O(n1315));
  LUT3 #(.INIT(8'h96)) lut_n1316 (.I0(n1303), .I1(n1306), .I2(n1307), .O(n1316));
  LUT3 #(.INIT(8'hE8)) lut_n1317 (.I0(n1312), .I1(n1315), .I2(n1316), .O(n1317));
  LUT3 #(.INIT(8'h96)) lut_n1318 (.I0(x501), .I1(x502), .I2(x503), .O(n1318));
  LUT3 #(.INIT(8'h96)) lut_n1319 (.I0(x504), .I1(x505), .I2(x506), .O(n1319));
  LUT5 #(.INIT(32'h96696996)) lut_n1320 (.I0(x495), .I1(x496), .I2(x497), .I3(n1313), .I4(n1314), .O(n1320));
  LUT3 #(.INIT(8'h96)) lut_n1321 (.I0(x507), .I1(x508), .I2(x509), .O(n1321));
  LUT3 #(.INIT(8'h96)) lut_n1322 (.I0(n1312), .I1(n1315), .I2(n1316), .O(n1322));
  LUT6 #(.INIT(64'hFFFEFEE8E8808000)) lut_n1323 (.I0(x510), .I1(n1318), .I2(n1319), .I3(n1320), .I4(n1321), .I5(n1322), .O(n1323));
  LUT3 #(.INIT(8'h96)) lut_n1324 (.I0(n1272), .I1(n1290), .I2(n1291), .O(n1324));
  LUT6 #(.INIT(64'hFFFEFEE8E8808000)) lut_n1325 (.I0(n1300), .I1(n1308), .I2(n1309), .I3(n1317), .I4(n1323), .I5(n1324), .O(n1325));
  LUT3 #(.INIT(8'h96)) lut_n1326 (.I0(n1097), .I1(n1175), .I2(n1176), .O(n1326));
  LUT6 #(.INIT(64'hFFFEFEE8E8808000)) lut_n1327 (.I0(n1215), .I1(n1253), .I2(n1254), .I3(n1292), .I4(n1325), .I5(n1326), .O(n1327));
  LUT6 #(.INIT(64'hFEEAEAA8EAA8A880)) lut_n1328 (.I0(n810), .I1(n888), .I2(n1018), .I3(n1019), .I4(n1177), .I5(n1327), .O(n1328));
  assign y0 = n1328;
endmodule
