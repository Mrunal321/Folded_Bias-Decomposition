`timescale 1ns/1ps
`default_nettype none

module tb_top;
  // 5025-bit input vector
  reg  [5024:0] x = 5025'b0;
  wire       y0;
  reg  [63:0] idx;

  // DUT instantiation
  top dut (
    .x0(x[0]), .x1(x[1]), .x2(x[2]), .x3(x[3]), .x4(x[4]), .x5(x[5]), .x6(x[6]), .x7(x[7]), .x8(x[8]), .x9(x[9]), .x10(x[10]), .x11(x[11]), .x12(x[12]), .x13(x[13]), .x14(x[14]), .x15(x[15]), .x16(x[16]), .x17(x[17]), .x18(x[18]), .x19(x[19]), .x20(x[20]), .x21(x[21]), .x22(x[22]), .x23(x[23]), .x24(x[24]), .x25(x[25]), .x26(x[26]), .x27(x[27]), .x28(x[28]), .x29(x[29]), .x30(x[30]), .x31(x[31]), .x32(x[32]), .x33(x[33]), .x34(x[34]), .x35(x[35]), .x36(x[36]), .x37(x[37]), .x38(x[38]), .x39(x[39]), .x40(x[40]), .x41(x[41]), .x42(x[42]), .x43(x[43]), .x44(x[44]), .x45(x[45]), .x46(x[46]), .x47(x[47]), .x48(x[48]), .x49(x[49]), .x50(x[50]), .x51(x[51]), .x52(x[52]), .x53(x[53]), .x54(x[54]), .x55(x[55]), .x56(x[56]), .x57(x[57]), .x58(x[58]), .x59(x[59]), .x60(x[60]), .x61(x[61]), .x62(x[62]), .x63(x[63]), .x64(x[64]), .x65(x[65]), .x66(x[66]), .x67(x[67]), .x68(x[68]), .x69(x[69]), .x70(x[70]), .x71(x[71]), .x72(x[72]), .x73(x[73]), .x74(x[74]), .x75(x[75]), .x76(x[76]), .x77(x[77]), .x78(x[78]), .x79(x[79]), .x80(x[80]), .x81(x[81]), .x82(x[82]), .x83(x[83]), .x84(x[84]), .x85(x[85]), .x86(x[86]), .x87(x[87]), .x88(x[88]), .x89(x[89]), .x90(x[90]), .x91(x[91]), .x92(x[92]), .x93(x[93]), .x94(x[94]), .x95(x[95]), .x96(x[96]), .x97(x[97]), .x98(x[98]), .x99(x[99]), .x100(x[100]), .x101(x[101]), .x102(x[102]), .x103(x[103]), .x104(x[104]), .x105(x[105]), .x106(x[106]), .x107(x[107]), .x108(x[108]), .x109(x[109]), .x110(x[110]), .x111(x[111]), .x112(x[112]), .x113(x[113]), .x114(x[114]), .x115(x[115]), .x116(x[116]), .x117(x[117]), .x118(x[118]), .x119(x[119]), .x120(x[120]), .x121(x[121]), .x122(x[122]), .x123(x[123]), .x124(x[124]), .x125(x[125]), .x126(x[126]), .x127(x[127]), .x128(x[128]), .x129(x[129]), .x130(x[130]), .x131(x[131]), .x132(x[132]), .x133(x[133]), .x134(x[134]), .x135(x[135]), .x136(x[136]), .x137(x[137]), .x138(x[138]), .x139(x[139]), .x140(x[140]), .x141(x[141]), .x142(x[142]), .x143(x[143]), .x144(x[144]), .x145(x[145]), .x146(x[146]), .x147(x[147]), .x148(x[148]), .x149(x[149]), .x150(x[150]), .x151(x[151]), .x152(x[152]), .x153(x[153]), .x154(x[154]), .x155(x[155]), .x156(x[156]), .x157(x[157]), .x158(x[158]), .x159(x[159]), .x160(x[160]), .x161(x[161]), .x162(x[162]), .x163(x[163]), .x164(x[164]), .x165(x[165]), .x166(x[166]), .x167(x[167]), .x168(x[168]), .x169(x[169]), .x170(x[170]), .x171(x[171]), .x172(x[172]), .x173(x[173]), .x174(x[174]), .x175(x[175]), .x176(x[176]), .x177(x[177]), .x178(x[178]), .x179(x[179]), .x180(x[180]), .x181(x[181]), .x182(x[182]), .x183(x[183]), .x184(x[184]), .x185(x[185]), .x186(x[186]), .x187(x[187]), .x188(x[188]), .x189(x[189]), .x190(x[190]), .x191(x[191]), .x192(x[192]), .x193(x[193]), .x194(x[194]), .x195(x[195]), .x196(x[196]), .x197(x[197]), .x198(x[198]), .x199(x[199]), .x200(x[200]), .x201(x[201]), .x202(x[202]), .x203(x[203]), .x204(x[204]), .x205(x[205]), .x206(x[206]), .x207(x[207]), .x208(x[208]), .x209(x[209]), .x210(x[210]), .x211(x[211]), .x212(x[212]), .x213(x[213]), .x214(x[214]), .x215(x[215]), .x216(x[216]), .x217(x[217]), .x218(x[218]), .x219(x[219]), .x220(x[220]), .x221(x[221]), .x222(x[222]), .x223(x[223]), .x224(x[224]), .x225(x[225]), .x226(x[226]), .x227(x[227]), .x228(x[228]), .x229(x[229]), .x230(x[230]), .x231(x[231]), .x232(x[232]), .x233(x[233]), .x234(x[234]), .x235(x[235]), .x236(x[236]), .x237(x[237]), .x238(x[238]), .x239(x[239]), .x240(x[240]), .x241(x[241]), .x242(x[242]), .x243(x[243]), .x244(x[244]), .x245(x[245]), .x246(x[246]), .x247(x[247]), .x248(x[248]), .x249(x[249]), .x250(x[250]), .x251(x[251]), .x252(x[252]), .x253(x[253]), .x254(x[254]), .x255(x[255]), .x256(x[256]), .x257(x[257]), .x258(x[258]), .x259(x[259]), .x260(x[260]), .x261(x[261]), .x262(x[262]), .x263(x[263]), .x264(x[264]), .x265(x[265]), .x266(x[266]), .x267(x[267]), .x268(x[268]), .x269(x[269]), .x270(x[270]), .x271(x[271]), .x272(x[272]), .x273(x[273]), .x274(x[274]), .x275(x[275]), .x276(x[276]), .x277(x[277]), .x278(x[278]), .x279(x[279]), .x280(x[280]), .x281(x[281]), .x282(x[282]), .x283(x[283]), .x284(x[284]), .x285(x[285]), .x286(x[286]), .x287(x[287]), .x288(x[288]), .x289(x[289]), .x290(x[290]), .x291(x[291]), .x292(x[292]), .x293(x[293]), .x294(x[294]), .x295(x[295]), .x296(x[296]), .x297(x[297]), .x298(x[298]), .x299(x[299]), .x300(x[300]), .x301(x[301]), .x302(x[302]), .x303(x[303]), .x304(x[304]), .x305(x[305]), .x306(x[306]), .x307(x[307]), .x308(x[308]), .x309(x[309]), .x310(x[310]), .x311(x[311]), .x312(x[312]), .x313(x[313]), .x314(x[314]), .x315(x[315]), .x316(x[316]), .x317(x[317]), .x318(x[318]), .x319(x[319]), .x320(x[320]), .x321(x[321]), .x322(x[322]), .x323(x[323]), .x324(x[324]), .x325(x[325]), .x326(x[326]), .x327(x[327]), .x328(x[328]), .x329(x[329]), .x330(x[330]), .x331(x[331]), .x332(x[332]), .x333(x[333]), .x334(x[334]), .x335(x[335]), .x336(x[336]), .x337(x[337]), .x338(x[338]), .x339(x[339]), .x340(x[340]), .x341(x[341]), .x342(x[342]), .x343(x[343]), .x344(x[344]), .x345(x[345]), .x346(x[346]), .x347(x[347]), .x348(x[348]), .x349(x[349]), .x350(x[350]), .x351(x[351]), .x352(x[352]), .x353(x[353]), .x354(x[354]), .x355(x[355]), .x356(x[356]), .x357(x[357]), .x358(x[358]), .x359(x[359]), .x360(x[360]), .x361(x[361]), .x362(x[362]), .x363(x[363]), .x364(x[364]), .x365(x[365]), .x366(x[366]), .x367(x[367]), .x368(x[368]), .x369(x[369]), .x370(x[370]), .x371(x[371]), .x372(x[372]), .x373(x[373]), .x374(x[374]), .x375(x[375]), .x376(x[376]), .x377(x[377]), .x378(x[378]), .x379(x[379]), .x380(x[380]), .x381(x[381]), .x382(x[382]), .x383(x[383]), .x384(x[384]), .x385(x[385]), .x386(x[386]), .x387(x[387]), .x388(x[388]), .x389(x[389]), .x390(x[390]), .x391(x[391]), .x392(x[392]), .x393(x[393]), .x394(x[394]), .x395(x[395]), .x396(x[396]), .x397(x[397]), .x398(x[398]), .x399(x[399]), .x400(x[400]), .x401(x[401]), .x402(x[402]), .x403(x[403]), .x404(x[404]), .x405(x[405]), .x406(x[406]), .x407(x[407]), .x408(x[408]), .x409(x[409]), .x410(x[410]), .x411(x[411]), .x412(x[412]), .x413(x[413]), .x414(x[414]), .x415(x[415]), .x416(x[416]), .x417(x[417]), .x418(x[418]), .x419(x[419]), .x420(x[420]), .x421(x[421]), .x422(x[422]), .x423(x[423]), .x424(x[424]), .x425(x[425]), .x426(x[426]), .x427(x[427]), .x428(x[428]), .x429(x[429]), .x430(x[430]), .x431(x[431]), .x432(x[432]), .x433(x[433]), .x434(x[434]), .x435(x[435]), .x436(x[436]), .x437(x[437]), .x438(x[438]), .x439(x[439]), .x440(x[440]), .x441(x[441]), .x442(x[442]), .x443(x[443]), .x444(x[444]), .x445(x[445]), .x446(x[446]), .x447(x[447]), .x448(x[448]), .x449(x[449]), .x450(x[450]), .x451(x[451]), .x452(x[452]), .x453(x[453]), .x454(x[454]), .x455(x[455]), .x456(x[456]), .x457(x[457]), .x458(x[458]), .x459(x[459]), .x460(x[460]), .x461(x[461]), .x462(x[462]), .x463(x[463]), .x464(x[464]), .x465(x[465]), .x466(x[466]), .x467(x[467]), .x468(x[468]), .x469(x[469]), .x470(x[470]), .x471(x[471]), .x472(x[472]), .x473(x[473]), .x474(x[474]), .x475(x[475]), .x476(x[476]), .x477(x[477]), .x478(x[478]), .x479(x[479]), .x480(x[480]), .x481(x[481]), .x482(x[482]), .x483(x[483]), .x484(x[484]), .x485(x[485]), .x486(x[486]), .x487(x[487]), .x488(x[488]), .x489(x[489]), .x490(x[490]), .x491(x[491]), .x492(x[492]), .x493(x[493]), .x494(x[494]), .x495(x[495]), .x496(x[496]), .x497(x[497]), .x498(x[498]), .x499(x[499]), .x500(x[500]), .x501(x[501]), .x502(x[502]), .x503(x[503]), .x504(x[504]), .x505(x[505]), .x506(x[506]), .x507(x[507]), .x508(x[508]), .x509(x[509]), .x510(x[510]), .x511(x[511]), .x512(x[512]), .x513(x[513]), .x514(x[514]), .x515(x[515]), .x516(x[516]), .x517(x[517]), .x518(x[518]), .x519(x[519]), .x520(x[520]), .x521(x[521]), .x522(x[522]), .x523(x[523]), .x524(x[524]), .x525(x[525]), .x526(x[526]), .x527(x[527]), .x528(x[528]), .x529(x[529]), .x530(x[530]), .x531(x[531]), .x532(x[532]), .x533(x[533]), .x534(x[534]), .x535(x[535]), .x536(x[536]), .x537(x[537]), .x538(x[538]), .x539(x[539]), .x540(x[540]), .x541(x[541]), .x542(x[542]), .x543(x[543]), .x544(x[544]), .x545(x[545]), .x546(x[546]), .x547(x[547]), .x548(x[548]), .x549(x[549]), .x550(x[550]), .x551(x[551]), .x552(x[552]), .x553(x[553]), .x554(x[554]), .x555(x[555]), .x556(x[556]), .x557(x[557]), .x558(x[558]), .x559(x[559]), .x560(x[560]), .x561(x[561]), .x562(x[562]), .x563(x[563]), .x564(x[564]), .x565(x[565]), .x566(x[566]), .x567(x[567]), .x568(x[568]), .x569(x[569]), .x570(x[570]), .x571(x[571]), .x572(x[572]), .x573(x[573]), .x574(x[574]), .x575(x[575]), .x576(x[576]), .x577(x[577]), .x578(x[578]), .x579(x[579]), .x580(x[580]), .x581(x[581]), .x582(x[582]), .x583(x[583]), .x584(x[584]), .x585(x[585]), .x586(x[586]), .x587(x[587]), .x588(x[588]), .x589(x[589]), .x590(x[590]), .x591(x[591]), .x592(x[592]), .x593(x[593]), .x594(x[594]), .x595(x[595]), .x596(x[596]), .x597(x[597]), .x598(x[598]), .x599(x[599]), .x600(x[600]), .x601(x[601]), .x602(x[602]), .x603(x[603]), .x604(x[604]), .x605(x[605]), .x606(x[606]), .x607(x[607]), .x608(x[608]), .x609(x[609]), .x610(x[610]), .x611(x[611]), .x612(x[612]), .x613(x[613]), .x614(x[614]), .x615(x[615]), .x616(x[616]), .x617(x[617]), .x618(x[618]), .x619(x[619]), .x620(x[620]), .x621(x[621]), .x622(x[622]), .x623(x[623]), .x624(x[624]), .x625(x[625]), .x626(x[626]), .x627(x[627]), .x628(x[628]), .x629(x[629]), .x630(x[630]), .x631(x[631]), .x632(x[632]), .x633(x[633]), .x634(x[634]), .x635(x[635]), .x636(x[636]), .x637(x[637]), .x638(x[638]), .x639(x[639]), .x640(x[640]), .x641(x[641]), .x642(x[642]), .x643(x[643]), .x644(x[644]), .x645(x[645]), .x646(x[646]), .x647(x[647]), .x648(x[648]), .x649(x[649]), .x650(x[650]), .x651(x[651]), .x652(x[652]), .x653(x[653]), .x654(x[654]), .x655(x[655]), .x656(x[656]), .x657(x[657]), .x658(x[658]), .x659(x[659]), .x660(x[660]), .x661(x[661]), .x662(x[662]), .x663(x[663]), .x664(x[664]), .x665(x[665]), .x666(x[666]), .x667(x[667]), .x668(x[668]), .x669(x[669]), .x670(x[670]), .x671(x[671]), .x672(x[672]), .x673(x[673]), .x674(x[674]), .x675(x[675]), .x676(x[676]), .x677(x[677]), .x678(x[678]), .x679(x[679]), .x680(x[680]), .x681(x[681]), .x682(x[682]), .x683(x[683]), .x684(x[684]), .x685(x[685]), .x686(x[686]), .x687(x[687]), .x688(x[688]), .x689(x[689]), .x690(x[690]), .x691(x[691]), .x692(x[692]), .x693(x[693]), .x694(x[694]), .x695(x[695]), .x696(x[696]), .x697(x[697]), .x698(x[698]), .x699(x[699]), .x700(x[700]), .x701(x[701]), .x702(x[702]), .x703(x[703]), .x704(x[704]), .x705(x[705]), .x706(x[706]), .x707(x[707]), .x708(x[708]), .x709(x[709]), .x710(x[710]), .x711(x[711]), .x712(x[712]), .x713(x[713]), .x714(x[714]), .x715(x[715]), .x716(x[716]), .x717(x[717]), .x718(x[718]), .x719(x[719]), .x720(x[720]), .x721(x[721]), .x722(x[722]), .x723(x[723]), .x724(x[724]), .x725(x[725]), .x726(x[726]), .x727(x[727]), .x728(x[728]), .x729(x[729]), .x730(x[730]), .x731(x[731]), .x732(x[732]), .x733(x[733]), .x734(x[734]), .x735(x[735]), .x736(x[736]), .x737(x[737]), .x738(x[738]), .x739(x[739]), .x740(x[740]), .x741(x[741]), .x742(x[742]), .x743(x[743]), .x744(x[744]), .x745(x[745]), .x746(x[746]), .x747(x[747]), .x748(x[748]), .x749(x[749]), .x750(x[750]), .x751(x[751]), .x752(x[752]), .x753(x[753]), .x754(x[754]), .x755(x[755]), .x756(x[756]), .x757(x[757]), .x758(x[758]), .x759(x[759]), .x760(x[760]), .x761(x[761]), .x762(x[762]), .x763(x[763]), .x764(x[764]), .x765(x[765]), .x766(x[766]), .x767(x[767]), .x768(x[768]), .x769(x[769]), .x770(x[770]), .x771(x[771]), .x772(x[772]), .x773(x[773]), .x774(x[774]), .x775(x[775]), .x776(x[776]), .x777(x[777]), .x778(x[778]), .x779(x[779]), .x780(x[780]), .x781(x[781]), .x782(x[782]), .x783(x[783]), .x784(x[784]), .x785(x[785]), .x786(x[786]), .x787(x[787]), .x788(x[788]), .x789(x[789]), .x790(x[790]), .x791(x[791]), .x792(x[792]), .x793(x[793]), .x794(x[794]), .x795(x[795]), .x796(x[796]), .x797(x[797]), .x798(x[798]), .x799(x[799]), .x800(x[800]), .x801(x[801]), .x802(x[802]), .x803(x[803]), .x804(x[804]), .x805(x[805]), .x806(x[806]), .x807(x[807]), .x808(x[808]), .x809(x[809]), .x810(x[810]), .x811(x[811]), .x812(x[812]), .x813(x[813]), .x814(x[814]), .x815(x[815]), .x816(x[816]), .x817(x[817]), .x818(x[818]), .x819(x[819]), .x820(x[820]), .x821(x[821]), .x822(x[822]), .x823(x[823]), .x824(x[824]), .x825(x[825]), .x826(x[826]), .x827(x[827]), .x828(x[828]), .x829(x[829]), .x830(x[830]), .x831(x[831]), .x832(x[832]), .x833(x[833]), .x834(x[834]), .x835(x[835]), .x836(x[836]), .x837(x[837]), .x838(x[838]), .x839(x[839]), .x840(x[840]), .x841(x[841]), .x842(x[842]), .x843(x[843]), .x844(x[844]), .x845(x[845]), .x846(x[846]), .x847(x[847]), .x848(x[848]), .x849(x[849]), .x850(x[850]), .x851(x[851]), .x852(x[852]), .x853(x[853]), .x854(x[854]), .x855(x[855]), .x856(x[856]), .x857(x[857]), .x858(x[858]), .x859(x[859]), .x860(x[860]), .x861(x[861]), .x862(x[862]), .x863(x[863]), .x864(x[864]), .x865(x[865]), .x866(x[866]), .x867(x[867]), .x868(x[868]), .x869(x[869]), .x870(x[870]), .x871(x[871]), .x872(x[872]), .x873(x[873]), .x874(x[874]), .x875(x[875]), .x876(x[876]), .x877(x[877]), .x878(x[878]), .x879(x[879]), .x880(x[880]), .x881(x[881]), .x882(x[882]), .x883(x[883]), .x884(x[884]), .x885(x[885]), .x886(x[886]), .x887(x[887]), .x888(x[888]), .x889(x[889]), .x890(x[890]), .x891(x[891]), .x892(x[892]), .x893(x[893]), .x894(x[894]), .x895(x[895]), .x896(x[896]), .x897(x[897]), .x898(x[898]), .x899(x[899]), .x900(x[900]), .x901(x[901]), .x902(x[902]), .x903(x[903]), .x904(x[904]), .x905(x[905]), .x906(x[906]), .x907(x[907]), .x908(x[908]), .x909(x[909]), .x910(x[910]), .x911(x[911]), .x912(x[912]), .x913(x[913]), .x914(x[914]), .x915(x[915]), .x916(x[916]), .x917(x[917]), .x918(x[918]), .x919(x[919]), .x920(x[920]), .x921(x[921]), .x922(x[922]), .x923(x[923]), .x924(x[924]), .x925(x[925]), .x926(x[926]), .x927(x[927]), .x928(x[928]), .x929(x[929]), .x930(x[930]), .x931(x[931]), .x932(x[932]), .x933(x[933]), .x934(x[934]), .x935(x[935]), .x936(x[936]), .x937(x[937]), .x938(x[938]), .x939(x[939]), .x940(x[940]), .x941(x[941]), .x942(x[942]), .x943(x[943]), .x944(x[944]), .x945(x[945]), .x946(x[946]), .x947(x[947]), .x948(x[948]), .x949(x[949]), .x950(x[950]), .x951(x[951]), .x952(x[952]), .x953(x[953]), .x954(x[954]), .x955(x[955]), .x956(x[956]), .x957(x[957]), .x958(x[958]), .x959(x[959]), .x960(x[960]), .x961(x[961]), .x962(x[962]), .x963(x[963]), .x964(x[964]), .x965(x[965]), .x966(x[966]), .x967(x[967]), .x968(x[968]), .x969(x[969]), .x970(x[970]), .x971(x[971]), .x972(x[972]), .x973(x[973]), .x974(x[974]), .x975(x[975]), .x976(x[976]), .x977(x[977]), .x978(x[978]), .x979(x[979]), .x980(x[980]), .x981(x[981]), .x982(x[982]), .x983(x[983]), .x984(x[984]), .x985(x[985]), .x986(x[986]), .x987(x[987]), .x988(x[988]), .x989(x[989]), .x990(x[990]), .x991(x[991]), .x992(x[992]), .x993(x[993]), .x994(x[994]), .x995(x[995]), .x996(x[996]), .x997(x[997]), .x998(x[998]), .x999(x[999]), .x1000(x[1000]), .x1001(x[1001]), .x1002(x[1002]), .x1003(x[1003]), .x1004(x[1004]), .x1005(x[1005]), .x1006(x[1006]), .x1007(x[1007]), .x1008(x[1008]), .x1009(x[1009]), .x1010(x[1010]), .x1011(x[1011]), .x1012(x[1012]), .x1013(x[1013]), .x1014(x[1014]), .x1015(x[1015]), .x1016(x[1016]), .x1017(x[1017]), .x1018(x[1018]), .x1019(x[1019]), .x1020(x[1020]), .x1021(x[1021]), .x1022(x[1022]), .x1023(x[1023]), .x1024(x[1024]), .x1025(x[1025]), .x1026(x[1026]), .x1027(x[1027]), .x1028(x[1028]), .x1029(x[1029]), .x1030(x[1030]), .x1031(x[1031]), .x1032(x[1032]), .x1033(x[1033]), .x1034(x[1034]), .x1035(x[1035]), .x1036(x[1036]), .x1037(x[1037]), .x1038(x[1038]), .x1039(x[1039]), .x1040(x[1040]), .x1041(x[1041]), .x1042(x[1042]), .x1043(x[1043]), .x1044(x[1044]), .x1045(x[1045]), .x1046(x[1046]), .x1047(x[1047]), .x1048(x[1048]), .x1049(x[1049]), .x1050(x[1050]), .x1051(x[1051]), .x1052(x[1052]), .x1053(x[1053]), .x1054(x[1054]), .x1055(x[1055]), .x1056(x[1056]), .x1057(x[1057]), .x1058(x[1058]), .x1059(x[1059]), .x1060(x[1060]), .x1061(x[1061]), .x1062(x[1062]), .x1063(x[1063]), .x1064(x[1064]), .x1065(x[1065]), .x1066(x[1066]), .x1067(x[1067]), .x1068(x[1068]), .x1069(x[1069]), .x1070(x[1070]), .x1071(x[1071]), .x1072(x[1072]), .x1073(x[1073]), .x1074(x[1074]), .x1075(x[1075]), .x1076(x[1076]), .x1077(x[1077]), .x1078(x[1078]), .x1079(x[1079]), .x1080(x[1080]), .x1081(x[1081]), .x1082(x[1082]), .x1083(x[1083]), .x1084(x[1084]), .x1085(x[1085]), .x1086(x[1086]), .x1087(x[1087]), .x1088(x[1088]), .x1089(x[1089]), .x1090(x[1090]), .x1091(x[1091]), .x1092(x[1092]), .x1093(x[1093]), .x1094(x[1094]), .x1095(x[1095]), .x1096(x[1096]), .x1097(x[1097]), .x1098(x[1098]), .x1099(x[1099]), .x1100(x[1100]), .x1101(x[1101]), .x1102(x[1102]), .x1103(x[1103]), .x1104(x[1104]), .x1105(x[1105]), .x1106(x[1106]), .x1107(x[1107]), .x1108(x[1108]), .x1109(x[1109]), .x1110(x[1110]), .x1111(x[1111]), .x1112(x[1112]), .x1113(x[1113]), .x1114(x[1114]), .x1115(x[1115]), .x1116(x[1116]), .x1117(x[1117]), .x1118(x[1118]), .x1119(x[1119]), .x1120(x[1120]), .x1121(x[1121]), .x1122(x[1122]), .x1123(x[1123]), .x1124(x[1124]), .x1125(x[1125]), .x1126(x[1126]), .x1127(x[1127]), .x1128(x[1128]), .x1129(x[1129]), .x1130(x[1130]), .x1131(x[1131]), .x1132(x[1132]), .x1133(x[1133]), .x1134(x[1134]), .x1135(x[1135]), .x1136(x[1136]), .x1137(x[1137]), .x1138(x[1138]), .x1139(x[1139]), .x1140(x[1140]), .x1141(x[1141]), .x1142(x[1142]), .x1143(x[1143]), .x1144(x[1144]), .x1145(x[1145]), .x1146(x[1146]), .x1147(x[1147]), .x1148(x[1148]), .x1149(x[1149]), .x1150(x[1150]), .x1151(x[1151]), .x1152(x[1152]), .x1153(x[1153]), .x1154(x[1154]), .x1155(x[1155]), .x1156(x[1156]), .x1157(x[1157]), .x1158(x[1158]), .x1159(x[1159]), .x1160(x[1160]), .x1161(x[1161]), .x1162(x[1162]), .x1163(x[1163]), .x1164(x[1164]), .x1165(x[1165]), .x1166(x[1166]), .x1167(x[1167]), .x1168(x[1168]), .x1169(x[1169]), .x1170(x[1170]), .x1171(x[1171]), .x1172(x[1172]), .x1173(x[1173]), .x1174(x[1174]), .x1175(x[1175]), .x1176(x[1176]), .x1177(x[1177]), .x1178(x[1178]), .x1179(x[1179]), .x1180(x[1180]), .x1181(x[1181]), .x1182(x[1182]), .x1183(x[1183]), .x1184(x[1184]), .x1185(x[1185]), .x1186(x[1186]), .x1187(x[1187]), .x1188(x[1188]), .x1189(x[1189]), .x1190(x[1190]), .x1191(x[1191]), .x1192(x[1192]), .x1193(x[1193]), .x1194(x[1194]), .x1195(x[1195]), .x1196(x[1196]), .x1197(x[1197]), .x1198(x[1198]), .x1199(x[1199]), .x1200(x[1200]), .x1201(x[1201]), .x1202(x[1202]), .x1203(x[1203]), .x1204(x[1204]), .x1205(x[1205]), .x1206(x[1206]), .x1207(x[1207]), .x1208(x[1208]), .x1209(x[1209]), .x1210(x[1210]), .x1211(x[1211]), .x1212(x[1212]), .x1213(x[1213]), .x1214(x[1214]), .x1215(x[1215]), .x1216(x[1216]), .x1217(x[1217]), .x1218(x[1218]), .x1219(x[1219]), .x1220(x[1220]), .x1221(x[1221]), .x1222(x[1222]), .x1223(x[1223]), .x1224(x[1224]), .x1225(x[1225]), .x1226(x[1226]), .x1227(x[1227]), .x1228(x[1228]), .x1229(x[1229]), .x1230(x[1230]), .x1231(x[1231]), .x1232(x[1232]), .x1233(x[1233]), .x1234(x[1234]), .x1235(x[1235]), .x1236(x[1236]), .x1237(x[1237]), .x1238(x[1238]), .x1239(x[1239]), .x1240(x[1240]), .x1241(x[1241]), .x1242(x[1242]), .x1243(x[1243]), .x1244(x[1244]), .x1245(x[1245]), .x1246(x[1246]), .x1247(x[1247]), .x1248(x[1248]), .x1249(x[1249]), .x1250(x[1250]), .x1251(x[1251]), .x1252(x[1252]), .x1253(x[1253]), .x1254(x[1254]), .x1255(x[1255]), .x1256(x[1256]), .x1257(x[1257]), .x1258(x[1258]), .x1259(x[1259]), .x1260(x[1260]), .x1261(x[1261]), .x1262(x[1262]), .x1263(x[1263]), .x1264(x[1264]), .x1265(x[1265]), .x1266(x[1266]), .x1267(x[1267]), .x1268(x[1268]), .x1269(x[1269]), .x1270(x[1270]), .x1271(x[1271]), .x1272(x[1272]), .x1273(x[1273]), .x1274(x[1274]), .x1275(x[1275]), .x1276(x[1276]), .x1277(x[1277]), .x1278(x[1278]), .x1279(x[1279]), .x1280(x[1280]), .x1281(x[1281]), .x1282(x[1282]), .x1283(x[1283]), .x1284(x[1284]), .x1285(x[1285]), .x1286(x[1286]), .x1287(x[1287]), .x1288(x[1288]), .x1289(x[1289]), .x1290(x[1290]), .x1291(x[1291]), .x1292(x[1292]), .x1293(x[1293]), .x1294(x[1294]), .x1295(x[1295]), .x1296(x[1296]), .x1297(x[1297]), .x1298(x[1298]), .x1299(x[1299]), .x1300(x[1300]), .x1301(x[1301]), .x1302(x[1302]), .x1303(x[1303]), .x1304(x[1304]), .x1305(x[1305]), .x1306(x[1306]), .x1307(x[1307]), .x1308(x[1308]), .x1309(x[1309]), .x1310(x[1310]), .x1311(x[1311]), .x1312(x[1312]), .x1313(x[1313]), .x1314(x[1314]), .x1315(x[1315]), .x1316(x[1316]), .x1317(x[1317]), .x1318(x[1318]), .x1319(x[1319]), .x1320(x[1320]), .x1321(x[1321]), .x1322(x[1322]), .x1323(x[1323]), .x1324(x[1324]), .x1325(x[1325]), .x1326(x[1326]), .x1327(x[1327]), .x1328(x[1328]), .x1329(x[1329]), .x1330(x[1330]), .x1331(x[1331]), .x1332(x[1332]), .x1333(x[1333]), .x1334(x[1334]), .x1335(x[1335]), .x1336(x[1336]), .x1337(x[1337]), .x1338(x[1338]), .x1339(x[1339]), .x1340(x[1340]), .x1341(x[1341]), .x1342(x[1342]), .x1343(x[1343]), .x1344(x[1344]), .x1345(x[1345]), .x1346(x[1346]), .x1347(x[1347]), .x1348(x[1348]), .x1349(x[1349]), .x1350(x[1350]), .x1351(x[1351]), .x1352(x[1352]), .x1353(x[1353]), .x1354(x[1354]), .x1355(x[1355]), .x1356(x[1356]), .x1357(x[1357]), .x1358(x[1358]), .x1359(x[1359]), .x1360(x[1360]), .x1361(x[1361]), .x1362(x[1362]), .x1363(x[1363]), .x1364(x[1364]), .x1365(x[1365]), .x1366(x[1366]), .x1367(x[1367]), .x1368(x[1368]), .x1369(x[1369]), .x1370(x[1370]), .x1371(x[1371]), .x1372(x[1372]), .x1373(x[1373]), .x1374(x[1374]), .x1375(x[1375]), .x1376(x[1376]), .x1377(x[1377]), .x1378(x[1378]), .x1379(x[1379]), .x1380(x[1380]), .x1381(x[1381]), .x1382(x[1382]), .x1383(x[1383]), .x1384(x[1384]), .x1385(x[1385]), .x1386(x[1386]), .x1387(x[1387]), .x1388(x[1388]), .x1389(x[1389]), .x1390(x[1390]), .x1391(x[1391]), .x1392(x[1392]), .x1393(x[1393]), .x1394(x[1394]), .x1395(x[1395]), .x1396(x[1396]), .x1397(x[1397]), .x1398(x[1398]), .x1399(x[1399]), .x1400(x[1400]), .x1401(x[1401]), .x1402(x[1402]), .x1403(x[1403]), .x1404(x[1404]), .x1405(x[1405]), .x1406(x[1406]), .x1407(x[1407]), .x1408(x[1408]), .x1409(x[1409]), .x1410(x[1410]), .x1411(x[1411]), .x1412(x[1412]), .x1413(x[1413]), .x1414(x[1414]), .x1415(x[1415]), .x1416(x[1416]), .x1417(x[1417]), .x1418(x[1418]), .x1419(x[1419]), .x1420(x[1420]), .x1421(x[1421]), .x1422(x[1422]), .x1423(x[1423]), .x1424(x[1424]), .x1425(x[1425]), .x1426(x[1426]), .x1427(x[1427]), .x1428(x[1428]), .x1429(x[1429]), .x1430(x[1430]), .x1431(x[1431]), .x1432(x[1432]), .x1433(x[1433]), .x1434(x[1434]), .x1435(x[1435]), .x1436(x[1436]), .x1437(x[1437]), .x1438(x[1438]), .x1439(x[1439]), .x1440(x[1440]), .x1441(x[1441]), .x1442(x[1442]), .x1443(x[1443]), .x1444(x[1444]), .x1445(x[1445]), .x1446(x[1446]), .x1447(x[1447]), .x1448(x[1448]), .x1449(x[1449]), .x1450(x[1450]), .x1451(x[1451]), .x1452(x[1452]), .x1453(x[1453]), .x1454(x[1454]), .x1455(x[1455]), .x1456(x[1456]), .x1457(x[1457]), .x1458(x[1458]), .x1459(x[1459]), .x1460(x[1460]), .x1461(x[1461]), .x1462(x[1462]), .x1463(x[1463]), .x1464(x[1464]), .x1465(x[1465]), .x1466(x[1466]), .x1467(x[1467]), .x1468(x[1468]), .x1469(x[1469]), .x1470(x[1470]), .x1471(x[1471]), .x1472(x[1472]), .x1473(x[1473]), .x1474(x[1474]), .x1475(x[1475]), .x1476(x[1476]), .x1477(x[1477]), .x1478(x[1478]), .x1479(x[1479]), .x1480(x[1480]), .x1481(x[1481]), .x1482(x[1482]), .x1483(x[1483]), .x1484(x[1484]), .x1485(x[1485]), .x1486(x[1486]), .x1487(x[1487]), .x1488(x[1488]), .x1489(x[1489]), .x1490(x[1490]), .x1491(x[1491]), .x1492(x[1492]), .x1493(x[1493]), .x1494(x[1494]), .x1495(x[1495]), .x1496(x[1496]), .x1497(x[1497]), .x1498(x[1498]), .x1499(x[1499]), .x1500(x[1500]), .x1501(x[1501]), .x1502(x[1502]), .x1503(x[1503]), .x1504(x[1504]), .x1505(x[1505]), .x1506(x[1506]), .x1507(x[1507]), .x1508(x[1508]), .x1509(x[1509]), .x1510(x[1510]), .x1511(x[1511]), .x1512(x[1512]), .x1513(x[1513]), .x1514(x[1514]), .x1515(x[1515]), .x1516(x[1516]), .x1517(x[1517]), .x1518(x[1518]), .x1519(x[1519]), .x1520(x[1520]), .x1521(x[1521]), .x1522(x[1522]), .x1523(x[1523]), .x1524(x[1524]), .x1525(x[1525]), .x1526(x[1526]), .x1527(x[1527]), .x1528(x[1528]), .x1529(x[1529]), .x1530(x[1530]), .x1531(x[1531]), .x1532(x[1532]), .x1533(x[1533]), .x1534(x[1534]), .x1535(x[1535]), .x1536(x[1536]), .x1537(x[1537]), .x1538(x[1538]), .x1539(x[1539]), .x1540(x[1540]), .x1541(x[1541]), .x1542(x[1542]), .x1543(x[1543]), .x1544(x[1544]), .x1545(x[1545]), .x1546(x[1546]), .x1547(x[1547]), .x1548(x[1548]), .x1549(x[1549]), .x1550(x[1550]), .x1551(x[1551]), .x1552(x[1552]), .x1553(x[1553]), .x1554(x[1554]), .x1555(x[1555]), .x1556(x[1556]), .x1557(x[1557]), .x1558(x[1558]), .x1559(x[1559]), .x1560(x[1560]), .x1561(x[1561]), .x1562(x[1562]), .x1563(x[1563]), .x1564(x[1564]), .x1565(x[1565]), .x1566(x[1566]), .x1567(x[1567]), .x1568(x[1568]), .x1569(x[1569]), .x1570(x[1570]), .x1571(x[1571]), .x1572(x[1572]), .x1573(x[1573]), .x1574(x[1574]), .x1575(x[1575]), .x1576(x[1576]), .x1577(x[1577]), .x1578(x[1578]), .x1579(x[1579]), .x1580(x[1580]), .x1581(x[1581]), .x1582(x[1582]), .x1583(x[1583]), .x1584(x[1584]), .x1585(x[1585]), .x1586(x[1586]), .x1587(x[1587]), .x1588(x[1588]), .x1589(x[1589]), .x1590(x[1590]), .x1591(x[1591]), .x1592(x[1592]), .x1593(x[1593]), .x1594(x[1594]), .x1595(x[1595]), .x1596(x[1596]), .x1597(x[1597]), .x1598(x[1598]), .x1599(x[1599]), .x1600(x[1600]), .x1601(x[1601]), .x1602(x[1602]), .x1603(x[1603]), .x1604(x[1604]), .x1605(x[1605]), .x1606(x[1606]), .x1607(x[1607]), .x1608(x[1608]), .x1609(x[1609]), .x1610(x[1610]), .x1611(x[1611]), .x1612(x[1612]), .x1613(x[1613]), .x1614(x[1614]), .x1615(x[1615]), .x1616(x[1616]), .x1617(x[1617]), .x1618(x[1618]), .x1619(x[1619]), .x1620(x[1620]), .x1621(x[1621]), .x1622(x[1622]), .x1623(x[1623]), .x1624(x[1624]), .x1625(x[1625]), .x1626(x[1626]), .x1627(x[1627]), .x1628(x[1628]), .x1629(x[1629]), .x1630(x[1630]), .x1631(x[1631]), .x1632(x[1632]), .x1633(x[1633]), .x1634(x[1634]), .x1635(x[1635]), .x1636(x[1636]), .x1637(x[1637]), .x1638(x[1638]), .x1639(x[1639]), .x1640(x[1640]), .x1641(x[1641]), .x1642(x[1642]), .x1643(x[1643]), .x1644(x[1644]), .x1645(x[1645]), .x1646(x[1646]), .x1647(x[1647]), .x1648(x[1648]), .x1649(x[1649]), .x1650(x[1650]), .x1651(x[1651]), .x1652(x[1652]), .x1653(x[1653]), .x1654(x[1654]), .x1655(x[1655]), .x1656(x[1656]), .x1657(x[1657]), .x1658(x[1658]), .x1659(x[1659]), .x1660(x[1660]), .x1661(x[1661]), .x1662(x[1662]), .x1663(x[1663]), .x1664(x[1664]), .x1665(x[1665]), .x1666(x[1666]), .x1667(x[1667]), .x1668(x[1668]), .x1669(x[1669]), .x1670(x[1670]), .x1671(x[1671]), .x1672(x[1672]), .x1673(x[1673]), .x1674(x[1674]), .x1675(x[1675]), .x1676(x[1676]), .x1677(x[1677]), .x1678(x[1678]), .x1679(x[1679]), .x1680(x[1680]), .x1681(x[1681]), .x1682(x[1682]), .x1683(x[1683]), .x1684(x[1684]), .x1685(x[1685]), .x1686(x[1686]), .x1687(x[1687]), .x1688(x[1688]), .x1689(x[1689]), .x1690(x[1690]), .x1691(x[1691]), .x1692(x[1692]), .x1693(x[1693]), .x1694(x[1694]), .x1695(x[1695]), .x1696(x[1696]), .x1697(x[1697]), .x1698(x[1698]), .x1699(x[1699]), .x1700(x[1700]), .x1701(x[1701]), .x1702(x[1702]), .x1703(x[1703]), .x1704(x[1704]), .x1705(x[1705]), .x1706(x[1706]), .x1707(x[1707]), .x1708(x[1708]), .x1709(x[1709]), .x1710(x[1710]), .x1711(x[1711]), .x1712(x[1712]), .x1713(x[1713]), .x1714(x[1714]), .x1715(x[1715]), .x1716(x[1716]), .x1717(x[1717]), .x1718(x[1718]), .x1719(x[1719]), .x1720(x[1720]), .x1721(x[1721]), .x1722(x[1722]), .x1723(x[1723]), .x1724(x[1724]), .x1725(x[1725]), .x1726(x[1726]), .x1727(x[1727]), .x1728(x[1728]), .x1729(x[1729]), .x1730(x[1730]), .x1731(x[1731]), .x1732(x[1732]), .x1733(x[1733]), .x1734(x[1734]), .x1735(x[1735]), .x1736(x[1736]), .x1737(x[1737]), .x1738(x[1738]), .x1739(x[1739]), .x1740(x[1740]), .x1741(x[1741]), .x1742(x[1742]), .x1743(x[1743]), .x1744(x[1744]), .x1745(x[1745]), .x1746(x[1746]), .x1747(x[1747]), .x1748(x[1748]), .x1749(x[1749]), .x1750(x[1750]), .x1751(x[1751]), .x1752(x[1752]), .x1753(x[1753]), .x1754(x[1754]), .x1755(x[1755]), .x1756(x[1756]), .x1757(x[1757]), .x1758(x[1758]), .x1759(x[1759]), .x1760(x[1760]), .x1761(x[1761]), .x1762(x[1762]), .x1763(x[1763]), .x1764(x[1764]), .x1765(x[1765]), .x1766(x[1766]), .x1767(x[1767]), .x1768(x[1768]), .x1769(x[1769]), .x1770(x[1770]), .x1771(x[1771]), .x1772(x[1772]), .x1773(x[1773]), .x1774(x[1774]), .x1775(x[1775]), .x1776(x[1776]), .x1777(x[1777]), .x1778(x[1778]), .x1779(x[1779]), .x1780(x[1780]), .x1781(x[1781]), .x1782(x[1782]), .x1783(x[1783]), .x1784(x[1784]), .x1785(x[1785]), .x1786(x[1786]), .x1787(x[1787]), .x1788(x[1788]), .x1789(x[1789]), .x1790(x[1790]), .x1791(x[1791]), .x1792(x[1792]), .x1793(x[1793]), .x1794(x[1794]), .x1795(x[1795]), .x1796(x[1796]), .x1797(x[1797]), .x1798(x[1798]), .x1799(x[1799]), .x1800(x[1800]), .x1801(x[1801]), .x1802(x[1802]), .x1803(x[1803]), .x1804(x[1804]), .x1805(x[1805]), .x1806(x[1806]), .x1807(x[1807]), .x1808(x[1808]), .x1809(x[1809]), .x1810(x[1810]), .x1811(x[1811]), .x1812(x[1812]), .x1813(x[1813]), .x1814(x[1814]), .x1815(x[1815]), .x1816(x[1816]), .x1817(x[1817]), .x1818(x[1818]), .x1819(x[1819]), .x1820(x[1820]), .x1821(x[1821]), .x1822(x[1822]), .x1823(x[1823]), .x1824(x[1824]), .x1825(x[1825]), .x1826(x[1826]), .x1827(x[1827]), .x1828(x[1828]), .x1829(x[1829]), .x1830(x[1830]), .x1831(x[1831]), .x1832(x[1832]), .x1833(x[1833]), .x1834(x[1834]), .x1835(x[1835]), .x1836(x[1836]), .x1837(x[1837]), .x1838(x[1838]), .x1839(x[1839]), .x1840(x[1840]), .x1841(x[1841]), .x1842(x[1842]), .x1843(x[1843]), .x1844(x[1844]), .x1845(x[1845]), .x1846(x[1846]), .x1847(x[1847]), .x1848(x[1848]), .x1849(x[1849]), .x1850(x[1850]), .x1851(x[1851]), .x1852(x[1852]), .x1853(x[1853]), .x1854(x[1854]), .x1855(x[1855]), .x1856(x[1856]), .x1857(x[1857]), .x1858(x[1858]), .x1859(x[1859]), .x1860(x[1860]), .x1861(x[1861]), .x1862(x[1862]), .x1863(x[1863]), .x1864(x[1864]), .x1865(x[1865]), .x1866(x[1866]), .x1867(x[1867]), .x1868(x[1868]), .x1869(x[1869]), .x1870(x[1870]), .x1871(x[1871]), .x1872(x[1872]), .x1873(x[1873]), .x1874(x[1874]), .x1875(x[1875]), .x1876(x[1876]), .x1877(x[1877]), .x1878(x[1878]), .x1879(x[1879]), .x1880(x[1880]), .x1881(x[1881]), .x1882(x[1882]), .x1883(x[1883]), .x1884(x[1884]), .x1885(x[1885]), .x1886(x[1886]), .x1887(x[1887]), .x1888(x[1888]), .x1889(x[1889]), .x1890(x[1890]), .x1891(x[1891]), .x1892(x[1892]), .x1893(x[1893]), .x1894(x[1894]), .x1895(x[1895]), .x1896(x[1896]), .x1897(x[1897]), .x1898(x[1898]), .x1899(x[1899]), .x1900(x[1900]), .x1901(x[1901]), .x1902(x[1902]), .x1903(x[1903]), .x1904(x[1904]), .x1905(x[1905]), .x1906(x[1906]), .x1907(x[1907]), .x1908(x[1908]), .x1909(x[1909]), .x1910(x[1910]), .x1911(x[1911]), .x1912(x[1912]), .x1913(x[1913]), .x1914(x[1914]), .x1915(x[1915]), .x1916(x[1916]), .x1917(x[1917]), .x1918(x[1918]), .x1919(x[1919]), .x1920(x[1920]), .x1921(x[1921]), .x1922(x[1922]), .x1923(x[1923]), .x1924(x[1924]), .x1925(x[1925]), .x1926(x[1926]), .x1927(x[1927]), .x1928(x[1928]), .x1929(x[1929]), .x1930(x[1930]), .x1931(x[1931]), .x1932(x[1932]), .x1933(x[1933]), .x1934(x[1934]), .x1935(x[1935]), .x1936(x[1936]), .x1937(x[1937]), .x1938(x[1938]), .x1939(x[1939]), .x1940(x[1940]), .x1941(x[1941]), .x1942(x[1942]), .x1943(x[1943]), .x1944(x[1944]), .x1945(x[1945]), .x1946(x[1946]), .x1947(x[1947]), .x1948(x[1948]), .x1949(x[1949]), .x1950(x[1950]), .x1951(x[1951]), .x1952(x[1952]), .x1953(x[1953]), .x1954(x[1954]), .x1955(x[1955]), .x1956(x[1956]), .x1957(x[1957]), .x1958(x[1958]), .x1959(x[1959]), .x1960(x[1960]), .x1961(x[1961]), .x1962(x[1962]), .x1963(x[1963]), .x1964(x[1964]), .x1965(x[1965]), .x1966(x[1966]), .x1967(x[1967]), .x1968(x[1968]), .x1969(x[1969]), .x1970(x[1970]), .x1971(x[1971]), .x1972(x[1972]), .x1973(x[1973]), .x1974(x[1974]), .x1975(x[1975]), .x1976(x[1976]), .x1977(x[1977]), .x1978(x[1978]), .x1979(x[1979]), .x1980(x[1980]), .x1981(x[1981]), .x1982(x[1982]), .x1983(x[1983]), .x1984(x[1984]), .x1985(x[1985]), .x1986(x[1986]), .x1987(x[1987]), .x1988(x[1988]), .x1989(x[1989]), .x1990(x[1990]), .x1991(x[1991]), .x1992(x[1992]), .x1993(x[1993]), .x1994(x[1994]), .x1995(x[1995]), .x1996(x[1996]), .x1997(x[1997]), .x1998(x[1998]), .x1999(x[1999]), .x2000(x[2000]), .x2001(x[2001]), .x2002(x[2002]), .x2003(x[2003]), .x2004(x[2004]), .x2005(x[2005]), .x2006(x[2006]), .x2007(x[2007]), .x2008(x[2008]), .x2009(x[2009]), .x2010(x[2010]), .x2011(x[2011]), .x2012(x[2012]), .x2013(x[2013]), .x2014(x[2014]), .x2015(x[2015]), .x2016(x[2016]), .x2017(x[2017]), .x2018(x[2018]), .x2019(x[2019]), .x2020(x[2020]), .x2021(x[2021]), .x2022(x[2022]), .x2023(x[2023]), .x2024(x[2024]), .x2025(x[2025]), .x2026(x[2026]), .x2027(x[2027]), .x2028(x[2028]), .x2029(x[2029]), .x2030(x[2030]), .x2031(x[2031]), .x2032(x[2032]), .x2033(x[2033]), .x2034(x[2034]), .x2035(x[2035]), .x2036(x[2036]), .x2037(x[2037]), .x2038(x[2038]), .x2039(x[2039]), .x2040(x[2040]), .x2041(x[2041]), .x2042(x[2042]), .x2043(x[2043]), .x2044(x[2044]), .x2045(x[2045]), .x2046(x[2046]), .x2047(x[2047]), .x2048(x[2048]), .x2049(x[2049]), .x2050(x[2050]), .x2051(x[2051]), .x2052(x[2052]), .x2053(x[2053]), .x2054(x[2054]), .x2055(x[2055]), .x2056(x[2056]), .x2057(x[2057]), .x2058(x[2058]), .x2059(x[2059]), .x2060(x[2060]), .x2061(x[2061]), .x2062(x[2062]), .x2063(x[2063]), .x2064(x[2064]), .x2065(x[2065]), .x2066(x[2066]), .x2067(x[2067]), .x2068(x[2068]), .x2069(x[2069]), .x2070(x[2070]), .x2071(x[2071]), .x2072(x[2072]), .x2073(x[2073]), .x2074(x[2074]), .x2075(x[2075]), .x2076(x[2076]), .x2077(x[2077]), .x2078(x[2078]), .x2079(x[2079]), .x2080(x[2080]), .x2081(x[2081]), .x2082(x[2082]), .x2083(x[2083]), .x2084(x[2084]), .x2085(x[2085]), .x2086(x[2086]), .x2087(x[2087]), .x2088(x[2088]), .x2089(x[2089]), .x2090(x[2090]), .x2091(x[2091]), .x2092(x[2092]), .x2093(x[2093]), .x2094(x[2094]), .x2095(x[2095]), .x2096(x[2096]), .x2097(x[2097]), .x2098(x[2098]), .x2099(x[2099]), .x2100(x[2100]), .x2101(x[2101]), .x2102(x[2102]), .x2103(x[2103]), .x2104(x[2104]), .x2105(x[2105]), .x2106(x[2106]), .x2107(x[2107]), .x2108(x[2108]), .x2109(x[2109]), .x2110(x[2110]), .x2111(x[2111]), .x2112(x[2112]), .x2113(x[2113]), .x2114(x[2114]), .x2115(x[2115]), .x2116(x[2116]), .x2117(x[2117]), .x2118(x[2118]), .x2119(x[2119]), .x2120(x[2120]), .x2121(x[2121]), .x2122(x[2122]), .x2123(x[2123]), .x2124(x[2124]), .x2125(x[2125]), .x2126(x[2126]), .x2127(x[2127]), .x2128(x[2128]), .x2129(x[2129]), .x2130(x[2130]), .x2131(x[2131]), .x2132(x[2132]), .x2133(x[2133]), .x2134(x[2134]), .x2135(x[2135]), .x2136(x[2136]), .x2137(x[2137]), .x2138(x[2138]), .x2139(x[2139]), .x2140(x[2140]), .x2141(x[2141]), .x2142(x[2142]), .x2143(x[2143]), .x2144(x[2144]), .x2145(x[2145]), .x2146(x[2146]), .x2147(x[2147]), .x2148(x[2148]), .x2149(x[2149]), .x2150(x[2150]), .x2151(x[2151]), .x2152(x[2152]), .x2153(x[2153]), .x2154(x[2154]), .x2155(x[2155]), .x2156(x[2156]), .x2157(x[2157]), .x2158(x[2158]), .x2159(x[2159]), .x2160(x[2160]), .x2161(x[2161]), .x2162(x[2162]), .x2163(x[2163]), .x2164(x[2164]), .x2165(x[2165]), .x2166(x[2166]), .x2167(x[2167]), .x2168(x[2168]), .x2169(x[2169]), .x2170(x[2170]), .x2171(x[2171]), .x2172(x[2172]), .x2173(x[2173]), .x2174(x[2174]), .x2175(x[2175]), .x2176(x[2176]), .x2177(x[2177]), .x2178(x[2178]), .x2179(x[2179]), .x2180(x[2180]), .x2181(x[2181]), .x2182(x[2182]), .x2183(x[2183]), .x2184(x[2184]), .x2185(x[2185]), .x2186(x[2186]), .x2187(x[2187]), .x2188(x[2188]), .x2189(x[2189]), .x2190(x[2190]), .x2191(x[2191]), .x2192(x[2192]), .x2193(x[2193]), .x2194(x[2194]), .x2195(x[2195]), .x2196(x[2196]), .x2197(x[2197]), .x2198(x[2198]), .x2199(x[2199]), .x2200(x[2200]), .x2201(x[2201]), .x2202(x[2202]), .x2203(x[2203]), .x2204(x[2204]), .x2205(x[2205]), .x2206(x[2206]), .x2207(x[2207]), .x2208(x[2208]), .x2209(x[2209]), .x2210(x[2210]), .x2211(x[2211]), .x2212(x[2212]), .x2213(x[2213]), .x2214(x[2214]), .x2215(x[2215]), .x2216(x[2216]), .x2217(x[2217]), .x2218(x[2218]), .x2219(x[2219]), .x2220(x[2220]), .x2221(x[2221]), .x2222(x[2222]), .x2223(x[2223]), .x2224(x[2224]), .x2225(x[2225]), .x2226(x[2226]), .x2227(x[2227]), .x2228(x[2228]), .x2229(x[2229]), .x2230(x[2230]), .x2231(x[2231]), .x2232(x[2232]), .x2233(x[2233]), .x2234(x[2234]), .x2235(x[2235]), .x2236(x[2236]), .x2237(x[2237]), .x2238(x[2238]), .x2239(x[2239]), .x2240(x[2240]), .x2241(x[2241]), .x2242(x[2242]), .x2243(x[2243]), .x2244(x[2244]), .x2245(x[2245]), .x2246(x[2246]), .x2247(x[2247]), .x2248(x[2248]), .x2249(x[2249]), .x2250(x[2250]), .x2251(x[2251]), .x2252(x[2252]), .x2253(x[2253]), .x2254(x[2254]), .x2255(x[2255]), .x2256(x[2256]), .x2257(x[2257]), .x2258(x[2258]), .x2259(x[2259]), .x2260(x[2260]), .x2261(x[2261]), .x2262(x[2262]), .x2263(x[2263]), .x2264(x[2264]), .x2265(x[2265]), .x2266(x[2266]), .x2267(x[2267]), .x2268(x[2268]), .x2269(x[2269]), .x2270(x[2270]), .x2271(x[2271]), .x2272(x[2272]), .x2273(x[2273]), .x2274(x[2274]), .x2275(x[2275]), .x2276(x[2276]), .x2277(x[2277]), .x2278(x[2278]), .x2279(x[2279]), .x2280(x[2280]), .x2281(x[2281]), .x2282(x[2282]), .x2283(x[2283]), .x2284(x[2284]), .x2285(x[2285]), .x2286(x[2286]), .x2287(x[2287]), .x2288(x[2288]), .x2289(x[2289]), .x2290(x[2290]), .x2291(x[2291]), .x2292(x[2292]), .x2293(x[2293]), .x2294(x[2294]), .x2295(x[2295]), .x2296(x[2296]), .x2297(x[2297]), .x2298(x[2298]), .x2299(x[2299]), .x2300(x[2300]), .x2301(x[2301]), .x2302(x[2302]), .x2303(x[2303]), .x2304(x[2304]), .x2305(x[2305]), .x2306(x[2306]), .x2307(x[2307]), .x2308(x[2308]), .x2309(x[2309]), .x2310(x[2310]), .x2311(x[2311]), .x2312(x[2312]), .x2313(x[2313]), .x2314(x[2314]), .x2315(x[2315]), .x2316(x[2316]), .x2317(x[2317]), .x2318(x[2318]), .x2319(x[2319]), .x2320(x[2320]), .x2321(x[2321]), .x2322(x[2322]), .x2323(x[2323]), .x2324(x[2324]), .x2325(x[2325]), .x2326(x[2326]), .x2327(x[2327]), .x2328(x[2328]), .x2329(x[2329]), .x2330(x[2330]), .x2331(x[2331]), .x2332(x[2332]), .x2333(x[2333]), .x2334(x[2334]), .x2335(x[2335]), .x2336(x[2336]), .x2337(x[2337]), .x2338(x[2338]), .x2339(x[2339]), .x2340(x[2340]), .x2341(x[2341]), .x2342(x[2342]), .x2343(x[2343]), .x2344(x[2344]), .x2345(x[2345]), .x2346(x[2346]), .x2347(x[2347]), .x2348(x[2348]), .x2349(x[2349]), .x2350(x[2350]), .x2351(x[2351]), .x2352(x[2352]), .x2353(x[2353]), .x2354(x[2354]), .x2355(x[2355]), .x2356(x[2356]), .x2357(x[2357]), .x2358(x[2358]), .x2359(x[2359]), .x2360(x[2360]), .x2361(x[2361]), .x2362(x[2362]), .x2363(x[2363]), .x2364(x[2364]), .x2365(x[2365]), .x2366(x[2366]), .x2367(x[2367]), .x2368(x[2368]), .x2369(x[2369]), .x2370(x[2370]), .x2371(x[2371]), .x2372(x[2372]), .x2373(x[2373]), .x2374(x[2374]), .x2375(x[2375]), .x2376(x[2376]), .x2377(x[2377]), .x2378(x[2378]), .x2379(x[2379]), .x2380(x[2380]), .x2381(x[2381]), .x2382(x[2382]), .x2383(x[2383]), .x2384(x[2384]), .x2385(x[2385]), .x2386(x[2386]), .x2387(x[2387]), .x2388(x[2388]), .x2389(x[2389]), .x2390(x[2390]), .x2391(x[2391]), .x2392(x[2392]), .x2393(x[2393]), .x2394(x[2394]), .x2395(x[2395]), .x2396(x[2396]), .x2397(x[2397]), .x2398(x[2398]), .x2399(x[2399]), .x2400(x[2400]), .x2401(x[2401]), .x2402(x[2402]), .x2403(x[2403]), .x2404(x[2404]), .x2405(x[2405]), .x2406(x[2406]), .x2407(x[2407]), .x2408(x[2408]), .x2409(x[2409]), .x2410(x[2410]), .x2411(x[2411]), .x2412(x[2412]), .x2413(x[2413]), .x2414(x[2414]), .x2415(x[2415]), .x2416(x[2416]), .x2417(x[2417]), .x2418(x[2418]), .x2419(x[2419]), .x2420(x[2420]), .x2421(x[2421]), .x2422(x[2422]), .x2423(x[2423]), .x2424(x[2424]), .x2425(x[2425]), .x2426(x[2426]), .x2427(x[2427]), .x2428(x[2428]), .x2429(x[2429]), .x2430(x[2430]), .x2431(x[2431]), .x2432(x[2432]), .x2433(x[2433]), .x2434(x[2434]), .x2435(x[2435]), .x2436(x[2436]), .x2437(x[2437]), .x2438(x[2438]), .x2439(x[2439]), .x2440(x[2440]), .x2441(x[2441]), .x2442(x[2442]), .x2443(x[2443]), .x2444(x[2444]), .x2445(x[2445]), .x2446(x[2446]), .x2447(x[2447]), .x2448(x[2448]), .x2449(x[2449]), .x2450(x[2450]), .x2451(x[2451]), .x2452(x[2452]), .x2453(x[2453]), .x2454(x[2454]), .x2455(x[2455]), .x2456(x[2456]), .x2457(x[2457]), .x2458(x[2458]), .x2459(x[2459]), .x2460(x[2460]), .x2461(x[2461]), .x2462(x[2462]), .x2463(x[2463]), .x2464(x[2464]), .x2465(x[2465]), .x2466(x[2466]), .x2467(x[2467]), .x2468(x[2468]), .x2469(x[2469]), .x2470(x[2470]), .x2471(x[2471]), .x2472(x[2472]), .x2473(x[2473]), .x2474(x[2474]), .x2475(x[2475]), .x2476(x[2476]), .x2477(x[2477]), .x2478(x[2478]), .x2479(x[2479]), .x2480(x[2480]), .x2481(x[2481]), .x2482(x[2482]), .x2483(x[2483]), .x2484(x[2484]), .x2485(x[2485]), .x2486(x[2486]), .x2487(x[2487]), .x2488(x[2488]), .x2489(x[2489]), .x2490(x[2490]), .x2491(x[2491]), .x2492(x[2492]), .x2493(x[2493]), .x2494(x[2494]), .x2495(x[2495]), .x2496(x[2496]), .x2497(x[2497]), .x2498(x[2498]), .x2499(x[2499]), .x2500(x[2500]), .x2501(x[2501]), .x2502(x[2502]), .x2503(x[2503]), .x2504(x[2504]), .x2505(x[2505]), .x2506(x[2506]), .x2507(x[2507]), .x2508(x[2508]), .x2509(x[2509]), .x2510(x[2510]), .x2511(x[2511]), .x2512(x[2512]), .x2513(x[2513]), .x2514(x[2514]), .x2515(x[2515]), .x2516(x[2516]), .x2517(x[2517]), .x2518(x[2518]), .x2519(x[2519]), .x2520(x[2520]), .x2521(x[2521]), .x2522(x[2522]), .x2523(x[2523]), .x2524(x[2524]), .x2525(x[2525]), .x2526(x[2526]), .x2527(x[2527]), .x2528(x[2528]), .x2529(x[2529]), .x2530(x[2530]), .x2531(x[2531]), .x2532(x[2532]), .x2533(x[2533]), .x2534(x[2534]), .x2535(x[2535]), .x2536(x[2536]), .x2537(x[2537]), .x2538(x[2538]), .x2539(x[2539]), .x2540(x[2540]), .x2541(x[2541]), .x2542(x[2542]), .x2543(x[2543]), .x2544(x[2544]), .x2545(x[2545]), .x2546(x[2546]), .x2547(x[2547]), .x2548(x[2548]), .x2549(x[2549]), .x2550(x[2550]), .x2551(x[2551]), .x2552(x[2552]), .x2553(x[2553]), .x2554(x[2554]), .x2555(x[2555]), .x2556(x[2556]), .x2557(x[2557]), .x2558(x[2558]), .x2559(x[2559]), .x2560(x[2560]), .x2561(x[2561]), .x2562(x[2562]), .x2563(x[2563]), .x2564(x[2564]), .x2565(x[2565]), .x2566(x[2566]), .x2567(x[2567]), .x2568(x[2568]), .x2569(x[2569]), .x2570(x[2570]), .x2571(x[2571]), .x2572(x[2572]), .x2573(x[2573]), .x2574(x[2574]), .x2575(x[2575]), .x2576(x[2576]), .x2577(x[2577]), .x2578(x[2578]), .x2579(x[2579]), .x2580(x[2580]), .x2581(x[2581]), .x2582(x[2582]), .x2583(x[2583]), .x2584(x[2584]), .x2585(x[2585]), .x2586(x[2586]), .x2587(x[2587]), .x2588(x[2588]), .x2589(x[2589]), .x2590(x[2590]), .x2591(x[2591]), .x2592(x[2592]), .x2593(x[2593]), .x2594(x[2594]), .x2595(x[2595]), .x2596(x[2596]), .x2597(x[2597]), .x2598(x[2598]), .x2599(x[2599]), .x2600(x[2600]), .x2601(x[2601]), .x2602(x[2602]), .x2603(x[2603]), .x2604(x[2604]), .x2605(x[2605]), .x2606(x[2606]), .x2607(x[2607]), .x2608(x[2608]), .x2609(x[2609]), .x2610(x[2610]), .x2611(x[2611]), .x2612(x[2612]), .x2613(x[2613]), .x2614(x[2614]), .x2615(x[2615]), .x2616(x[2616]), .x2617(x[2617]), .x2618(x[2618]), .x2619(x[2619]), .x2620(x[2620]), .x2621(x[2621]), .x2622(x[2622]), .x2623(x[2623]), .x2624(x[2624]), .x2625(x[2625]), .x2626(x[2626]), .x2627(x[2627]), .x2628(x[2628]), .x2629(x[2629]), .x2630(x[2630]), .x2631(x[2631]), .x2632(x[2632]), .x2633(x[2633]), .x2634(x[2634]), .x2635(x[2635]), .x2636(x[2636]), .x2637(x[2637]), .x2638(x[2638]), .x2639(x[2639]), .x2640(x[2640]), .x2641(x[2641]), .x2642(x[2642]), .x2643(x[2643]), .x2644(x[2644]), .x2645(x[2645]), .x2646(x[2646]), .x2647(x[2647]), .x2648(x[2648]), .x2649(x[2649]), .x2650(x[2650]), .x2651(x[2651]), .x2652(x[2652]), .x2653(x[2653]), .x2654(x[2654]), .x2655(x[2655]), .x2656(x[2656]), .x2657(x[2657]), .x2658(x[2658]), .x2659(x[2659]), .x2660(x[2660]), .x2661(x[2661]), .x2662(x[2662]), .x2663(x[2663]), .x2664(x[2664]), .x2665(x[2665]), .x2666(x[2666]), .x2667(x[2667]), .x2668(x[2668]), .x2669(x[2669]), .x2670(x[2670]), .x2671(x[2671]), .x2672(x[2672]), .x2673(x[2673]), .x2674(x[2674]), .x2675(x[2675]), .x2676(x[2676]), .x2677(x[2677]), .x2678(x[2678]), .x2679(x[2679]), .x2680(x[2680]), .x2681(x[2681]), .x2682(x[2682]), .x2683(x[2683]), .x2684(x[2684]), .x2685(x[2685]), .x2686(x[2686]), .x2687(x[2687]), .x2688(x[2688]), .x2689(x[2689]), .x2690(x[2690]), .x2691(x[2691]), .x2692(x[2692]), .x2693(x[2693]), .x2694(x[2694]), .x2695(x[2695]), .x2696(x[2696]), .x2697(x[2697]), .x2698(x[2698]), .x2699(x[2699]), .x2700(x[2700]), .x2701(x[2701]), .x2702(x[2702]), .x2703(x[2703]), .x2704(x[2704]), .x2705(x[2705]), .x2706(x[2706]), .x2707(x[2707]), .x2708(x[2708]), .x2709(x[2709]), .x2710(x[2710]), .x2711(x[2711]), .x2712(x[2712]), .x2713(x[2713]), .x2714(x[2714]), .x2715(x[2715]), .x2716(x[2716]), .x2717(x[2717]), .x2718(x[2718]), .x2719(x[2719]), .x2720(x[2720]), .x2721(x[2721]), .x2722(x[2722]), .x2723(x[2723]), .x2724(x[2724]), .x2725(x[2725]), .x2726(x[2726]), .x2727(x[2727]), .x2728(x[2728]), .x2729(x[2729]), .x2730(x[2730]), .x2731(x[2731]), .x2732(x[2732]), .x2733(x[2733]), .x2734(x[2734]), .x2735(x[2735]), .x2736(x[2736]), .x2737(x[2737]), .x2738(x[2738]), .x2739(x[2739]), .x2740(x[2740]), .x2741(x[2741]), .x2742(x[2742]), .x2743(x[2743]), .x2744(x[2744]), .x2745(x[2745]), .x2746(x[2746]), .x2747(x[2747]), .x2748(x[2748]), .x2749(x[2749]), .x2750(x[2750]), .x2751(x[2751]), .x2752(x[2752]), .x2753(x[2753]), .x2754(x[2754]), .x2755(x[2755]), .x2756(x[2756]), .x2757(x[2757]), .x2758(x[2758]), .x2759(x[2759]), .x2760(x[2760]), .x2761(x[2761]), .x2762(x[2762]), .x2763(x[2763]), .x2764(x[2764]), .x2765(x[2765]), .x2766(x[2766]), .x2767(x[2767]), .x2768(x[2768]), .x2769(x[2769]), .x2770(x[2770]), .x2771(x[2771]), .x2772(x[2772]), .x2773(x[2773]), .x2774(x[2774]), .x2775(x[2775]), .x2776(x[2776]), .x2777(x[2777]), .x2778(x[2778]), .x2779(x[2779]), .x2780(x[2780]), .x2781(x[2781]), .x2782(x[2782]), .x2783(x[2783]), .x2784(x[2784]), .x2785(x[2785]), .x2786(x[2786]), .x2787(x[2787]), .x2788(x[2788]), .x2789(x[2789]), .x2790(x[2790]), .x2791(x[2791]), .x2792(x[2792]), .x2793(x[2793]), .x2794(x[2794]), .x2795(x[2795]), .x2796(x[2796]), .x2797(x[2797]), .x2798(x[2798]), .x2799(x[2799]), .x2800(x[2800]), .x2801(x[2801]), .x2802(x[2802]), .x2803(x[2803]), .x2804(x[2804]), .x2805(x[2805]), .x2806(x[2806]), .x2807(x[2807]), .x2808(x[2808]), .x2809(x[2809]), .x2810(x[2810]), .x2811(x[2811]), .x2812(x[2812]), .x2813(x[2813]), .x2814(x[2814]), .x2815(x[2815]), .x2816(x[2816]), .x2817(x[2817]), .x2818(x[2818]), .x2819(x[2819]), .x2820(x[2820]), .x2821(x[2821]), .x2822(x[2822]), .x2823(x[2823]), .x2824(x[2824]), .x2825(x[2825]), .x2826(x[2826]), .x2827(x[2827]), .x2828(x[2828]), .x2829(x[2829]), .x2830(x[2830]), .x2831(x[2831]), .x2832(x[2832]), .x2833(x[2833]), .x2834(x[2834]), .x2835(x[2835]), .x2836(x[2836]), .x2837(x[2837]), .x2838(x[2838]), .x2839(x[2839]), .x2840(x[2840]), .x2841(x[2841]), .x2842(x[2842]), .x2843(x[2843]), .x2844(x[2844]), .x2845(x[2845]), .x2846(x[2846]), .x2847(x[2847]), .x2848(x[2848]), .x2849(x[2849]), .x2850(x[2850]), .x2851(x[2851]), .x2852(x[2852]), .x2853(x[2853]), .x2854(x[2854]), .x2855(x[2855]), .x2856(x[2856]), .x2857(x[2857]), .x2858(x[2858]), .x2859(x[2859]), .x2860(x[2860]), .x2861(x[2861]), .x2862(x[2862]), .x2863(x[2863]), .x2864(x[2864]), .x2865(x[2865]), .x2866(x[2866]), .x2867(x[2867]), .x2868(x[2868]), .x2869(x[2869]), .x2870(x[2870]), .x2871(x[2871]), .x2872(x[2872]), .x2873(x[2873]), .x2874(x[2874]), .x2875(x[2875]), .x2876(x[2876]), .x2877(x[2877]), .x2878(x[2878]), .x2879(x[2879]), .x2880(x[2880]), .x2881(x[2881]), .x2882(x[2882]), .x2883(x[2883]), .x2884(x[2884]), .x2885(x[2885]), .x2886(x[2886]), .x2887(x[2887]), .x2888(x[2888]), .x2889(x[2889]), .x2890(x[2890]), .x2891(x[2891]), .x2892(x[2892]), .x2893(x[2893]), .x2894(x[2894]), .x2895(x[2895]), .x2896(x[2896]), .x2897(x[2897]), .x2898(x[2898]), .x2899(x[2899]), .x2900(x[2900]), .x2901(x[2901]), .x2902(x[2902]), .x2903(x[2903]), .x2904(x[2904]), .x2905(x[2905]), .x2906(x[2906]), .x2907(x[2907]), .x2908(x[2908]), .x2909(x[2909]), .x2910(x[2910]), .x2911(x[2911]), .x2912(x[2912]), .x2913(x[2913]), .x2914(x[2914]), .x2915(x[2915]), .x2916(x[2916]), .x2917(x[2917]), .x2918(x[2918]), .x2919(x[2919]), .x2920(x[2920]), .x2921(x[2921]), .x2922(x[2922]), .x2923(x[2923]), .x2924(x[2924]), .x2925(x[2925]), .x2926(x[2926]), .x2927(x[2927]), .x2928(x[2928]), .x2929(x[2929]), .x2930(x[2930]), .x2931(x[2931]), .x2932(x[2932]), .x2933(x[2933]), .x2934(x[2934]), .x2935(x[2935]), .x2936(x[2936]), .x2937(x[2937]), .x2938(x[2938]), .x2939(x[2939]), .x2940(x[2940]), .x2941(x[2941]), .x2942(x[2942]), .x2943(x[2943]), .x2944(x[2944]), .x2945(x[2945]), .x2946(x[2946]), .x2947(x[2947]), .x2948(x[2948]), .x2949(x[2949]), .x2950(x[2950]), .x2951(x[2951]), .x2952(x[2952]), .x2953(x[2953]), .x2954(x[2954]), .x2955(x[2955]), .x2956(x[2956]), .x2957(x[2957]), .x2958(x[2958]), .x2959(x[2959]), .x2960(x[2960]), .x2961(x[2961]), .x2962(x[2962]), .x2963(x[2963]), .x2964(x[2964]), .x2965(x[2965]), .x2966(x[2966]), .x2967(x[2967]), .x2968(x[2968]), .x2969(x[2969]), .x2970(x[2970]), .x2971(x[2971]), .x2972(x[2972]), .x2973(x[2973]), .x2974(x[2974]), .x2975(x[2975]), .x2976(x[2976]), .x2977(x[2977]), .x2978(x[2978]), .x2979(x[2979]), .x2980(x[2980]), .x2981(x[2981]), .x2982(x[2982]), .x2983(x[2983]), .x2984(x[2984]), .x2985(x[2985]), .x2986(x[2986]), .x2987(x[2987]), .x2988(x[2988]), .x2989(x[2989]), .x2990(x[2990]), .x2991(x[2991]), .x2992(x[2992]), .x2993(x[2993]), .x2994(x[2994]), .x2995(x[2995]), .x2996(x[2996]), .x2997(x[2997]), .x2998(x[2998]), .x2999(x[2999]), .x3000(x[3000]), .x3001(x[3001]), .x3002(x[3002]), .x3003(x[3003]), .x3004(x[3004]), .x3005(x[3005]), .x3006(x[3006]), .x3007(x[3007]), .x3008(x[3008]), .x3009(x[3009]), .x3010(x[3010]), .x3011(x[3011]), .x3012(x[3012]), .x3013(x[3013]), .x3014(x[3014]), .x3015(x[3015]), .x3016(x[3016]), .x3017(x[3017]), .x3018(x[3018]), .x3019(x[3019]), .x3020(x[3020]), .x3021(x[3021]), .x3022(x[3022]), .x3023(x[3023]), .x3024(x[3024]), .x3025(x[3025]), .x3026(x[3026]), .x3027(x[3027]), .x3028(x[3028]), .x3029(x[3029]), .x3030(x[3030]), .x3031(x[3031]), .x3032(x[3032]), .x3033(x[3033]), .x3034(x[3034]), .x3035(x[3035]), .x3036(x[3036]), .x3037(x[3037]), .x3038(x[3038]), .x3039(x[3039]), .x3040(x[3040]), .x3041(x[3041]), .x3042(x[3042]), .x3043(x[3043]), .x3044(x[3044]), .x3045(x[3045]), .x3046(x[3046]), .x3047(x[3047]), .x3048(x[3048]), .x3049(x[3049]), .x3050(x[3050]), .x3051(x[3051]), .x3052(x[3052]), .x3053(x[3053]), .x3054(x[3054]), .x3055(x[3055]), .x3056(x[3056]), .x3057(x[3057]), .x3058(x[3058]), .x3059(x[3059]), .x3060(x[3060]), .x3061(x[3061]), .x3062(x[3062]), .x3063(x[3063]), .x3064(x[3064]), .x3065(x[3065]), .x3066(x[3066]), .x3067(x[3067]), .x3068(x[3068]), .x3069(x[3069]), .x3070(x[3070]), .x3071(x[3071]), .x3072(x[3072]), .x3073(x[3073]), .x3074(x[3074]), .x3075(x[3075]), .x3076(x[3076]), .x3077(x[3077]), .x3078(x[3078]), .x3079(x[3079]), .x3080(x[3080]), .x3081(x[3081]), .x3082(x[3082]), .x3083(x[3083]), .x3084(x[3084]), .x3085(x[3085]), .x3086(x[3086]), .x3087(x[3087]), .x3088(x[3088]), .x3089(x[3089]), .x3090(x[3090]), .x3091(x[3091]), .x3092(x[3092]), .x3093(x[3093]), .x3094(x[3094]), .x3095(x[3095]), .x3096(x[3096]), .x3097(x[3097]), .x3098(x[3098]), .x3099(x[3099]), .x3100(x[3100]), .x3101(x[3101]), .x3102(x[3102]), .x3103(x[3103]), .x3104(x[3104]), .x3105(x[3105]), .x3106(x[3106]), .x3107(x[3107]), .x3108(x[3108]), .x3109(x[3109]), .x3110(x[3110]), .x3111(x[3111]), .x3112(x[3112]), .x3113(x[3113]), .x3114(x[3114]), .x3115(x[3115]), .x3116(x[3116]), .x3117(x[3117]), .x3118(x[3118]), .x3119(x[3119]), .x3120(x[3120]), .x3121(x[3121]), .x3122(x[3122]), .x3123(x[3123]), .x3124(x[3124]), .x3125(x[3125]), .x3126(x[3126]), .x3127(x[3127]), .x3128(x[3128]), .x3129(x[3129]), .x3130(x[3130]), .x3131(x[3131]), .x3132(x[3132]), .x3133(x[3133]), .x3134(x[3134]), .x3135(x[3135]), .x3136(x[3136]), .x3137(x[3137]), .x3138(x[3138]), .x3139(x[3139]), .x3140(x[3140]), .x3141(x[3141]), .x3142(x[3142]), .x3143(x[3143]), .x3144(x[3144]), .x3145(x[3145]), .x3146(x[3146]), .x3147(x[3147]), .x3148(x[3148]), .x3149(x[3149]), .x3150(x[3150]), .x3151(x[3151]), .x3152(x[3152]), .x3153(x[3153]), .x3154(x[3154]), .x3155(x[3155]), .x3156(x[3156]), .x3157(x[3157]), .x3158(x[3158]), .x3159(x[3159]), .x3160(x[3160]), .x3161(x[3161]), .x3162(x[3162]), .x3163(x[3163]), .x3164(x[3164]), .x3165(x[3165]), .x3166(x[3166]), .x3167(x[3167]), .x3168(x[3168]), .x3169(x[3169]), .x3170(x[3170]), .x3171(x[3171]), .x3172(x[3172]), .x3173(x[3173]), .x3174(x[3174]), .x3175(x[3175]), .x3176(x[3176]), .x3177(x[3177]), .x3178(x[3178]), .x3179(x[3179]), .x3180(x[3180]), .x3181(x[3181]), .x3182(x[3182]), .x3183(x[3183]), .x3184(x[3184]), .x3185(x[3185]), .x3186(x[3186]), .x3187(x[3187]), .x3188(x[3188]), .x3189(x[3189]), .x3190(x[3190]), .x3191(x[3191]), .x3192(x[3192]), .x3193(x[3193]), .x3194(x[3194]), .x3195(x[3195]), .x3196(x[3196]), .x3197(x[3197]), .x3198(x[3198]), .x3199(x[3199]), .x3200(x[3200]), .x3201(x[3201]), .x3202(x[3202]), .x3203(x[3203]), .x3204(x[3204]), .x3205(x[3205]), .x3206(x[3206]), .x3207(x[3207]), .x3208(x[3208]), .x3209(x[3209]), .x3210(x[3210]), .x3211(x[3211]), .x3212(x[3212]), .x3213(x[3213]), .x3214(x[3214]), .x3215(x[3215]), .x3216(x[3216]), .x3217(x[3217]), .x3218(x[3218]), .x3219(x[3219]), .x3220(x[3220]), .x3221(x[3221]), .x3222(x[3222]), .x3223(x[3223]), .x3224(x[3224]), .x3225(x[3225]), .x3226(x[3226]), .x3227(x[3227]), .x3228(x[3228]), .x3229(x[3229]), .x3230(x[3230]), .x3231(x[3231]), .x3232(x[3232]), .x3233(x[3233]), .x3234(x[3234]), .x3235(x[3235]), .x3236(x[3236]), .x3237(x[3237]), .x3238(x[3238]), .x3239(x[3239]), .x3240(x[3240]), .x3241(x[3241]), .x3242(x[3242]), .x3243(x[3243]), .x3244(x[3244]), .x3245(x[3245]), .x3246(x[3246]), .x3247(x[3247]), .x3248(x[3248]), .x3249(x[3249]), .x3250(x[3250]), .x3251(x[3251]), .x3252(x[3252]), .x3253(x[3253]), .x3254(x[3254]), .x3255(x[3255]), .x3256(x[3256]), .x3257(x[3257]), .x3258(x[3258]), .x3259(x[3259]), .x3260(x[3260]), .x3261(x[3261]), .x3262(x[3262]), .x3263(x[3263]), .x3264(x[3264]), .x3265(x[3265]), .x3266(x[3266]), .x3267(x[3267]), .x3268(x[3268]), .x3269(x[3269]), .x3270(x[3270]), .x3271(x[3271]), .x3272(x[3272]), .x3273(x[3273]), .x3274(x[3274]), .x3275(x[3275]), .x3276(x[3276]), .x3277(x[3277]), .x3278(x[3278]), .x3279(x[3279]), .x3280(x[3280]), .x3281(x[3281]), .x3282(x[3282]), .x3283(x[3283]), .x3284(x[3284]), .x3285(x[3285]), .x3286(x[3286]), .x3287(x[3287]), .x3288(x[3288]), .x3289(x[3289]), .x3290(x[3290]), .x3291(x[3291]), .x3292(x[3292]), .x3293(x[3293]), .x3294(x[3294]), .x3295(x[3295]), .x3296(x[3296]), .x3297(x[3297]), .x3298(x[3298]), .x3299(x[3299]), .x3300(x[3300]), .x3301(x[3301]), .x3302(x[3302]), .x3303(x[3303]), .x3304(x[3304]), .x3305(x[3305]), .x3306(x[3306]), .x3307(x[3307]), .x3308(x[3308]), .x3309(x[3309]), .x3310(x[3310]), .x3311(x[3311]), .x3312(x[3312]), .x3313(x[3313]), .x3314(x[3314]), .x3315(x[3315]), .x3316(x[3316]), .x3317(x[3317]), .x3318(x[3318]), .x3319(x[3319]), .x3320(x[3320]), .x3321(x[3321]), .x3322(x[3322]), .x3323(x[3323]), .x3324(x[3324]), .x3325(x[3325]), .x3326(x[3326]), .x3327(x[3327]), .x3328(x[3328]), .x3329(x[3329]), .x3330(x[3330]), .x3331(x[3331]), .x3332(x[3332]), .x3333(x[3333]), .x3334(x[3334]), .x3335(x[3335]), .x3336(x[3336]), .x3337(x[3337]), .x3338(x[3338]), .x3339(x[3339]), .x3340(x[3340]), .x3341(x[3341]), .x3342(x[3342]), .x3343(x[3343]), .x3344(x[3344]), .x3345(x[3345]), .x3346(x[3346]), .x3347(x[3347]), .x3348(x[3348]), .x3349(x[3349]), .x3350(x[3350]), .x3351(x[3351]), .x3352(x[3352]), .x3353(x[3353]), .x3354(x[3354]), .x3355(x[3355]), .x3356(x[3356]), .x3357(x[3357]), .x3358(x[3358]), .x3359(x[3359]), .x3360(x[3360]), .x3361(x[3361]), .x3362(x[3362]), .x3363(x[3363]), .x3364(x[3364]), .x3365(x[3365]), .x3366(x[3366]), .x3367(x[3367]), .x3368(x[3368]), .x3369(x[3369]), .x3370(x[3370]), .x3371(x[3371]), .x3372(x[3372]), .x3373(x[3373]), .x3374(x[3374]), .x3375(x[3375]), .x3376(x[3376]), .x3377(x[3377]), .x3378(x[3378]), .x3379(x[3379]), .x3380(x[3380]), .x3381(x[3381]), .x3382(x[3382]), .x3383(x[3383]), .x3384(x[3384]), .x3385(x[3385]), .x3386(x[3386]), .x3387(x[3387]), .x3388(x[3388]), .x3389(x[3389]), .x3390(x[3390]), .x3391(x[3391]), .x3392(x[3392]), .x3393(x[3393]), .x3394(x[3394]), .x3395(x[3395]), .x3396(x[3396]), .x3397(x[3397]), .x3398(x[3398]), .x3399(x[3399]), .x3400(x[3400]), .x3401(x[3401]), .x3402(x[3402]), .x3403(x[3403]), .x3404(x[3404]), .x3405(x[3405]), .x3406(x[3406]), .x3407(x[3407]), .x3408(x[3408]), .x3409(x[3409]), .x3410(x[3410]), .x3411(x[3411]), .x3412(x[3412]), .x3413(x[3413]), .x3414(x[3414]), .x3415(x[3415]), .x3416(x[3416]), .x3417(x[3417]), .x3418(x[3418]), .x3419(x[3419]), .x3420(x[3420]), .x3421(x[3421]), .x3422(x[3422]), .x3423(x[3423]), .x3424(x[3424]), .x3425(x[3425]), .x3426(x[3426]), .x3427(x[3427]), .x3428(x[3428]), .x3429(x[3429]), .x3430(x[3430]), .x3431(x[3431]), .x3432(x[3432]), .x3433(x[3433]), .x3434(x[3434]), .x3435(x[3435]), .x3436(x[3436]), .x3437(x[3437]), .x3438(x[3438]), .x3439(x[3439]), .x3440(x[3440]), .x3441(x[3441]), .x3442(x[3442]), .x3443(x[3443]), .x3444(x[3444]), .x3445(x[3445]), .x3446(x[3446]), .x3447(x[3447]), .x3448(x[3448]), .x3449(x[3449]), .x3450(x[3450]), .x3451(x[3451]), .x3452(x[3452]), .x3453(x[3453]), .x3454(x[3454]), .x3455(x[3455]), .x3456(x[3456]), .x3457(x[3457]), .x3458(x[3458]), .x3459(x[3459]), .x3460(x[3460]), .x3461(x[3461]), .x3462(x[3462]), .x3463(x[3463]), .x3464(x[3464]), .x3465(x[3465]), .x3466(x[3466]), .x3467(x[3467]), .x3468(x[3468]), .x3469(x[3469]), .x3470(x[3470]), .x3471(x[3471]), .x3472(x[3472]), .x3473(x[3473]), .x3474(x[3474]), .x3475(x[3475]), .x3476(x[3476]), .x3477(x[3477]), .x3478(x[3478]), .x3479(x[3479]), .x3480(x[3480]), .x3481(x[3481]), .x3482(x[3482]), .x3483(x[3483]), .x3484(x[3484]), .x3485(x[3485]), .x3486(x[3486]), .x3487(x[3487]), .x3488(x[3488]), .x3489(x[3489]), .x3490(x[3490]), .x3491(x[3491]), .x3492(x[3492]), .x3493(x[3493]), .x3494(x[3494]), .x3495(x[3495]), .x3496(x[3496]), .x3497(x[3497]), .x3498(x[3498]), .x3499(x[3499]), .x3500(x[3500]), .x3501(x[3501]), .x3502(x[3502]), .x3503(x[3503]), .x3504(x[3504]), .x3505(x[3505]), .x3506(x[3506]), .x3507(x[3507]), .x3508(x[3508]), .x3509(x[3509]), .x3510(x[3510]), .x3511(x[3511]), .x3512(x[3512]), .x3513(x[3513]), .x3514(x[3514]), .x3515(x[3515]), .x3516(x[3516]), .x3517(x[3517]), .x3518(x[3518]), .x3519(x[3519]), .x3520(x[3520]), .x3521(x[3521]), .x3522(x[3522]), .x3523(x[3523]), .x3524(x[3524]), .x3525(x[3525]), .x3526(x[3526]), .x3527(x[3527]), .x3528(x[3528]), .x3529(x[3529]), .x3530(x[3530]), .x3531(x[3531]), .x3532(x[3532]), .x3533(x[3533]), .x3534(x[3534]), .x3535(x[3535]), .x3536(x[3536]), .x3537(x[3537]), .x3538(x[3538]), .x3539(x[3539]), .x3540(x[3540]), .x3541(x[3541]), .x3542(x[3542]), .x3543(x[3543]), .x3544(x[3544]), .x3545(x[3545]), .x3546(x[3546]), .x3547(x[3547]), .x3548(x[3548]), .x3549(x[3549]), .x3550(x[3550]), .x3551(x[3551]), .x3552(x[3552]), .x3553(x[3553]), .x3554(x[3554]), .x3555(x[3555]), .x3556(x[3556]), .x3557(x[3557]), .x3558(x[3558]), .x3559(x[3559]), .x3560(x[3560]), .x3561(x[3561]), .x3562(x[3562]), .x3563(x[3563]), .x3564(x[3564]), .x3565(x[3565]), .x3566(x[3566]), .x3567(x[3567]), .x3568(x[3568]), .x3569(x[3569]), .x3570(x[3570]), .x3571(x[3571]), .x3572(x[3572]), .x3573(x[3573]), .x3574(x[3574]), .x3575(x[3575]), .x3576(x[3576]), .x3577(x[3577]), .x3578(x[3578]), .x3579(x[3579]), .x3580(x[3580]), .x3581(x[3581]), .x3582(x[3582]), .x3583(x[3583]), .x3584(x[3584]), .x3585(x[3585]), .x3586(x[3586]), .x3587(x[3587]), .x3588(x[3588]), .x3589(x[3589]), .x3590(x[3590]), .x3591(x[3591]), .x3592(x[3592]), .x3593(x[3593]), .x3594(x[3594]), .x3595(x[3595]), .x3596(x[3596]), .x3597(x[3597]), .x3598(x[3598]), .x3599(x[3599]), .x3600(x[3600]), .x3601(x[3601]), .x3602(x[3602]), .x3603(x[3603]), .x3604(x[3604]), .x3605(x[3605]), .x3606(x[3606]), .x3607(x[3607]), .x3608(x[3608]), .x3609(x[3609]), .x3610(x[3610]), .x3611(x[3611]), .x3612(x[3612]), .x3613(x[3613]), .x3614(x[3614]), .x3615(x[3615]), .x3616(x[3616]), .x3617(x[3617]), .x3618(x[3618]), .x3619(x[3619]), .x3620(x[3620]), .x3621(x[3621]), .x3622(x[3622]), .x3623(x[3623]), .x3624(x[3624]), .x3625(x[3625]), .x3626(x[3626]), .x3627(x[3627]), .x3628(x[3628]), .x3629(x[3629]), .x3630(x[3630]), .x3631(x[3631]), .x3632(x[3632]), .x3633(x[3633]), .x3634(x[3634]), .x3635(x[3635]), .x3636(x[3636]), .x3637(x[3637]), .x3638(x[3638]), .x3639(x[3639]), .x3640(x[3640]), .x3641(x[3641]), .x3642(x[3642]), .x3643(x[3643]), .x3644(x[3644]), .x3645(x[3645]), .x3646(x[3646]), .x3647(x[3647]), .x3648(x[3648]), .x3649(x[3649]), .x3650(x[3650]), .x3651(x[3651]), .x3652(x[3652]), .x3653(x[3653]), .x3654(x[3654]), .x3655(x[3655]), .x3656(x[3656]), .x3657(x[3657]), .x3658(x[3658]), .x3659(x[3659]), .x3660(x[3660]), .x3661(x[3661]), .x3662(x[3662]), .x3663(x[3663]), .x3664(x[3664]), .x3665(x[3665]), .x3666(x[3666]), .x3667(x[3667]), .x3668(x[3668]), .x3669(x[3669]), .x3670(x[3670]), .x3671(x[3671]), .x3672(x[3672]), .x3673(x[3673]), .x3674(x[3674]), .x3675(x[3675]), .x3676(x[3676]), .x3677(x[3677]), .x3678(x[3678]), .x3679(x[3679]), .x3680(x[3680]), .x3681(x[3681]), .x3682(x[3682]), .x3683(x[3683]), .x3684(x[3684]), .x3685(x[3685]), .x3686(x[3686]), .x3687(x[3687]), .x3688(x[3688]), .x3689(x[3689]), .x3690(x[3690]), .x3691(x[3691]), .x3692(x[3692]), .x3693(x[3693]), .x3694(x[3694]), .x3695(x[3695]), .x3696(x[3696]), .x3697(x[3697]), .x3698(x[3698]), .x3699(x[3699]), .x3700(x[3700]), .x3701(x[3701]), .x3702(x[3702]), .x3703(x[3703]), .x3704(x[3704]), .x3705(x[3705]), .x3706(x[3706]), .x3707(x[3707]), .x3708(x[3708]), .x3709(x[3709]), .x3710(x[3710]), .x3711(x[3711]), .x3712(x[3712]), .x3713(x[3713]), .x3714(x[3714]), .x3715(x[3715]), .x3716(x[3716]), .x3717(x[3717]), .x3718(x[3718]), .x3719(x[3719]), .x3720(x[3720]), .x3721(x[3721]), .x3722(x[3722]), .x3723(x[3723]), .x3724(x[3724]), .x3725(x[3725]), .x3726(x[3726]), .x3727(x[3727]), .x3728(x[3728]), .x3729(x[3729]), .x3730(x[3730]), .x3731(x[3731]), .x3732(x[3732]), .x3733(x[3733]), .x3734(x[3734]), .x3735(x[3735]), .x3736(x[3736]), .x3737(x[3737]), .x3738(x[3738]), .x3739(x[3739]), .x3740(x[3740]), .x3741(x[3741]), .x3742(x[3742]), .x3743(x[3743]), .x3744(x[3744]), .x3745(x[3745]), .x3746(x[3746]), .x3747(x[3747]), .x3748(x[3748]), .x3749(x[3749]), .x3750(x[3750]), .x3751(x[3751]), .x3752(x[3752]), .x3753(x[3753]), .x3754(x[3754]), .x3755(x[3755]), .x3756(x[3756]), .x3757(x[3757]), .x3758(x[3758]), .x3759(x[3759]), .x3760(x[3760]), .x3761(x[3761]), .x3762(x[3762]), .x3763(x[3763]), .x3764(x[3764]), .x3765(x[3765]), .x3766(x[3766]), .x3767(x[3767]), .x3768(x[3768]), .x3769(x[3769]), .x3770(x[3770]), .x3771(x[3771]), .x3772(x[3772]), .x3773(x[3773]), .x3774(x[3774]), .x3775(x[3775]), .x3776(x[3776]), .x3777(x[3777]), .x3778(x[3778]), .x3779(x[3779]), .x3780(x[3780]), .x3781(x[3781]), .x3782(x[3782]), .x3783(x[3783]), .x3784(x[3784]), .x3785(x[3785]), .x3786(x[3786]), .x3787(x[3787]), .x3788(x[3788]), .x3789(x[3789]), .x3790(x[3790]), .x3791(x[3791]), .x3792(x[3792]), .x3793(x[3793]), .x3794(x[3794]), .x3795(x[3795]), .x3796(x[3796]), .x3797(x[3797]), .x3798(x[3798]), .x3799(x[3799]), .x3800(x[3800]), .x3801(x[3801]), .x3802(x[3802]), .x3803(x[3803]), .x3804(x[3804]), .x3805(x[3805]), .x3806(x[3806]), .x3807(x[3807]), .x3808(x[3808]), .x3809(x[3809]), .x3810(x[3810]), .x3811(x[3811]), .x3812(x[3812]), .x3813(x[3813]), .x3814(x[3814]), .x3815(x[3815]), .x3816(x[3816]), .x3817(x[3817]), .x3818(x[3818]), .x3819(x[3819]), .x3820(x[3820]), .x3821(x[3821]), .x3822(x[3822]), .x3823(x[3823]), .x3824(x[3824]), .x3825(x[3825]), .x3826(x[3826]), .x3827(x[3827]), .x3828(x[3828]), .x3829(x[3829]), .x3830(x[3830]), .x3831(x[3831]), .x3832(x[3832]), .x3833(x[3833]), .x3834(x[3834]), .x3835(x[3835]), .x3836(x[3836]), .x3837(x[3837]), .x3838(x[3838]), .x3839(x[3839]), .x3840(x[3840]), .x3841(x[3841]), .x3842(x[3842]), .x3843(x[3843]), .x3844(x[3844]), .x3845(x[3845]), .x3846(x[3846]), .x3847(x[3847]), .x3848(x[3848]), .x3849(x[3849]), .x3850(x[3850]), .x3851(x[3851]), .x3852(x[3852]), .x3853(x[3853]), .x3854(x[3854]), .x3855(x[3855]), .x3856(x[3856]), .x3857(x[3857]), .x3858(x[3858]), .x3859(x[3859]), .x3860(x[3860]), .x3861(x[3861]), .x3862(x[3862]), .x3863(x[3863]), .x3864(x[3864]), .x3865(x[3865]), .x3866(x[3866]), .x3867(x[3867]), .x3868(x[3868]), .x3869(x[3869]), .x3870(x[3870]), .x3871(x[3871]), .x3872(x[3872]), .x3873(x[3873]), .x3874(x[3874]), .x3875(x[3875]), .x3876(x[3876]), .x3877(x[3877]), .x3878(x[3878]), .x3879(x[3879]), .x3880(x[3880]), .x3881(x[3881]), .x3882(x[3882]), .x3883(x[3883]), .x3884(x[3884]), .x3885(x[3885]), .x3886(x[3886]), .x3887(x[3887]), .x3888(x[3888]), .x3889(x[3889]), .x3890(x[3890]), .x3891(x[3891]), .x3892(x[3892]), .x3893(x[3893]), .x3894(x[3894]), .x3895(x[3895]), .x3896(x[3896]), .x3897(x[3897]), .x3898(x[3898]), .x3899(x[3899]), .x3900(x[3900]), .x3901(x[3901]), .x3902(x[3902]), .x3903(x[3903]), .x3904(x[3904]), .x3905(x[3905]), .x3906(x[3906]), .x3907(x[3907]), .x3908(x[3908]), .x3909(x[3909]), .x3910(x[3910]), .x3911(x[3911]), .x3912(x[3912]), .x3913(x[3913]), .x3914(x[3914]), .x3915(x[3915]), .x3916(x[3916]), .x3917(x[3917]), .x3918(x[3918]), .x3919(x[3919]), .x3920(x[3920]), .x3921(x[3921]), .x3922(x[3922]), .x3923(x[3923]), .x3924(x[3924]), .x3925(x[3925]), .x3926(x[3926]), .x3927(x[3927]), .x3928(x[3928]), .x3929(x[3929]), .x3930(x[3930]), .x3931(x[3931]), .x3932(x[3932]), .x3933(x[3933]), .x3934(x[3934]), .x3935(x[3935]), .x3936(x[3936]), .x3937(x[3937]), .x3938(x[3938]), .x3939(x[3939]), .x3940(x[3940]), .x3941(x[3941]), .x3942(x[3942]), .x3943(x[3943]), .x3944(x[3944]), .x3945(x[3945]), .x3946(x[3946]), .x3947(x[3947]), .x3948(x[3948]), .x3949(x[3949]), .x3950(x[3950]), .x3951(x[3951]), .x3952(x[3952]), .x3953(x[3953]), .x3954(x[3954]), .x3955(x[3955]), .x3956(x[3956]), .x3957(x[3957]), .x3958(x[3958]), .x3959(x[3959]), .x3960(x[3960]), .x3961(x[3961]), .x3962(x[3962]), .x3963(x[3963]), .x3964(x[3964]), .x3965(x[3965]), .x3966(x[3966]), .x3967(x[3967]), .x3968(x[3968]), .x3969(x[3969]), .x3970(x[3970]), .x3971(x[3971]), .x3972(x[3972]), .x3973(x[3973]), .x3974(x[3974]), .x3975(x[3975]), .x3976(x[3976]), .x3977(x[3977]), .x3978(x[3978]), .x3979(x[3979]), .x3980(x[3980]), .x3981(x[3981]), .x3982(x[3982]), .x3983(x[3983]), .x3984(x[3984]), .x3985(x[3985]), .x3986(x[3986]), .x3987(x[3987]), .x3988(x[3988]), .x3989(x[3989]), .x3990(x[3990]), .x3991(x[3991]), .x3992(x[3992]), .x3993(x[3993]), .x3994(x[3994]), .x3995(x[3995]), .x3996(x[3996]), .x3997(x[3997]), .x3998(x[3998]), .x3999(x[3999]), .x4000(x[4000]), .x4001(x[4001]), .x4002(x[4002]), .x4003(x[4003]), .x4004(x[4004]), .x4005(x[4005]), .x4006(x[4006]), .x4007(x[4007]), .x4008(x[4008]), .x4009(x[4009]), .x4010(x[4010]), .x4011(x[4011]), .x4012(x[4012]), .x4013(x[4013]), .x4014(x[4014]), .x4015(x[4015]), .x4016(x[4016]), .x4017(x[4017]), .x4018(x[4018]), .x4019(x[4019]), .x4020(x[4020]), .x4021(x[4021]), .x4022(x[4022]), .x4023(x[4023]), .x4024(x[4024]), .x4025(x[4025]), .x4026(x[4026]), .x4027(x[4027]), .x4028(x[4028]), .x4029(x[4029]), .x4030(x[4030]), .x4031(x[4031]), .x4032(x[4032]), .x4033(x[4033]), .x4034(x[4034]), .x4035(x[4035]), .x4036(x[4036]), .x4037(x[4037]), .x4038(x[4038]), .x4039(x[4039]), .x4040(x[4040]), .x4041(x[4041]), .x4042(x[4042]), .x4043(x[4043]), .x4044(x[4044]), .x4045(x[4045]), .x4046(x[4046]), .x4047(x[4047]), .x4048(x[4048]), .x4049(x[4049]), .x4050(x[4050]), .x4051(x[4051]), .x4052(x[4052]), .x4053(x[4053]), .x4054(x[4054]), .x4055(x[4055]), .x4056(x[4056]), .x4057(x[4057]), .x4058(x[4058]), .x4059(x[4059]), .x4060(x[4060]), .x4061(x[4061]), .x4062(x[4062]), .x4063(x[4063]), .x4064(x[4064]), .x4065(x[4065]), .x4066(x[4066]), .x4067(x[4067]), .x4068(x[4068]), .x4069(x[4069]), .x4070(x[4070]), .x4071(x[4071]), .x4072(x[4072]), .x4073(x[4073]), .x4074(x[4074]), .x4075(x[4075]), .x4076(x[4076]), .x4077(x[4077]), .x4078(x[4078]), .x4079(x[4079]), .x4080(x[4080]), .x4081(x[4081]), .x4082(x[4082]), .x4083(x[4083]), .x4084(x[4084]), .x4085(x[4085]), .x4086(x[4086]), .x4087(x[4087]), .x4088(x[4088]), .x4089(x[4089]), .x4090(x[4090]), .x4091(x[4091]), .x4092(x[4092]), .x4093(x[4093]), .x4094(x[4094]), .x4095(x[4095]), .x4096(x[4096]), .x4097(x[4097]), .x4098(x[4098]), .x4099(x[4099]), .x4100(x[4100]), .x4101(x[4101]), .x4102(x[4102]), .x4103(x[4103]), .x4104(x[4104]), .x4105(x[4105]), .x4106(x[4106]), .x4107(x[4107]), .x4108(x[4108]), .x4109(x[4109]), .x4110(x[4110]), .x4111(x[4111]), .x4112(x[4112]), .x4113(x[4113]), .x4114(x[4114]), .x4115(x[4115]), .x4116(x[4116]), .x4117(x[4117]), .x4118(x[4118]), .x4119(x[4119]), .x4120(x[4120]), .x4121(x[4121]), .x4122(x[4122]), .x4123(x[4123]), .x4124(x[4124]), .x4125(x[4125]), .x4126(x[4126]), .x4127(x[4127]), .x4128(x[4128]), .x4129(x[4129]), .x4130(x[4130]), .x4131(x[4131]), .x4132(x[4132]), .x4133(x[4133]), .x4134(x[4134]), .x4135(x[4135]), .x4136(x[4136]), .x4137(x[4137]), .x4138(x[4138]), .x4139(x[4139]), .x4140(x[4140]), .x4141(x[4141]), .x4142(x[4142]), .x4143(x[4143]), .x4144(x[4144]), .x4145(x[4145]), .x4146(x[4146]), .x4147(x[4147]), .x4148(x[4148]), .x4149(x[4149]), .x4150(x[4150]), .x4151(x[4151]), .x4152(x[4152]), .x4153(x[4153]), .x4154(x[4154]), .x4155(x[4155]), .x4156(x[4156]), .x4157(x[4157]), .x4158(x[4158]), .x4159(x[4159]), .x4160(x[4160]), .x4161(x[4161]), .x4162(x[4162]), .x4163(x[4163]), .x4164(x[4164]), .x4165(x[4165]), .x4166(x[4166]), .x4167(x[4167]), .x4168(x[4168]), .x4169(x[4169]), .x4170(x[4170]), .x4171(x[4171]), .x4172(x[4172]), .x4173(x[4173]), .x4174(x[4174]), .x4175(x[4175]), .x4176(x[4176]), .x4177(x[4177]), .x4178(x[4178]), .x4179(x[4179]), .x4180(x[4180]), .x4181(x[4181]), .x4182(x[4182]), .x4183(x[4183]), .x4184(x[4184]), .x4185(x[4185]), .x4186(x[4186]), .x4187(x[4187]), .x4188(x[4188]), .x4189(x[4189]), .x4190(x[4190]), .x4191(x[4191]), .x4192(x[4192]), .x4193(x[4193]), .x4194(x[4194]), .x4195(x[4195]), .x4196(x[4196]), .x4197(x[4197]), .x4198(x[4198]), .x4199(x[4199]), .x4200(x[4200]), .x4201(x[4201]), .x4202(x[4202]), .x4203(x[4203]), .x4204(x[4204]), .x4205(x[4205]), .x4206(x[4206]), .x4207(x[4207]), .x4208(x[4208]), .x4209(x[4209]), .x4210(x[4210]), .x4211(x[4211]), .x4212(x[4212]), .x4213(x[4213]), .x4214(x[4214]), .x4215(x[4215]), .x4216(x[4216]), .x4217(x[4217]), .x4218(x[4218]), .x4219(x[4219]), .x4220(x[4220]), .x4221(x[4221]), .x4222(x[4222]), .x4223(x[4223]), .x4224(x[4224]), .x4225(x[4225]), .x4226(x[4226]), .x4227(x[4227]), .x4228(x[4228]), .x4229(x[4229]), .x4230(x[4230]), .x4231(x[4231]), .x4232(x[4232]), .x4233(x[4233]), .x4234(x[4234]), .x4235(x[4235]), .x4236(x[4236]), .x4237(x[4237]), .x4238(x[4238]), .x4239(x[4239]), .x4240(x[4240]), .x4241(x[4241]), .x4242(x[4242]), .x4243(x[4243]), .x4244(x[4244]), .x4245(x[4245]), .x4246(x[4246]), .x4247(x[4247]), .x4248(x[4248]), .x4249(x[4249]), .x4250(x[4250]), .x4251(x[4251]), .x4252(x[4252]), .x4253(x[4253]), .x4254(x[4254]), .x4255(x[4255]), .x4256(x[4256]), .x4257(x[4257]), .x4258(x[4258]), .x4259(x[4259]), .x4260(x[4260]), .x4261(x[4261]), .x4262(x[4262]), .x4263(x[4263]), .x4264(x[4264]), .x4265(x[4265]), .x4266(x[4266]), .x4267(x[4267]), .x4268(x[4268]), .x4269(x[4269]), .x4270(x[4270]), .x4271(x[4271]), .x4272(x[4272]), .x4273(x[4273]), .x4274(x[4274]), .x4275(x[4275]), .x4276(x[4276]), .x4277(x[4277]), .x4278(x[4278]), .x4279(x[4279]), .x4280(x[4280]), .x4281(x[4281]), .x4282(x[4282]), .x4283(x[4283]), .x4284(x[4284]), .x4285(x[4285]), .x4286(x[4286]), .x4287(x[4287]), .x4288(x[4288]), .x4289(x[4289]), .x4290(x[4290]), .x4291(x[4291]), .x4292(x[4292]), .x4293(x[4293]), .x4294(x[4294]), .x4295(x[4295]), .x4296(x[4296]), .x4297(x[4297]), .x4298(x[4298]), .x4299(x[4299]), .x4300(x[4300]), .x4301(x[4301]), .x4302(x[4302]), .x4303(x[4303]), .x4304(x[4304]), .x4305(x[4305]), .x4306(x[4306]), .x4307(x[4307]), .x4308(x[4308]), .x4309(x[4309]), .x4310(x[4310]), .x4311(x[4311]), .x4312(x[4312]), .x4313(x[4313]), .x4314(x[4314]), .x4315(x[4315]), .x4316(x[4316]), .x4317(x[4317]), .x4318(x[4318]), .x4319(x[4319]), .x4320(x[4320]), .x4321(x[4321]), .x4322(x[4322]), .x4323(x[4323]), .x4324(x[4324]), .x4325(x[4325]), .x4326(x[4326]), .x4327(x[4327]), .x4328(x[4328]), .x4329(x[4329]), .x4330(x[4330]), .x4331(x[4331]), .x4332(x[4332]), .x4333(x[4333]), .x4334(x[4334]), .x4335(x[4335]), .x4336(x[4336]), .x4337(x[4337]), .x4338(x[4338]), .x4339(x[4339]), .x4340(x[4340]), .x4341(x[4341]), .x4342(x[4342]), .x4343(x[4343]), .x4344(x[4344]), .x4345(x[4345]), .x4346(x[4346]), .x4347(x[4347]), .x4348(x[4348]), .x4349(x[4349]), .x4350(x[4350]), .x4351(x[4351]), .x4352(x[4352]), .x4353(x[4353]), .x4354(x[4354]), .x4355(x[4355]), .x4356(x[4356]), .x4357(x[4357]), .x4358(x[4358]), .x4359(x[4359]), .x4360(x[4360]), .x4361(x[4361]), .x4362(x[4362]), .x4363(x[4363]), .x4364(x[4364]), .x4365(x[4365]), .x4366(x[4366]), .x4367(x[4367]), .x4368(x[4368]), .x4369(x[4369]), .x4370(x[4370]), .x4371(x[4371]), .x4372(x[4372]), .x4373(x[4373]), .x4374(x[4374]), .x4375(x[4375]), .x4376(x[4376]), .x4377(x[4377]), .x4378(x[4378]), .x4379(x[4379]), .x4380(x[4380]), .x4381(x[4381]), .x4382(x[4382]), .x4383(x[4383]), .x4384(x[4384]), .x4385(x[4385]), .x4386(x[4386]), .x4387(x[4387]), .x4388(x[4388]), .x4389(x[4389]), .x4390(x[4390]), .x4391(x[4391]), .x4392(x[4392]), .x4393(x[4393]), .x4394(x[4394]), .x4395(x[4395]), .x4396(x[4396]), .x4397(x[4397]), .x4398(x[4398]), .x4399(x[4399]), .x4400(x[4400]), .x4401(x[4401]), .x4402(x[4402]), .x4403(x[4403]), .x4404(x[4404]), .x4405(x[4405]), .x4406(x[4406]), .x4407(x[4407]), .x4408(x[4408]), .x4409(x[4409]), .x4410(x[4410]), .x4411(x[4411]), .x4412(x[4412]), .x4413(x[4413]), .x4414(x[4414]), .x4415(x[4415]), .x4416(x[4416]), .x4417(x[4417]), .x4418(x[4418]), .x4419(x[4419]), .x4420(x[4420]), .x4421(x[4421]), .x4422(x[4422]), .x4423(x[4423]), .x4424(x[4424]), .x4425(x[4425]), .x4426(x[4426]), .x4427(x[4427]), .x4428(x[4428]), .x4429(x[4429]), .x4430(x[4430]), .x4431(x[4431]), .x4432(x[4432]), .x4433(x[4433]), .x4434(x[4434]), .x4435(x[4435]), .x4436(x[4436]), .x4437(x[4437]), .x4438(x[4438]), .x4439(x[4439]), .x4440(x[4440]), .x4441(x[4441]), .x4442(x[4442]), .x4443(x[4443]), .x4444(x[4444]), .x4445(x[4445]), .x4446(x[4446]), .x4447(x[4447]), .x4448(x[4448]), .x4449(x[4449]), .x4450(x[4450]), .x4451(x[4451]), .x4452(x[4452]), .x4453(x[4453]), .x4454(x[4454]), .x4455(x[4455]), .x4456(x[4456]), .x4457(x[4457]), .x4458(x[4458]), .x4459(x[4459]), .x4460(x[4460]), .x4461(x[4461]), .x4462(x[4462]), .x4463(x[4463]), .x4464(x[4464]), .x4465(x[4465]), .x4466(x[4466]), .x4467(x[4467]), .x4468(x[4468]), .x4469(x[4469]), .x4470(x[4470]), .x4471(x[4471]), .x4472(x[4472]), .x4473(x[4473]), .x4474(x[4474]), .x4475(x[4475]), .x4476(x[4476]), .x4477(x[4477]), .x4478(x[4478]), .x4479(x[4479]), .x4480(x[4480]), .x4481(x[4481]), .x4482(x[4482]), .x4483(x[4483]), .x4484(x[4484]), .x4485(x[4485]), .x4486(x[4486]), .x4487(x[4487]), .x4488(x[4488]), .x4489(x[4489]), .x4490(x[4490]), .x4491(x[4491]), .x4492(x[4492]), .x4493(x[4493]), .x4494(x[4494]), .x4495(x[4495]), .x4496(x[4496]), .x4497(x[4497]), .x4498(x[4498]), .x4499(x[4499]), .x4500(x[4500]), .x4501(x[4501]), .x4502(x[4502]), .x4503(x[4503]), .x4504(x[4504]), .x4505(x[4505]), .x4506(x[4506]), .x4507(x[4507]), .x4508(x[4508]), .x4509(x[4509]), .x4510(x[4510]), .x4511(x[4511]), .x4512(x[4512]), .x4513(x[4513]), .x4514(x[4514]), .x4515(x[4515]), .x4516(x[4516]), .x4517(x[4517]), .x4518(x[4518]), .x4519(x[4519]), .x4520(x[4520]), .x4521(x[4521]), .x4522(x[4522]), .x4523(x[4523]), .x4524(x[4524]), .x4525(x[4525]), .x4526(x[4526]), .x4527(x[4527]), .x4528(x[4528]), .x4529(x[4529]), .x4530(x[4530]), .x4531(x[4531]), .x4532(x[4532]), .x4533(x[4533]), .x4534(x[4534]), .x4535(x[4535]), .x4536(x[4536]), .x4537(x[4537]), .x4538(x[4538]), .x4539(x[4539]), .x4540(x[4540]), .x4541(x[4541]), .x4542(x[4542]), .x4543(x[4543]), .x4544(x[4544]), .x4545(x[4545]), .x4546(x[4546]), .x4547(x[4547]), .x4548(x[4548]), .x4549(x[4549]), .x4550(x[4550]), .x4551(x[4551]), .x4552(x[4552]), .x4553(x[4553]), .x4554(x[4554]), .x4555(x[4555]), .x4556(x[4556]), .x4557(x[4557]), .x4558(x[4558]), .x4559(x[4559]), .x4560(x[4560]), .x4561(x[4561]), .x4562(x[4562]), .x4563(x[4563]), .x4564(x[4564]), .x4565(x[4565]), .x4566(x[4566]), .x4567(x[4567]), .x4568(x[4568]), .x4569(x[4569]), .x4570(x[4570]), .x4571(x[4571]), .x4572(x[4572]), .x4573(x[4573]), .x4574(x[4574]), .x4575(x[4575]), .x4576(x[4576]), .x4577(x[4577]), .x4578(x[4578]), .x4579(x[4579]), .x4580(x[4580]), .x4581(x[4581]), .x4582(x[4582]), .x4583(x[4583]), .x4584(x[4584]), .x4585(x[4585]), .x4586(x[4586]), .x4587(x[4587]), .x4588(x[4588]), .x4589(x[4589]), .x4590(x[4590]), .x4591(x[4591]), .x4592(x[4592]), .x4593(x[4593]), .x4594(x[4594]), .x4595(x[4595]), .x4596(x[4596]), .x4597(x[4597]), .x4598(x[4598]), .x4599(x[4599]), .x4600(x[4600]), .x4601(x[4601]), .x4602(x[4602]), .x4603(x[4603]), .x4604(x[4604]), .x4605(x[4605]), .x4606(x[4606]), .x4607(x[4607]), .x4608(x[4608]), .x4609(x[4609]), .x4610(x[4610]), .x4611(x[4611]), .x4612(x[4612]), .x4613(x[4613]), .x4614(x[4614]), .x4615(x[4615]), .x4616(x[4616]), .x4617(x[4617]), .x4618(x[4618]), .x4619(x[4619]), .x4620(x[4620]), .x4621(x[4621]), .x4622(x[4622]), .x4623(x[4623]), .x4624(x[4624]), .x4625(x[4625]), .x4626(x[4626]), .x4627(x[4627]), .x4628(x[4628]), .x4629(x[4629]), .x4630(x[4630]), .x4631(x[4631]), .x4632(x[4632]), .x4633(x[4633]), .x4634(x[4634]), .x4635(x[4635]), .x4636(x[4636]), .x4637(x[4637]), .x4638(x[4638]), .x4639(x[4639]), .x4640(x[4640]), .x4641(x[4641]), .x4642(x[4642]), .x4643(x[4643]), .x4644(x[4644]), .x4645(x[4645]), .x4646(x[4646]), .x4647(x[4647]), .x4648(x[4648]), .x4649(x[4649]), .x4650(x[4650]), .x4651(x[4651]), .x4652(x[4652]), .x4653(x[4653]), .x4654(x[4654]), .x4655(x[4655]), .x4656(x[4656]), .x4657(x[4657]), .x4658(x[4658]), .x4659(x[4659]), .x4660(x[4660]), .x4661(x[4661]), .x4662(x[4662]), .x4663(x[4663]), .x4664(x[4664]), .x4665(x[4665]), .x4666(x[4666]), .x4667(x[4667]), .x4668(x[4668]), .x4669(x[4669]), .x4670(x[4670]), .x4671(x[4671]), .x4672(x[4672]), .x4673(x[4673]), .x4674(x[4674]), .x4675(x[4675]), .x4676(x[4676]), .x4677(x[4677]), .x4678(x[4678]), .x4679(x[4679]), .x4680(x[4680]), .x4681(x[4681]), .x4682(x[4682]), .x4683(x[4683]), .x4684(x[4684]), .x4685(x[4685]), .x4686(x[4686]), .x4687(x[4687]), .x4688(x[4688]), .x4689(x[4689]), .x4690(x[4690]), .x4691(x[4691]), .x4692(x[4692]), .x4693(x[4693]), .x4694(x[4694]), .x4695(x[4695]), .x4696(x[4696]), .x4697(x[4697]), .x4698(x[4698]), .x4699(x[4699]), .x4700(x[4700]), .x4701(x[4701]), .x4702(x[4702]), .x4703(x[4703]), .x4704(x[4704]), .x4705(x[4705]), .x4706(x[4706]), .x4707(x[4707]), .x4708(x[4708]), .x4709(x[4709]), .x4710(x[4710]), .x4711(x[4711]), .x4712(x[4712]), .x4713(x[4713]), .x4714(x[4714]), .x4715(x[4715]), .x4716(x[4716]), .x4717(x[4717]), .x4718(x[4718]), .x4719(x[4719]), .x4720(x[4720]), .x4721(x[4721]), .x4722(x[4722]), .x4723(x[4723]), .x4724(x[4724]), .x4725(x[4725]), .x4726(x[4726]), .x4727(x[4727]), .x4728(x[4728]), .x4729(x[4729]), .x4730(x[4730]), .x4731(x[4731]), .x4732(x[4732]), .x4733(x[4733]), .x4734(x[4734]), .x4735(x[4735]), .x4736(x[4736]), .x4737(x[4737]), .x4738(x[4738]), .x4739(x[4739]), .x4740(x[4740]), .x4741(x[4741]), .x4742(x[4742]), .x4743(x[4743]), .x4744(x[4744]), .x4745(x[4745]), .x4746(x[4746]), .x4747(x[4747]), .x4748(x[4748]), .x4749(x[4749]), .x4750(x[4750]), .x4751(x[4751]), .x4752(x[4752]), .x4753(x[4753]), .x4754(x[4754]), .x4755(x[4755]), .x4756(x[4756]), .x4757(x[4757]), .x4758(x[4758]), .x4759(x[4759]), .x4760(x[4760]), .x4761(x[4761]), .x4762(x[4762]), .x4763(x[4763]), .x4764(x[4764]), .x4765(x[4765]), .x4766(x[4766]), .x4767(x[4767]), .x4768(x[4768]), .x4769(x[4769]), .x4770(x[4770]), .x4771(x[4771]), .x4772(x[4772]), .x4773(x[4773]), .x4774(x[4774]), .x4775(x[4775]), .x4776(x[4776]), .x4777(x[4777]), .x4778(x[4778]), .x4779(x[4779]), .x4780(x[4780]), .x4781(x[4781]), .x4782(x[4782]), .x4783(x[4783]), .x4784(x[4784]), .x4785(x[4785]), .x4786(x[4786]), .x4787(x[4787]), .x4788(x[4788]), .x4789(x[4789]), .x4790(x[4790]), .x4791(x[4791]), .x4792(x[4792]), .x4793(x[4793]), .x4794(x[4794]), .x4795(x[4795]), .x4796(x[4796]), .x4797(x[4797]), .x4798(x[4798]), .x4799(x[4799]), .x4800(x[4800]), .x4801(x[4801]), .x4802(x[4802]), .x4803(x[4803]), .x4804(x[4804]), .x4805(x[4805]), .x4806(x[4806]), .x4807(x[4807]), .x4808(x[4808]), .x4809(x[4809]), .x4810(x[4810]), .x4811(x[4811]), .x4812(x[4812]), .x4813(x[4813]), .x4814(x[4814]), .x4815(x[4815]), .x4816(x[4816]), .x4817(x[4817]), .x4818(x[4818]), .x4819(x[4819]), .x4820(x[4820]), .x4821(x[4821]), .x4822(x[4822]), .x4823(x[4823]), .x4824(x[4824]), .x4825(x[4825]), .x4826(x[4826]), .x4827(x[4827]), .x4828(x[4828]), .x4829(x[4829]), .x4830(x[4830]), .x4831(x[4831]), .x4832(x[4832]), .x4833(x[4833]), .x4834(x[4834]), .x4835(x[4835]), .x4836(x[4836]), .x4837(x[4837]), .x4838(x[4838]), .x4839(x[4839]), .x4840(x[4840]), .x4841(x[4841]), .x4842(x[4842]), .x4843(x[4843]), .x4844(x[4844]), .x4845(x[4845]), .x4846(x[4846]), .x4847(x[4847]), .x4848(x[4848]), .x4849(x[4849]), .x4850(x[4850]), .x4851(x[4851]), .x4852(x[4852]), .x4853(x[4853]), .x4854(x[4854]), .x4855(x[4855]), .x4856(x[4856]), .x4857(x[4857]), .x4858(x[4858]), .x4859(x[4859]), .x4860(x[4860]), .x4861(x[4861]), .x4862(x[4862]), .x4863(x[4863]), .x4864(x[4864]), .x4865(x[4865]), .x4866(x[4866]), .x4867(x[4867]), .x4868(x[4868]), .x4869(x[4869]), .x4870(x[4870]), .x4871(x[4871]), .x4872(x[4872]), .x4873(x[4873]), .x4874(x[4874]), .x4875(x[4875]), .x4876(x[4876]), .x4877(x[4877]), .x4878(x[4878]), .x4879(x[4879]), .x4880(x[4880]), .x4881(x[4881]), .x4882(x[4882]), .x4883(x[4883]), .x4884(x[4884]), .x4885(x[4885]), .x4886(x[4886]), .x4887(x[4887]), .x4888(x[4888]), .x4889(x[4889]), .x4890(x[4890]), .x4891(x[4891]), .x4892(x[4892]), .x4893(x[4893]), .x4894(x[4894]), .x4895(x[4895]), .x4896(x[4896]), .x4897(x[4897]), .x4898(x[4898]), .x4899(x[4899]), .x4900(x[4900]), .x4901(x[4901]), .x4902(x[4902]), .x4903(x[4903]), .x4904(x[4904]), .x4905(x[4905]), .x4906(x[4906]), .x4907(x[4907]), .x4908(x[4908]), .x4909(x[4909]), .x4910(x[4910]), .x4911(x[4911]), .x4912(x[4912]), .x4913(x[4913]), .x4914(x[4914]), .x4915(x[4915]), .x4916(x[4916]), .x4917(x[4917]), .x4918(x[4918]), .x4919(x[4919]), .x4920(x[4920]), .x4921(x[4921]), .x4922(x[4922]), .x4923(x[4923]), .x4924(x[4924]), .x4925(x[4925]), .x4926(x[4926]), .x4927(x[4927]), .x4928(x[4928]), .x4929(x[4929]), .x4930(x[4930]), .x4931(x[4931]), .x4932(x[4932]), .x4933(x[4933]), .x4934(x[4934]), .x4935(x[4935]), .x4936(x[4936]), .x4937(x[4937]), .x4938(x[4938]), .x4939(x[4939]), .x4940(x[4940]), .x4941(x[4941]), .x4942(x[4942]), .x4943(x[4943]), .x4944(x[4944]), .x4945(x[4945]), .x4946(x[4946]), .x4947(x[4947]), .x4948(x[4948]), .x4949(x[4949]), .x4950(x[4950]), .x4951(x[4951]), .x4952(x[4952]), .x4953(x[4953]), .x4954(x[4954]), .x4955(x[4955]), .x4956(x[4956]), .x4957(x[4957]), .x4958(x[4958]), .x4959(x[4959]), .x4960(x[4960]), .x4961(x[4961]), .x4962(x[4962]), .x4963(x[4963]), .x4964(x[4964]), .x4965(x[4965]), .x4966(x[4966]), .x4967(x[4967]), .x4968(x[4968]), .x4969(x[4969]), .x4970(x[4970]), .x4971(x[4971]), .x4972(x[4972]), .x4973(x[4973]), .x4974(x[4974]), .x4975(x[4975]), .x4976(x[4976]), .x4977(x[4977]), .x4978(x[4978]), .x4979(x[4979]), .x4980(x[4980]), .x4981(x[4981]), .x4982(x[4982]), .x4983(x[4983]), .x4984(x[4984]), .x4985(x[4985]), .x4986(x[4986]), .x4987(x[4987]), .x4988(x[4988]), .x4989(x[4989]), .x4990(x[4990]), .x4991(x[4991]), .x4992(x[4992]), .x4993(x[4993]), .x4994(x[4994]), .x4995(x[4995]), .x4996(x[4996]), .x4997(x[4997]), .x4998(x[4998]), .x4999(x[4999]), .x5000(x[5000]), .x5001(x[5001]), .x5002(x[5002]), .x5003(x[5003]), .x5004(x[5004]), .x5005(x[5005]), .x5006(x[5006]), .x5007(x[5007]), .x5008(x[5008]), .x5009(x[5009]), .x5010(x[5010]), .x5011(x[5011]), .x5012(x[5012]), .x5013(x[5013]), .x5014(x[5014]), .x5015(x[5015]), .x5016(x[5016]), .x5017(x[5017]), .x5018(x[5018]), .x5019(x[5019]), .x5020(x[5020]), .x5021(x[5021]), .x5022(x[5022]), .x5023(x[5023]), .x5024(x[5024]),
    .y0(y0)
  );

  // Optional reference function (majority reference for sanity check)
  function [12:0] popcount(input [5024:0] v);
    integer i; reg [12:0] c;
    begin
      c = 0;
      for (i = 0; i < 5025; i = i + 1)
        c = c + v[i];
      popcount = c;
    end
  endfunction

  // Reference majority: at least 2513 ones
  wire y_ref = (popcount(x) >= 2513);

  localparam [63:0] TOTAL_VECTORS = 64'd4739452898216418547201653797763595860957428722528977235532895354610283334595157992601954763893350737531098159036292099891217849718658132949599338305423909899252433568409523604296927531388595995903212328377859293925028196664665449850920047372460929548959622342553774931470029996136721692487549847800783165669065600283216761882728648823088672849767761096787054409317648768673870046197091729852874525071048417569058029910574146116161366297222991158549940296605431801079820504387040532005678479769096620906801991999931319916541911339092108224127155815316085299843959201857069250074266999672661907812994957711857222227385566463837903557701706172013317028659878977488721010157415572005239921821872642128383718566810743592190387800338965309406435642999976013852377063915568381663822154853706240880713672399028318733383264792633014849194780378227897156978938757328083522020917300464403999534043883489380242875421456525648278512104832460583690257724803208284252160095154337085117492746715082940721986813303177842688134816866983859627735702246922741856296160056654162807679644176131822175861244568214031779577836287324457834556298882134763531751909360525557572719095658843766275014763096181817096664181823043722510021319610830579781988247221574674180784741135629303528577581367198572085824120663747784090886290823216458725893664233566807777314155339529598238740914418234871716424282967739043062987444191457487347008423479118751929185205742311071535373987016939985312505575666322649798388484889607881003797682733554107154432;

  initial begin
    $display("Time | x5024 x5023 x5022 x5021 x5020 x5019 x5018 x5017 x5016 x5015 x5014 x5013 x5012 x5011 x5010 x5009 x5008 x5007 x5006 x5005 x5004 x5003 x5002 x5001 x5000 x4999 x4998 x4997 x4996 x4995 x4994 x4993 x4992 x4991 x4990 x4989 x4988 x4987 x4986 x4985 x4984 x4983 x4982 x4981 x4980 x4979 x4978 x4977 x4976 x4975 x4974 x4973 x4972 x4971 x4970 x4969 x4968 x4967 x4966 x4965 x4964 x4963 x4962 x4961 x4960 x4959 x4958 x4957 x4956 x4955 x4954 x4953 x4952 x4951 x4950 x4949 x4948 x4947 x4946 x4945 x4944 x4943 x4942 x4941 x4940 x4939 x4938 x4937 x4936 x4935 x4934 x4933 x4932 x4931 x4930 x4929 x4928 x4927 x4926 x4925 x4924 x4923 x4922 x4921 x4920 x4919 x4918 x4917 x4916 x4915 x4914 x4913 x4912 x4911 x4910 x4909 x4908 x4907 x4906 x4905 x4904 x4903 x4902 x4901 x4900 x4899 x4898 x4897 x4896 x4895 x4894 x4893 x4892 x4891 x4890 x4889 x4888 x4887 x4886 x4885 x4884 x4883 x4882 x4881 x4880 x4879 x4878 x4877 x4876 x4875 x4874 x4873 x4872 x4871 x4870 x4869 x4868 x4867 x4866 x4865 x4864 x4863 x4862 x4861 x4860 x4859 x4858 x4857 x4856 x4855 x4854 x4853 x4852 x4851 x4850 x4849 x4848 x4847 x4846 x4845 x4844 x4843 x4842 x4841 x4840 x4839 x4838 x4837 x4836 x4835 x4834 x4833 x4832 x4831 x4830 x4829 x4828 x4827 x4826 x4825 x4824 x4823 x4822 x4821 x4820 x4819 x4818 x4817 x4816 x4815 x4814 x4813 x4812 x4811 x4810 x4809 x4808 x4807 x4806 x4805 x4804 x4803 x4802 x4801 x4800 x4799 x4798 x4797 x4796 x4795 x4794 x4793 x4792 x4791 x4790 x4789 x4788 x4787 x4786 x4785 x4784 x4783 x4782 x4781 x4780 x4779 x4778 x4777 x4776 x4775 x4774 x4773 x4772 x4771 x4770 x4769 x4768 x4767 x4766 x4765 x4764 x4763 x4762 x4761 x4760 x4759 x4758 x4757 x4756 x4755 x4754 x4753 x4752 x4751 x4750 x4749 x4748 x4747 x4746 x4745 x4744 x4743 x4742 x4741 x4740 x4739 x4738 x4737 x4736 x4735 x4734 x4733 x4732 x4731 x4730 x4729 x4728 x4727 x4726 x4725 x4724 x4723 x4722 x4721 x4720 x4719 x4718 x4717 x4716 x4715 x4714 x4713 x4712 x4711 x4710 x4709 x4708 x4707 x4706 x4705 x4704 x4703 x4702 x4701 x4700 x4699 x4698 x4697 x4696 x4695 x4694 x4693 x4692 x4691 x4690 x4689 x4688 x4687 x4686 x4685 x4684 x4683 x4682 x4681 x4680 x4679 x4678 x4677 x4676 x4675 x4674 x4673 x4672 x4671 x4670 x4669 x4668 x4667 x4666 x4665 x4664 x4663 x4662 x4661 x4660 x4659 x4658 x4657 x4656 x4655 x4654 x4653 x4652 x4651 x4650 x4649 x4648 x4647 x4646 x4645 x4644 x4643 x4642 x4641 x4640 x4639 x4638 x4637 x4636 x4635 x4634 x4633 x4632 x4631 x4630 x4629 x4628 x4627 x4626 x4625 x4624 x4623 x4622 x4621 x4620 x4619 x4618 x4617 x4616 x4615 x4614 x4613 x4612 x4611 x4610 x4609 x4608 x4607 x4606 x4605 x4604 x4603 x4602 x4601 x4600 x4599 x4598 x4597 x4596 x4595 x4594 x4593 x4592 x4591 x4590 x4589 x4588 x4587 x4586 x4585 x4584 x4583 x4582 x4581 x4580 x4579 x4578 x4577 x4576 x4575 x4574 x4573 x4572 x4571 x4570 x4569 x4568 x4567 x4566 x4565 x4564 x4563 x4562 x4561 x4560 x4559 x4558 x4557 x4556 x4555 x4554 x4553 x4552 x4551 x4550 x4549 x4548 x4547 x4546 x4545 x4544 x4543 x4542 x4541 x4540 x4539 x4538 x4537 x4536 x4535 x4534 x4533 x4532 x4531 x4530 x4529 x4528 x4527 x4526 x4525 x4524 x4523 x4522 x4521 x4520 x4519 x4518 x4517 x4516 x4515 x4514 x4513 x4512 x4511 x4510 x4509 x4508 x4507 x4506 x4505 x4504 x4503 x4502 x4501 x4500 x4499 x4498 x4497 x4496 x4495 x4494 x4493 x4492 x4491 x4490 x4489 x4488 x4487 x4486 x4485 x4484 x4483 x4482 x4481 x4480 x4479 x4478 x4477 x4476 x4475 x4474 x4473 x4472 x4471 x4470 x4469 x4468 x4467 x4466 x4465 x4464 x4463 x4462 x4461 x4460 x4459 x4458 x4457 x4456 x4455 x4454 x4453 x4452 x4451 x4450 x4449 x4448 x4447 x4446 x4445 x4444 x4443 x4442 x4441 x4440 x4439 x4438 x4437 x4436 x4435 x4434 x4433 x4432 x4431 x4430 x4429 x4428 x4427 x4426 x4425 x4424 x4423 x4422 x4421 x4420 x4419 x4418 x4417 x4416 x4415 x4414 x4413 x4412 x4411 x4410 x4409 x4408 x4407 x4406 x4405 x4404 x4403 x4402 x4401 x4400 x4399 x4398 x4397 x4396 x4395 x4394 x4393 x4392 x4391 x4390 x4389 x4388 x4387 x4386 x4385 x4384 x4383 x4382 x4381 x4380 x4379 x4378 x4377 x4376 x4375 x4374 x4373 x4372 x4371 x4370 x4369 x4368 x4367 x4366 x4365 x4364 x4363 x4362 x4361 x4360 x4359 x4358 x4357 x4356 x4355 x4354 x4353 x4352 x4351 x4350 x4349 x4348 x4347 x4346 x4345 x4344 x4343 x4342 x4341 x4340 x4339 x4338 x4337 x4336 x4335 x4334 x4333 x4332 x4331 x4330 x4329 x4328 x4327 x4326 x4325 x4324 x4323 x4322 x4321 x4320 x4319 x4318 x4317 x4316 x4315 x4314 x4313 x4312 x4311 x4310 x4309 x4308 x4307 x4306 x4305 x4304 x4303 x4302 x4301 x4300 x4299 x4298 x4297 x4296 x4295 x4294 x4293 x4292 x4291 x4290 x4289 x4288 x4287 x4286 x4285 x4284 x4283 x4282 x4281 x4280 x4279 x4278 x4277 x4276 x4275 x4274 x4273 x4272 x4271 x4270 x4269 x4268 x4267 x4266 x4265 x4264 x4263 x4262 x4261 x4260 x4259 x4258 x4257 x4256 x4255 x4254 x4253 x4252 x4251 x4250 x4249 x4248 x4247 x4246 x4245 x4244 x4243 x4242 x4241 x4240 x4239 x4238 x4237 x4236 x4235 x4234 x4233 x4232 x4231 x4230 x4229 x4228 x4227 x4226 x4225 x4224 x4223 x4222 x4221 x4220 x4219 x4218 x4217 x4216 x4215 x4214 x4213 x4212 x4211 x4210 x4209 x4208 x4207 x4206 x4205 x4204 x4203 x4202 x4201 x4200 x4199 x4198 x4197 x4196 x4195 x4194 x4193 x4192 x4191 x4190 x4189 x4188 x4187 x4186 x4185 x4184 x4183 x4182 x4181 x4180 x4179 x4178 x4177 x4176 x4175 x4174 x4173 x4172 x4171 x4170 x4169 x4168 x4167 x4166 x4165 x4164 x4163 x4162 x4161 x4160 x4159 x4158 x4157 x4156 x4155 x4154 x4153 x4152 x4151 x4150 x4149 x4148 x4147 x4146 x4145 x4144 x4143 x4142 x4141 x4140 x4139 x4138 x4137 x4136 x4135 x4134 x4133 x4132 x4131 x4130 x4129 x4128 x4127 x4126 x4125 x4124 x4123 x4122 x4121 x4120 x4119 x4118 x4117 x4116 x4115 x4114 x4113 x4112 x4111 x4110 x4109 x4108 x4107 x4106 x4105 x4104 x4103 x4102 x4101 x4100 x4099 x4098 x4097 x4096 x4095 x4094 x4093 x4092 x4091 x4090 x4089 x4088 x4087 x4086 x4085 x4084 x4083 x4082 x4081 x4080 x4079 x4078 x4077 x4076 x4075 x4074 x4073 x4072 x4071 x4070 x4069 x4068 x4067 x4066 x4065 x4064 x4063 x4062 x4061 x4060 x4059 x4058 x4057 x4056 x4055 x4054 x4053 x4052 x4051 x4050 x4049 x4048 x4047 x4046 x4045 x4044 x4043 x4042 x4041 x4040 x4039 x4038 x4037 x4036 x4035 x4034 x4033 x4032 x4031 x4030 x4029 x4028 x4027 x4026 x4025 x4024 x4023 x4022 x4021 x4020 x4019 x4018 x4017 x4016 x4015 x4014 x4013 x4012 x4011 x4010 x4009 x4008 x4007 x4006 x4005 x4004 x4003 x4002 x4001 x4000 x3999 x3998 x3997 x3996 x3995 x3994 x3993 x3992 x3991 x3990 x3989 x3988 x3987 x3986 x3985 x3984 x3983 x3982 x3981 x3980 x3979 x3978 x3977 x3976 x3975 x3974 x3973 x3972 x3971 x3970 x3969 x3968 x3967 x3966 x3965 x3964 x3963 x3962 x3961 x3960 x3959 x3958 x3957 x3956 x3955 x3954 x3953 x3952 x3951 x3950 x3949 x3948 x3947 x3946 x3945 x3944 x3943 x3942 x3941 x3940 x3939 x3938 x3937 x3936 x3935 x3934 x3933 x3932 x3931 x3930 x3929 x3928 x3927 x3926 x3925 x3924 x3923 x3922 x3921 x3920 x3919 x3918 x3917 x3916 x3915 x3914 x3913 x3912 x3911 x3910 x3909 x3908 x3907 x3906 x3905 x3904 x3903 x3902 x3901 x3900 x3899 x3898 x3897 x3896 x3895 x3894 x3893 x3892 x3891 x3890 x3889 x3888 x3887 x3886 x3885 x3884 x3883 x3882 x3881 x3880 x3879 x3878 x3877 x3876 x3875 x3874 x3873 x3872 x3871 x3870 x3869 x3868 x3867 x3866 x3865 x3864 x3863 x3862 x3861 x3860 x3859 x3858 x3857 x3856 x3855 x3854 x3853 x3852 x3851 x3850 x3849 x3848 x3847 x3846 x3845 x3844 x3843 x3842 x3841 x3840 x3839 x3838 x3837 x3836 x3835 x3834 x3833 x3832 x3831 x3830 x3829 x3828 x3827 x3826 x3825 x3824 x3823 x3822 x3821 x3820 x3819 x3818 x3817 x3816 x3815 x3814 x3813 x3812 x3811 x3810 x3809 x3808 x3807 x3806 x3805 x3804 x3803 x3802 x3801 x3800 x3799 x3798 x3797 x3796 x3795 x3794 x3793 x3792 x3791 x3790 x3789 x3788 x3787 x3786 x3785 x3784 x3783 x3782 x3781 x3780 x3779 x3778 x3777 x3776 x3775 x3774 x3773 x3772 x3771 x3770 x3769 x3768 x3767 x3766 x3765 x3764 x3763 x3762 x3761 x3760 x3759 x3758 x3757 x3756 x3755 x3754 x3753 x3752 x3751 x3750 x3749 x3748 x3747 x3746 x3745 x3744 x3743 x3742 x3741 x3740 x3739 x3738 x3737 x3736 x3735 x3734 x3733 x3732 x3731 x3730 x3729 x3728 x3727 x3726 x3725 x3724 x3723 x3722 x3721 x3720 x3719 x3718 x3717 x3716 x3715 x3714 x3713 x3712 x3711 x3710 x3709 x3708 x3707 x3706 x3705 x3704 x3703 x3702 x3701 x3700 x3699 x3698 x3697 x3696 x3695 x3694 x3693 x3692 x3691 x3690 x3689 x3688 x3687 x3686 x3685 x3684 x3683 x3682 x3681 x3680 x3679 x3678 x3677 x3676 x3675 x3674 x3673 x3672 x3671 x3670 x3669 x3668 x3667 x3666 x3665 x3664 x3663 x3662 x3661 x3660 x3659 x3658 x3657 x3656 x3655 x3654 x3653 x3652 x3651 x3650 x3649 x3648 x3647 x3646 x3645 x3644 x3643 x3642 x3641 x3640 x3639 x3638 x3637 x3636 x3635 x3634 x3633 x3632 x3631 x3630 x3629 x3628 x3627 x3626 x3625 x3624 x3623 x3622 x3621 x3620 x3619 x3618 x3617 x3616 x3615 x3614 x3613 x3612 x3611 x3610 x3609 x3608 x3607 x3606 x3605 x3604 x3603 x3602 x3601 x3600 x3599 x3598 x3597 x3596 x3595 x3594 x3593 x3592 x3591 x3590 x3589 x3588 x3587 x3586 x3585 x3584 x3583 x3582 x3581 x3580 x3579 x3578 x3577 x3576 x3575 x3574 x3573 x3572 x3571 x3570 x3569 x3568 x3567 x3566 x3565 x3564 x3563 x3562 x3561 x3560 x3559 x3558 x3557 x3556 x3555 x3554 x3553 x3552 x3551 x3550 x3549 x3548 x3547 x3546 x3545 x3544 x3543 x3542 x3541 x3540 x3539 x3538 x3537 x3536 x3535 x3534 x3533 x3532 x3531 x3530 x3529 x3528 x3527 x3526 x3525 x3524 x3523 x3522 x3521 x3520 x3519 x3518 x3517 x3516 x3515 x3514 x3513 x3512 x3511 x3510 x3509 x3508 x3507 x3506 x3505 x3504 x3503 x3502 x3501 x3500 x3499 x3498 x3497 x3496 x3495 x3494 x3493 x3492 x3491 x3490 x3489 x3488 x3487 x3486 x3485 x3484 x3483 x3482 x3481 x3480 x3479 x3478 x3477 x3476 x3475 x3474 x3473 x3472 x3471 x3470 x3469 x3468 x3467 x3466 x3465 x3464 x3463 x3462 x3461 x3460 x3459 x3458 x3457 x3456 x3455 x3454 x3453 x3452 x3451 x3450 x3449 x3448 x3447 x3446 x3445 x3444 x3443 x3442 x3441 x3440 x3439 x3438 x3437 x3436 x3435 x3434 x3433 x3432 x3431 x3430 x3429 x3428 x3427 x3426 x3425 x3424 x3423 x3422 x3421 x3420 x3419 x3418 x3417 x3416 x3415 x3414 x3413 x3412 x3411 x3410 x3409 x3408 x3407 x3406 x3405 x3404 x3403 x3402 x3401 x3400 x3399 x3398 x3397 x3396 x3395 x3394 x3393 x3392 x3391 x3390 x3389 x3388 x3387 x3386 x3385 x3384 x3383 x3382 x3381 x3380 x3379 x3378 x3377 x3376 x3375 x3374 x3373 x3372 x3371 x3370 x3369 x3368 x3367 x3366 x3365 x3364 x3363 x3362 x3361 x3360 x3359 x3358 x3357 x3356 x3355 x3354 x3353 x3352 x3351 x3350 x3349 x3348 x3347 x3346 x3345 x3344 x3343 x3342 x3341 x3340 x3339 x3338 x3337 x3336 x3335 x3334 x3333 x3332 x3331 x3330 x3329 x3328 x3327 x3326 x3325 x3324 x3323 x3322 x3321 x3320 x3319 x3318 x3317 x3316 x3315 x3314 x3313 x3312 x3311 x3310 x3309 x3308 x3307 x3306 x3305 x3304 x3303 x3302 x3301 x3300 x3299 x3298 x3297 x3296 x3295 x3294 x3293 x3292 x3291 x3290 x3289 x3288 x3287 x3286 x3285 x3284 x3283 x3282 x3281 x3280 x3279 x3278 x3277 x3276 x3275 x3274 x3273 x3272 x3271 x3270 x3269 x3268 x3267 x3266 x3265 x3264 x3263 x3262 x3261 x3260 x3259 x3258 x3257 x3256 x3255 x3254 x3253 x3252 x3251 x3250 x3249 x3248 x3247 x3246 x3245 x3244 x3243 x3242 x3241 x3240 x3239 x3238 x3237 x3236 x3235 x3234 x3233 x3232 x3231 x3230 x3229 x3228 x3227 x3226 x3225 x3224 x3223 x3222 x3221 x3220 x3219 x3218 x3217 x3216 x3215 x3214 x3213 x3212 x3211 x3210 x3209 x3208 x3207 x3206 x3205 x3204 x3203 x3202 x3201 x3200 x3199 x3198 x3197 x3196 x3195 x3194 x3193 x3192 x3191 x3190 x3189 x3188 x3187 x3186 x3185 x3184 x3183 x3182 x3181 x3180 x3179 x3178 x3177 x3176 x3175 x3174 x3173 x3172 x3171 x3170 x3169 x3168 x3167 x3166 x3165 x3164 x3163 x3162 x3161 x3160 x3159 x3158 x3157 x3156 x3155 x3154 x3153 x3152 x3151 x3150 x3149 x3148 x3147 x3146 x3145 x3144 x3143 x3142 x3141 x3140 x3139 x3138 x3137 x3136 x3135 x3134 x3133 x3132 x3131 x3130 x3129 x3128 x3127 x3126 x3125 x3124 x3123 x3122 x3121 x3120 x3119 x3118 x3117 x3116 x3115 x3114 x3113 x3112 x3111 x3110 x3109 x3108 x3107 x3106 x3105 x3104 x3103 x3102 x3101 x3100 x3099 x3098 x3097 x3096 x3095 x3094 x3093 x3092 x3091 x3090 x3089 x3088 x3087 x3086 x3085 x3084 x3083 x3082 x3081 x3080 x3079 x3078 x3077 x3076 x3075 x3074 x3073 x3072 x3071 x3070 x3069 x3068 x3067 x3066 x3065 x3064 x3063 x3062 x3061 x3060 x3059 x3058 x3057 x3056 x3055 x3054 x3053 x3052 x3051 x3050 x3049 x3048 x3047 x3046 x3045 x3044 x3043 x3042 x3041 x3040 x3039 x3038 x3037 x3036 x3035 x3034 x3033 x3032 x3031 x3030 x3029 x3028 x3027 x3026 x3025 x3024 x3023 x3022 x3021 x3020 x3019 x3018 x3017 x3016 x3015 x3014 x3013 x3012 x3011 x3010 x3009 x3008 x3007 x3006 x3005 x3004 x3003 x3002 x3001 x3000 x2999 x2998 x2997 x2996 x2995 x2994 x2993 x2992 x2991 x2990 x2989 x2988 x2987 x2986 x2985 x2984 x2983 x2982 x2981 x2980 x2979 x2978 x2977 x2976 x2975 x2974 x2973 x2972 x2971 x2970 x2969 x2968 x2967 x2966 x2965 x2964 x2963 x2962 x2961 x2960 x2959 x2958 x2957 x2956 x2955 x2954 x2953 x2952 x2951 x2950 x2949 x2948 x2947 x2946 x2945 x2944 x2943 x2942 x2941 x2940 x2939 x2938 x2937 x2936 x2935 x2934 x2933 x2932 x2931 x2930 x2929 x2928 x2927 x2926 x2925 x2924 x2923 x2922 x2921 x2920 x2919 x2918 x2917 x2916 x2915 x2914 x2913 x2912 x2911 x2910 x2909 x2908 x2907 x2906 x2905 x2904 x2903 x2902 x2901 x2900 x2899 x2898 x2897 x2896 x2895 x2894 x2893 x2892 x2891 x2890 x2889 x2888 x2887 x2886 x2885 x2884 x2883 x2882 x2881 x2880 x2879 x2878 x2877 x2876 x2875 x2874 x2873 x2872 x2871 x2870 x2869 x2868 x2867 x2866 x2865 x2864 x2863 x2862 x2861 x2860 x2859 x2858 x2857 x2856 x2855 x2854 x2853 x2852 x2851 x2850 x2849 x2848 x2847 x2846 x2845 x2844 x2843 x2842 x2841 x2840 x2839 x2838 x2837 x2836 x2835 x2834 x2833 x2832 x2831 x2830 x2829 x2828 x2827 x2826 x2825 x2824 x2823 x2822 x2821 x2820 x2819 x2818 x2817 x2816 x2815 x2814 x2813 x2812 x2811 x2810 x2809 x2808 x2807 x2806 x2805 x2804 x2803 x2802 x2801 x2800 x2799 x2798 x2797 x2796 x2795 x2794 x2793 x2792 x2791 x2790 x2789 x2788 x2787 x2786 x2785 x2784 x2783 x2782 x2781 x2780 x2779 x2778 x2777 x2776 x2775 x2774 x2773 x2772 x2771 x2770 x2769 x2768 x2767 x2766 x2765 x2764 x2763 x2762 x2761 x2760 x2759 x2758 x2757 x2756 x2755 x2754 x2753 x2752 x2751 x2750 x2749 x2748 x2747 x2746 x2745 x2744 x2743 x2742 x2741 x2740 x2739 x2738 x2737 x2736 x2735 x2734 x2733 x2732 x2731 x2730 x2729 x2728 x2727 x2726 x2725 x2724 x2723 x2722 x2721 x2720 x2719 x2718 x2717 x2716 x2715 x2714 x2713 x2712 x2711 x2710 x2709 x2708 x2707 x2706 x2705 x2704 x2703 x2702 x2701 x2700 x2699 x2698 x2697 x2696 x2695 x2694 x2693 x2692 x2691 x2690 x2689 x2688 x2687 x2686 x2685 x2684 x2683 x2682 x2681 x2680 x2679 x2678 x2677 x2676 x2675 x2674 x2673 x2672 x2671 x2670 x2669 x2668 x2667 x2666 x2665 x2664 x2663 x2662 x2661 x2660 x2659 x2658 x2657 x2656 x2655 x2654 x2653 x2652 x2651 x2650 x2649 x2648 x2647 x2646 x2645 x2644 x2643 x2642 x2641 x2640 x2639 x2638 x2637 x2636 x2635 x2634 x2633 x2632 x2631 x2630 x2629 x2628 x2627 x2626 x2625 x2624 x2623 x2622 x2621 x2620 x2619 x2618 x2617 x2616 x2615 x2614 x2613 x2612 x2611 x2610 x2609 x2608 x2607 x2606 x2605 x2604 x2603 x2602 x2601 x2600 x2599 x2598 x2597 x2596 x2595 x2594 x2593 x2592 x2591 x2590 x2589 x2588 x2587 x2586 x2585 x2584 x2583 x2582 x2581 x2580 x2579 x2578 x2577 x2576 x2575 x2574 x2573 x2572 x2571 x2570 x2569 x2568 x2567 x2566 x2565 x2564 x2563 x2562 x2561 x2560 x2559 x2558 x2557 x2556 x2555 x2554 x2553 x2552 x2551 x2550 x2549 x2548 x2547 x2546 x2545 x2544 x2543 x2542 x2541 x2540 x2539 x2538 x2537 x2536 x2535 x2534 x2533 x2532 x2531 x2530 x2529 x2528 x2527 x2526 x2525 x2524 x2523 x2522 x2521 x2520 x2519 x2518 x2517 x2516 x2515 x2514 x2513 x2512 x2511 x2510 x2509 x2508 x2507 x2506 x2505 x2504 x2503 x2502 x2501 x2500 x2499 x2498 x2497 x2496 x2495 x2494 x2493 x2492 x2491 x2490 x2489 x2488 x2487 x2486 x2485 x2484 x2483 x2482 x2481 x2480 x2479 x2478 x2477 x2476 x2475 x2474 x2473 x2472 x2471 x2470 x2469 x2468 x2467 x2466 x2465 x2464 x2463 x2462 x2461 x2460 x2459 x2458 x2457 x2456 x2455 x2454 x2453 x2452 x2451 x2450 x2449 x2448 x2447 x2446 x2445 x2444 x2443 x2442 x2441 x2440 x2439 x2438 x2437 x2436 x2435 x2434 x2433 x2432 x2431 x2430 x2429 x2428 x2427 x2426 x2425 x2424 x2423 x2422 x2421 x2420 x2419 x2418 x2417 x2416 x2415 x2414 x2413 x2412 x2411 x2410 x2409 x2408 x2407 x2406 x2405 x2404 x2403 x2402 x2401 x2400 x2399 x2398 x2397 x2396 x2395 x2394 x2393 x2392 x2391 x2390 x2389 x2388 x2387 x2386 x2385 x2384 x2383 x2382 x2381 x2380 x2379 x2378 x2377 x2376 x2375 x2374 x2373 x2372 x2371 x2370 x2369 x2368 x2367 x2366 x2365 x2364 x2363 x2362 x2361 x2360 x2359 x2358 x2357 x2356 x2355 x2354 x2353 x2352 x2351 x2350 x2349 x2348 x2347 x2346 x2345 x2344 x2343 x2342 x2341 x2340 x2339 x2338 x2337 x2336 x2335 x2334 x2333 x2332 x2331 x2330 x2329 x2328 x2327 x2326 x2325 x2324 x2323 x2322 x2321 x2320 x2319 x2318 x2317 x2316 x2315 x2314 x2313 x2312 x2311 x2310 x2309 x2308 x2307 x2306 x2305 x2304 x2303 x2302 x2301 x2300 x2299 x2298 x2297 x2296 x2295 x2294 x2293 x2292 x2291 x2290 x2289 x2288 x2287 x2286 x2285 x2284 x2283 x2282 x2281 x2280 x2279 x2278 x2277 x2276 x2275 x2274 x2273 x2272 x2271 x2270 x2269 x2268 x2267 x2266 x2265 x2264 x2263 x2262 x2261 x2260 x2259 x2258 x2257 x2256 x2255 x2254 x2253 x2252 x2251 x2250 x2249 x2248 x2247 x2246 x2245 x2244 x2243 x2242 x2241 x2240 x2239 x2238 x2237 x2236 x2235 x2234 x2233 x2232 x2231 x2230 x2229 x2228 x2227 x2226 x2225 x2224 x2223 x2222 x2221 x2220 x2219 x2218 x2217 x2216 x2215 x2214 x2213 x2212 x2211 x2210 x2209 x2208 x2207 x2206 x2205 x2204 x2203 x2202 x2201 x2200 x2199 x2198 x2197 x2196 x2195 x2194 x2193 x2192 x2191 x2190 x2189 x2188 x2187 x2186 x2185 x2184 x2183 x2182 x2181 x2180 x2179 x2178 x2177 x2176 x2175 x2174 x2173 x2172 x2171 x2170 x2169 x2168 x2167 x2166 x2165 x2164 x2163 x2162 x2161 x2160 x2159 x2158 x2157 x2156 x2155 x2154 x2153 x2152 x2151 x2150 x2149 x2148 x2147 x2146 x2145 x2144 x2143 x2142 x2141 x2140 x2139 x2138 x2137 x2136 x2135 x2134 x2133 x2132 x2131 x2130 x2129 x2128 x2127 x2126 x2125 x2124 x2123 x2122 x2121 x2120 x2119 x2118 x2117 x2116 x2115 x2114 x2113 x2112 x2111 x2110 x2109 x2108 x2107 x2106 x2105 x2104 x2103 x2102 x2101 x2100 x2099 x2098 x2097 x2096 x2095 x2094 x2093 x2092 x2091 x2090 x2089 x2088 x2087 x2086 x2085 x2084 x2083 x2082 x2081 x2080 x2079 x2078 x2077 x2076 x2075 x2074 x2073 x2072 x2071 x2070 x2069 x2068 x2067 x2066 x2065 x2064 x2063 x2062 x2061 x2060 x2059 x2058 x2057 x2056 x2055 x2054 x2053 x2052 x2051 x2050 x2049 x2048 x2047 x2046 x2045 x2044 x2043 x2042 x2041 x2040 x2039 x2038 x2037 x2036 x2035 x2034 x2033 x2032 x2031 x2030 x2029 x2028 x2027 x2026 x2025 x2024 x2023 x2022 x2021 x2020 x2019 x2018 x2017 x2016 x2015 x2014 x2013 x2012 x2011 x2010 x2009 x2008 x2007 x2006 x2005 x2004 x2003 x2002 x2001 x2000 x1999 x1998 x1997 x1996 x1995 x1994 x1993 x1992 x1991 x1990 x1989 x1988 x1987 x1986 x1985 x1984 x1983 x1982 x1981 x1980 x1979 x1978 x1977 x1976 x1975 x1974 x1973 x1972 x1971 x1970 x1969 x1968 x1967 x1966 x1965 x1964 x1963 x1962 x1961 x1960 x1959 x1958 x1957 x1956 x1955 x1954 x1953 x1952 x1951 x1950 x1949 x1948 x1947 x1946 x1945 x1944 x1943 x1942 x1941 x1940 x1939 x1938 x1937 x1936 x1935 x1934 x1933 x1932 x1931 x1930 x1929 x1928 x1927 x1926 x1925 x1924 x1923 x1922 x1921 x1920 x1919 x1918 x1917 x1916 x1915 x1914 x1913 x1912 x1911 x1910 x1909 x1908 x1907 x1906 x1905 x1904 x1903 x1902 x1901 x1900 x1899 x1898 x1897 x1896 x1895 x1894 x1893 x1892 x1891 x1890 x1889 x1888 x1887 x1886 x1885 x1884 x1883 x1882 x1881 x1880 x1879 x1878 x1877 x1876 x1875 x1874 x1873 x1872 x1871 x1870 x1869 x1868 x1867 x1866 x1865 x1864 x1863 x1862 x1861 x1860 x1859 x1858 x1857 x1856 x1855 x1854 x1853 x1852 x1851 x1850 x1849 x1848 x1847 x1846 x1845 x1844 x1843 x1842 x1841 x1840 x1839 x1838 x1837 x1836 x1835 x1834 x1833 x1832 x1831 x1830 x1829 x1828 x1827 x1826 x1825 x1824 x1823 x1822 x1821 x1820 x1819 x1818 x1817 x1816 x1815 x1814 x1813 x1812 x1811 x1810 x1809 x1808 x1807 x1806 x1805 x1804 x1803 x1802 x1801 x1800 x1799 x1798 x1797 x1796 x1795 x1794 x1793 x1792 x1791 x1790 x1789 x1788 x1787 x1786 x1785 x1784 x1783 x1782 x1781 x1780 x1779 x1778 x1777 x1776 x1775 x1774 x1773 x1772 x1771 x1770 x1769 x1768 x1767 x1766 x1765 x1764 x1763 x1762 x1761 x1760 x1759 x1758 x1757 x1756 x1755 x1754 x1753 x1752 x1751 x1750 x1749 x1748 x1747 x1746 x1745 x1744 x1743 x1742 x1741 x1740 x1739 x1738 x1737 x1736 x1735 x1734 x1733 x1732 x1731 x1730 x1729 x1728 x1727 x1726 x1725 x1724 x1723 x1722 x1721 x1720 x1719 x1718 x1717 x1716 x1715 x1714 x1713 x1712 x1711 x1710 x1709 x1708 x1707 x1706 x1705 x1704 x1703 x1702 x1701 x1700 x1699 x1698 x1697 x1696 x1695 x1694 x1693 x1692 x1691 x1690 x1689 x1688 x1687 x1686 x1685 x1684 x1683 x1682 x1681 x1680 x1679 x1678 x1677 x1676 x1675 x1674 x1673 x1672 x1671 x1670 x1669 x1668 x1667 x1666 x1665 x1664 x1663 x1662 x1661 x1660 x1659 x1658 x1657 x1656 x1655 x1654 x1653 x1652 x1651 x1650 x1649 x1648 x1647 x1646 x1645 x1644 x1643 x1642 x1641 x1640 x1639 x1638 x1637 x1636 x1635 x1634 x1633 x1632 x1631 x1630 x1629 x1628 x1627 x1626 x1625 x1624 x1623 x1622 x1621 x1620 x1619 x1618 x1617 x1616 x1615 x1614 x1613 x1612 x1611 x1610 x1609 x1608 x1607 x1606 x1605 x1604 x1603 x1602 x1601 x1600 x1599 x1598 x1597 x1596 x1595 x1594 x1593 x1592 x1591 x1590 x1589 x1588 x1587 x1586 x1585 x1584 x1583 x1582 x1581 x1580 x1579 x1578 x1577 x1576 x1575 x1574 x1573 x1572 x1571 x1570 x1569 x1568 x1567 x1566 x1565 x1564 x1563 x1562 x1561 x1560 x1559 x1558 x1557 x1556 x1555 x1554 x1553 x1552 x1551 x1550 x1549 x1548 x1547 x1546 x1545 x1544 x1543 x1542 x1541 x1540 x1539 x1538 x1537 x1536 x1535 x1534 x1533 x1532 x1531 x1530 x1529 x1528 x1527 x1526 x1525 x1524 x1523 x1522 x1521 x1520 x1519 x1518 x1517 x1516 x1515 x1514 x1513 x1512 x1511 x1510 x1509 x1508 x1507 x1506 x1505 x1504 x1503 x1502 x1501 x1500 x1499 x1498 x1497 x1496 x1495 x1494 x1493 x1492 x1491 x1490 x1489 x1488 x1487 x1486 x1485 x1484 x1483 x1482 x1481 x1480 x1479 x1478 x1477 x1476 x1475 x1474 x1473 x1472 x1471 x1470 x1469 x1468 x1467 x1466 x1465 x1464 x1463 x1462 x1461 x1460 x1459 x1458 x1457 x1456 x1455 x1454 x1453 x1452 x1451 x1450 x1449 x1448 x1447 x1446 x1445 x1444 x1443 x1442 x1441 x1440 x1439 x1438 x1437 x1436 x1435 x1434 x1433 x1432 x1431 x1430 x1429 x1428 x1427 x1426 x1425 x1424 x1423 x1422 x1421 x1420 x1419 x1418 x1417 x1416 x1415 x1414 x1413 x1412 x1411 x1410 x1409 x1408 x1407 x1406 x1405 x1404 x1403 x1402 x1401 x1400 x1399 x1398 x1397 x1396 x1395 x1394 x1393 x1392 x1391 x1390 x1389 x1388 x1387 x1386 x1385 x1384 x1383 x1382 x1381 x1380 x1379 x1378 x1377 x1376 x1375 x1374 x1373 x1372 x1371 x1370 x1369 x1368 x1367 x1366 x1365 x1364 x1363 x1362 x1361 x1360 x1359 x1358 x1357 x1356 x1355 x1354 x1353 x1352 x1351 x1350 x1349 x1348 x1347 x1346 x1345 x1344 x1343 x1342 x1341 x1340 x1339 x1338 x1337 x1336 x1335 x1334 x1333 x1332 x1331 x1330 x1329 x1328 x1327 x1326 x1325 x1324 x1323 x1322 x1321 x1320 x1319 x1318 x1317 x1316 x1315 x1314 x1313 x1312 x1311 x1310 x1309 x1308 x1307 x1306 x1305 x1304 x1303 x1302 x1301 x1300 x1299 x1298 x1297 x1296 x1295 x1294 x1293 x1292 x1291 x1290 x1289 x1288 x1287 x1286 x1285 x1284 x1283 x1282 x1281 x1280 x1279 x1278 x1277 x1276 x1275 x1274 x1273 x1272 x1271 x1270 x1269 x1268 x1267 x1266 x1265 x1264 x1263 x1262 x1261 x1260 x1259 x1258 x1257 x1256 x1255 x1254 x1253 x1252 x1251 x1250 x1249 x1248 x1247 x1246 x1245 x1244 x1243 x1242 x1241 x1240 x1239 x1238 x1237 x1236 x1235 x1234 x1233 x1232 x1231 x1230 x1229 x1228 x1227 x1226 x1225 x1224 x1223 x1222 x1221 x1220 x1219 x1218 x1217 x1216 x1215 x1214 x1213 x1212 x1211 x1210 x1209 x1208 x1207 x1206 x1205 x1204 x1203 x1202 x1201 x1200 x1199 x1198 x1197 x1196 x1195 x1194 x1193 x1192 x1191 x1190 x1189 x1188 x1187 x1186 x1185 x1184 x1183 x1182 x1181 x1180 x1179 x1178 x1177 x1176 x1175 x1174 x1173 x1172 x1171 x1170 x1169 x1168 x1167 x1166 x1165 x1164 x1163 x1162 x1161 x1160 x1159 x1158 x1157 x1156 x1155 x1154 x1153 x1152 x1151 x1150 x1149 x1148 x1147 x1146 x1145 x1144 x1143 x1142 x1141 x1140 x1139 x1138 x1137 x1136 x1135 x1134 x1133 x1132 x1131 x1130 x1129 x1128 x1127 x1126 x1125 x1124 x1123 x1122 x1121 x1120 x1119 x1118 x1117 x1116 x1115 x1114 x1113 x1112 x1111 x1110 x1109 x1108 x1107 x1106 x1105 x1104 x1103 x1102 x1101 x1100 x1099 x1098 x1097 x1096 x1095 x1094 x1093 x1092 x1091 x1090 x1089 x1088 x1087 x1086 x1085 x1084 x1083 x1082 x1081 x1080 x1079 x1078 x1077 x1076 x1075 x1074 x1073 x1072 x1071 x1070 x1069 x1068 x1067 x1066 x1065 x1064 x1063 x1062 x1061 x1060 x1059 x1058 x1057 x1056 x1055 x1054 x1053 x1052 x1051 x1050 x1049 x1048 x1047 x1046 x1045 x1044 x1043 x1042 x1041 x1040 x1039 x1038 x1037 x1036 x1035 x1034 x1033 x1032 x1031 x1030 x1029 x1028 x1027 x1026 x1025 x1024 x1023 x1022 x1021 x1020 x1019 x1018 x1017 x1016 x1015 x1014 x1013 x1012 x1011 x1010 x1009 x1008 x1007 x1006 x1005 x1004 x1003 x1002 x1001 x1000 x999 x998 x997 x996 x995 x994 x993 x992 x991 x990 x989 x988 x987 x986 x985 x984 x983 x982 x981 x980 x979 x978 x977 x976 x975 x974 x973 x972 x971 x970 x969 x968 x967 x966 x965 x964 x963 x962 x961 x960 x959 x958 x957 x956 x955 x954 x953 x952 x951 x950 x949 x948 x947 x946 x945 x944 x943 x942 x941 x940 x939 x938 x937 x936 x935 x934 x933 x932 x931 x930 x929 x928 x927 x926 x925 x924 x923 x922 x921 x920 x919 x918 x917 x916 x915 x914 x913 x912 x911 x910 x909 x908 x907 x906 x905 x904 x903 x902 x901 x900 x899 x898 x897 x896 x895 x894 x893 x892 x891 x890 x889 x888 x887 x886 x885 x884 x883 x882 x881 x880 x879 x878 x877 x876 x875 x874 x873 x872 x871 x870 x869 x868 x867 x866 x865 x864 x863 x862 x861 x860 x859 x858 x857 x856 x855 x854 x853 x852 x851 x850 x849 x848 x847 x846 x845 x844 x843 x842 x841 x840 x839 x838 x837 x836 x835 x834 x833 x832 x831 x830 x829 x828 x827 x826 x825 x824 x823 x822 x821 x820 x819 x818 x817 x816 x815 x814 x813 x812 x811 x810 x809 x808 x807 x806 x805 x804 x803 x802 x801 x800 x799 x798 x797 x796 x795 x794 x793 x792 x791 x790 x789 x788 x787 x786 x785 x784 x783 x782 x781 x780 x779 x778 x777 x776 x775 x774 x773 x772 x771 x770 x769 x768 x767 x766 x765 x764 x763 x762 x761 x760 x759 x758 x757 x756 x755 x754 x753 x752 x751 x750 x749 x748 x747 x746 x745 x744 x743 x742 x741 x740 x739 x738 x737 x736 x735 x734 x733 x732 x731 x730 x729 x728 x727 x726 x725 x724 x723 x722 x721 x720 x719 x718 x717 x716 x715 x714 x713 x712 x711 x710 x709 x708 x707 x706 x705 x704 x703 x702 x701 x700 x699 x698 x697 x696 x695 x694 x693 x692 x691 x690 x689 x688 x687 x686 x685 x684 x683 x682 x681 x680 x679 x678 x677 x676 x675 x674 x673 x672 x671 x670 x669 x668 x667 x666 x665 x664 x663 x662 x661 x660 x659 x658 x657 x656 x655 x654 x653 x652 x651 x650 x649 x648 x647 x646 x645 x644 x643 x642 x641 x640 x639 x638 x637 x636 x635 x634 x633 x632 x631 x630 x629 x628 x627 x626 x625 x624 x623 x622 x621 x620 x619 x618 x617 x616 x615 x614 x613 x612 x611 x610 x609 x608 x607 x606 x605 x604 x603 x602 x601 x600 x599 x598 x597 x596 x595 x594 x593 x592 x591 x590 x589 x588 x587 x586 x585 x584 x583 x582 x581 x580 x579 x578 x577 x576 x575 x574 x573 x572 x571 x570 x569 x568 x567 x566 x565 x564 x563 x562 x561 x560 x559 x558 x557 x556 x555 x554 x553 x552 x551 x550 x549 x548 x547 x546 x545 x544 x543 x542 x541 x540 x539 x538 x537 x536 x535 x534 x533 x532 x531 x530 x529 x528 x527 x526 x525 x524 x523 x522 x521 x520 x519 x518 x517 x516 x515 x514 x513 x512 x511 x510 x509 x508 x507 x506 x505 x504 x503 x502 x501 x500 x499 x498 x497 x496 x495 x494 x493 x492 x491 x490 x489 x488 x487 x486 x485 x484 x483 x482 x481 x480 x479 x478 x477 x476 x475 x474 x473 x472 x471 x470 x469 x468 x467 x466 x465 x464 x463 x462 x461 x460 x459 x458 x457 x456 x455 x454 x453 x452 x451 x450 x449 x448 x447 x446 x445 x444 x443 x442 x441 x440 x439 x438 x437 x436 x435 x434 x433 x432 x431 x430 x429 x428 x427 x426 x425 x424 x423 x422 x421 x420 x419 x418 x417 x416 x415 x414 x413 x412 x411 x410 x409 x408 x407 x406 x405 x404 x403 x402 x401 x400 x399 x398 x397 x396 x395 x394 x393 x392 x391 x390 x389 x388 x387 x386 x385 x384 x383 x382 x381 x380 x379 x378 x377 x376 x375 x374 x373 x372 x371 x370 x369 x368 x367 x366 x365 x364 x363 x362 x361 x360 x359 x358 x357 x356 x355 x354 x353 x352 x351 x350 x349 x348 x347 x346 x345 x344 x343 x342 x341 x340 x339 x338 x337 x336 x335 x334 x333 x332 x331 x330 x329 x328 x327 x326 x325 x324 x323 x322 x321 x320 x319 x318 x317 x316 x315 x314 x313 x312 x311 x310 x309 x308 x307 x306 x305 x304 x303 x302 x301 x300 x299 x298 x297 x296 x295 x294 x293 x292 x291 x290 x289 x288 x287 x286 x285 x284 x283 x282 x281 x280 x279 x278 x277 x276 x275 x274 x273 x272 x271 x270 x269 x268 x267 x266 x265 x264 x263 x262 x261 x260 x259 x258 x257 x256 x255 x254 x253 x252 x251 x250 x249 x248 x247 x246 x245 x244 x243 x242 x241 x240 x239 x238 x237 x236 x235 x234 x233 x232 x231 x230 x229 x228 x227 x226 x225 x224 x223 x222 x221 x220 x219 x218 x217 x216 x215 x214 x213 x212 x211 x210 x209 x208 x207 x206 x205 x204 x203 x202 x201 x200 x199 x198 x197 x196 x195 x194 x193 x192 x191 x190 x189 x188 x187 x186 x185 x184 x183 x182 x181 x180 x179 x178 x177 x176 x175 x174 x173 x172 x171 x170 x169 x168 x167 x166 x165 x164 x163 x162 x161 x160 x159 x158 x157 x156 x155 x154 x153 x152 x151 x150 x149 x148 x147 x146 x145 x144 x143 x142 x141 x140 x139 x138 x137 x136 x135 x134 x133 x132 x131 x130 x129 x128 x127 x126 x125 x124 x123 x122 x121 x120 x119 x118 x117 x116 x115 x114 x113 x112 x111 x110 x109 x108 x107 x106 x105 x104 x103 x102 x101 x100 x99 x98 x97 x96 x95 x94 x93 x92 x91 x90 x89 x88 x87 x86 x85 x84 x83 x82 x81 x80 x79 x78 x77 x76 x75 x74 x73 x72 x71 x70 x69 x68 x67 x66 x65 x64 x63 x62 x61 x60 x59 x58 x57 x56 x55 x54 x53 x52 x51 x50 x49 x48 x47 x46 x45 x44 x43 x42 x41 x40 x39 x38 x37 x36 x35 x34 x33 x32 x31 x30 x29 x28 x27 x26 x25 x24 x23 x22 x21 x20 x19 x18 x17 x16 x15 x14 x13 x12 x11 x10 x9 x8 x7 x6 x5 x4 x3 x2 x1 x0 | y0 (DUT) y_ref (Maj5025)");
    $display("---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------");
    // Loop through all 4739452898216418547201653797763595860957428722528977235532895354610283334595157992601954763893350737531098159036292099891217849718658132949599338305423909899252433568409523604296927531388595995903212328377859293925028196664665449850920047372460929548959622342553774931470029996136721692487549847800783165669065600283216761882728648823088672849767761096787054409317648768673870046197091729852874525071048417569058029910574146116161366297222991158549940296605431801079820504387040532005678479769096620906801991999931319916541911339092108224127155815316085299843959201857069250074266999672661907812994957711857222227385566463837903557701706172013317028659878977488721010157415572005239921821872642128383718566810743592190387800338965309406435642999976013852377063915568381663822154853706240880713672399028318733383264792633014849194780378227897156978938757328083522020917300464403999534043883489380242875421456525648278512104832460583690257724803208284252160095154337085117492746715082940721986813303177842688134816866983859627735702246922741856296160056654162807679644176131822175861244568214031779577836287324457834556298882134763531751909360525557572719095658843766275014763096181817096664181823043722510021319610830579781988247221574674180784741135629303528577581367198572085824120663747784090886290823216458725893664233566807777314155339529598238740914418234871716424282967739043062987444191457487347008423479118751929185205742311071535373987016939985312505575666322649798388484889607881003797682733554107154432 combinations
    for (idx = 0; idx < TOTAL_VECTORS; idx = idx + 1) begin
      x = idx[5024:0];
      #10 $display("%4t |  %b  |   %b       %b",
                   $time, x, y0, y_ref);
    end
    #10 $finish;
  end

  // Optional mismatch check
  always #1 if (^x !== 1'bx && y0 !== y_ref)
    $display("Mismatch at t=%0t x=%b HW=%0d y0=%0b ref=%0b",
             $time, x, popcount(x), y0, y_ref);

endmodule

`default_nettype wire
