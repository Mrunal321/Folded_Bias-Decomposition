`timescale 1ns/1ps
`default_nettype none

module tb_top;
  // 3001-bit input vector
  reg  [3000:0] x = 3001'b0;
  wire       y0;
  reg  [63:0] idx;

  // DUT instantiation
  top dut (
    .x0(x[0]), .x1(x[1]), .x2(x[2]), .x3(x[3]), .x4(x[4]), .x5(x[5]), .x6(x[6]), .x7(x[7]), .x8(x[8]), .x9(x[9]), .x10(x[10]), .x11(x[11]), .x12(x[12]), .x13(x[13]), .x14(x[14]), .x15(x[15]), .x16(x[16]), .x17(x[17]), .x18(x[18]), .x19(x[19]), .x20(x[20]), .x21(x[21]), .x22(x[22]), .x23(x[23]), .x24(x[24]), .x25(x[25]), .x26(x[26]), .x27(x[27]), .x28(x[28]), .x29(x[29]), .x30(x[30]), .x31(x[31]), .x32(x[32]), .x33(x[33]), .x34(x[34]), .x35(x[35]), .x36(x[36]), .x37(x[37]), .x38(x[38]), .x39(x[39]), .x40(x[40]), .x41(x[41]), .x42(x[42]), .x43(x[43]), .x44(x[44]), .x45(x[45]), .x46(x[46]), .x47(x[47]), .x48(x[48]), .x49(x[49]), .x50(x[50]), .x51(x[51]), .x52(x[52]), .x53(x[53]), .x54(x[54]), .x55(x[55]), .x56(x[56]), .x57(x[57]), .x58(x[58]), .x59(x[59]), .x60(x[60]), .x61(x[61]), .x62(x[62]), .x63(x[63]), .x64(x[64]), .x65(x[65]), .x66(x[66]), .x67(x[67]), .x68(x[68]), .x69(x[69]), .x70(x[70]), .x71(x[71]), .x72(x[72]), .x73(x[73]), .x74(x[74]), .x75(x[75]), .x76(x[76]), .x77(x[77]), .x78(x[78]), .x79(x[79]), .x80(x[80]), .x81(x[81]), .x82(x[82]), .x83(x[83]), .x84(x[84]), .x85(x[85]), .x86(x[86]), .x87(x[87]), .x88(x[88]), .x89(x[89]), .x90(x[90]), .x91(x[91]), .x92(x[92]), .x93(x[93]), .x94(x[94]), .x95(x[95]), .x96(x[96]), .x97(x[97]), .x98(x[98]), .x99(x[99]), .x100(x[100]), .x101(x[101]), .x102(x[102]), .x103(x[103]), .x104(x[104]), .x105(x[105]), .x106(x[106]), .x107(x[107]), .x108(x[108]), .x109(x[109]), .x110(x[110]), .x111(x[111]), .x112(x[112]), .x113(x[113]), .x114(x[114]), .x115(x[115]), .x116(x[116]), .x117(x[117]), .x118(x[118]), .x119(x[119]), .x120(x[120]), .x121(x[121]), .x122(x[122]), .x123(x[123]), .x124(x[124]), .x125(x[125]), .x126(x[126]), .x127(x[127]), .x128(x[128]), .x129(x[129]), .x130(x[130]), .x131(x[131]), .x132(x[132]), .x133(x[133]), .x134(x[134]), .x135(x[135]), .x136(x[136]), .x137(x[137]), .x138(x[138]), .x139(x[139]), .x140(x[140]), .x141(x[141]), .x142(x[142]), .x143(x[143]), .x144(x[144]), .x145(x[145]), .x146(x[146]), .x147(x[147]), .x148(x[148]), .x149(x[149]), .x150(x[150]), .x151(x[151]), .x152(x[152]), .x153(x[153]), .x154(x[154]), .x155(x[155]), .x156(x[156]), .x157(x[157]), .x158(x[158]), .x159(x[159]), .x160(x[160]), .x161(x[161]), .x162(x[162]), .x163(x[163]), .x164(x[164]), .x165(x[165]), .x166(x[166]), .x167(x[167]), .x168(x[168]), .x169(x[169]), .x170(x[170]), .x171(x[171]), .x172(x[172]), .x173(x[173]), .x174(x[174]), .x175(x[175]), .x176(x[176]), .x177(x[177]), .x178(x[178]), .x179(x[179]), .x180(x[180]), .x181(x[181]), .x182(x[182]), .x183(x[183]), .x184(x[184]), .x185(x[185]), .x186(x[186]), .x187(x[187]), .x188(x[188]), .x189(x[189]), .x190(x[190]), .x191(x[191]), .x192(x[192]), .x193(x[193]), .x194(x[194]), .x195(x[195]), .x196(x[196]), .x197(x[197]), .x198(x[198]), .x199(x[199]), .x200(x[200]), .x201(x[201]), .x202(x[202]), .x203(x[203]), .x204(x[204]), .x205(x[205]), .x206(x[206]), .x207(x[207]), .x208(x[208]), .x209(x[209]), .x210(x[210]), .x211(x[211]), .x212(x[212]), .x213(x[213]), .x214(x[214]), .x215(x[215]), .x216(x[216]), .x217(x[217]), .x218(x[218]), .x219(x[219]), .x220(x[220]), .x221(x[221]), .x222(x[222]), .x223(x[223]), .x224(x[224]), .x225(x[225]), .x226(x[226]), .x227(x[227]), .x228(x[228]), .x229(x[229]), .x230(x[230]), .x231(x[231]), .x232(x[232]), .x233(x[233]), .x234(x[234]), .x235(x[235]), .x236(x[236]), .x237(x[237]), .x238(x[238]), .x239(x[239]), .x240(x[240]), .x241(x[241]), .x242(x[242]), .x243(x[243]), .x244(x[244]), .x245(x[245]), .x246(x[246]), .x247(x[247]), .x248(x[248]), .x249(x[249]), .x250(x[250]), .x251(x[251]), .x252(x[252]), .x253(x[253]), .x254(x[254]), .x255(x[255]), .x256(x[256]), .x257(x[257]), .x258(x[258]), .x259(x[259]), .x260(x[260]), .x261(x[261]), .x262(x[262]), .x263(x[263]), .x264(x[264]), .x265(x[265]), .x266(x[266]), .x267(x[267]), .x268(x[268]), .x269(x[269]), .x270(x[270]), .x271(x[271]), .x272(x[272]), .x273(x[273]), .x274(x[274]), .x275(x[275]), .x276(x[276]), .x277(x[277]), .x278(x[278]), .x279(x[279]), .x280(x[280]), .x281(x[281]), .x282(x[282]), .x283(x[283]), .x284(x[284]), .x285(x[285]), .x286(x[286]), .x287(x[287]), .x288(x[288]), .x289(x[289]), .x290(x[290]), .x291(x[291]), .x292(x[292]), .x293(x[293]), .x294(x[294]), .x295(x[295]), .x296(x[296]), .x297(x[297]), .x298(x[298]), .x299(x[299]), .x300(x[300]), .x301(x[301]), .x302(x[302]), .x303(x[303]), .x304(x[304]), .x305(x[305]), .x306(x[306]), .x307(x[307]), .x308(x[308]), .x309(x[309]), .x310(x[310]), .x311(x[311]), .x312(x[312]), .x313(x[313]), .x314(x[314]), .x315(x[315]), .x316(x[316]), .x317(x[317]), .x318(x[318]), .x319(x[319]), .x320(x[320]), .x321(x[321]), .x322(x[322]), .x323(x[323]), .x324(x[324]), .x325(x[325]), .x326(x[326]), .x327(x[327]), .x328(x[328]), .x329(x[329]), .x330(x[330]), .x331(x[331]), .x332(x[332]), .x333(x[333]), .x334(x[334]), .x335(x[335]), .x336(x[336]), .x337(x[337]), .x338(x[338]), .x339(x[339]), .x340(x[340]), .x341(x[341]), .x342(x[342]), .x343(x[343]), .x344(x[344]), .x345(x[345]), .x346(x[346]), .x347(x[347]), .x348(x[348]), .x349(x[349]), .x350(x[350]), .x351(x[351]), .x352(x[352]), .x353(x[353]), .x354(x[354]), .x355(x[355]), .x356(x[356]), .x357(x[357]), .x358(x[358]), .x359(x[359]), .x360(x[360]), .x361(x[361]), .x362(x[362]), .x363(x[363]), .x364(x[364]), .x365(x[365]), .x366(x[366]), .x367(x[367]), .x368(x[368]), .x369(x[369]), .x370(x[370]), .x371(x[371]), .x372(x[372]), .x373(x[373]), .x374(x[374]), .x375(x[375]), .x376(x[376]), .x377(x[377]), .x378(x[378]), .x379(x[379]), .x380(x[380]), .x381(x[381]), .x382(x[382]), .x383(x[383]), .x384(x[384]), .x385(x[385]), .x386(x[386]), .x387(x[387]), .x388(x[388]), .x389(x[389]), .x390(x[390]), .x391(x[391]), .x392(x[392]), .x393(x[393]), .x394(x[394]), .x395(x[395]), .x396(x[396]), .x397(x[397]), .x398(x[398]), .x399(x[399]), .x400(x[400]), .x401(x[401]), .x402(x[402]), .x403(x[403]), .x404(x[404]), .x405(x[405]), .x406(x[406]), .x407(x[407]), .x408(x[408]), .x409(x[409]), .x410(x[410]), .x411(x[411]), .x412(x[412]), .x413(x[413]), .x414(x[414]), .x415(x[415]), .x416(x[416]), .x417(x[417]), .x418(x[418]), .x419(x[419]), .x420(x[420]), .x421(x[421]), .x422(x[422]), .x423(x[423]), .x424(x[424]), .x425(x[425]), .x426(x[426]), .x427(x[427]), .x428(x[428]), .x429(x[429]), .x430(x[430]), .x431(x[431]), .x432(x[432]), .x433(x[433]), .x434(x[434]), .x435(x[435]), .x436(x[436]), .x437(x[437]), .x438(x[438]), .x439(x[439]), .x440(x[440]), .x441(x[441]), .x442(x[442]), .x443(x[443]), .x444(x[444]), .x445(x[445]), .x446(x[446]), .x447(x[447]), .x448(x[448]), .x449(x[449]), .x450(x[450]), .x451(x[451]), .x452(x[452]), .x453(x[453]), .x454(x[454]), .x455(x[455]), .x456(x[456]), .x457(x[457]), .x458(x[458]), .x459(x[459]), .x460(x[460]), .x461(x[461]), .x462(x[462]), .x463(x[463]), .x464(x[464]), .x465(x[465]), .x466(x[466]), .x467(x[467]), .x468(x[468]), .x469(x[469]), .x470(x[470]), .x471(x[471]), .x472(x[472]), .x473(x[473]), .x474(x[474]), .x475(x[475]), .x476(x[476]), .x477(x[477]), .x478(x[478]), .x479(x[479]), .x480(x[480]), .x481(x[481]), .x482(x[482]), .x483(x[483]), .x484(x[484]), .x485(x[485]), .x486(x[486]), .x487(x[487]), .x488(x[488]), .x489(x[489]), .x490(x[490]), .x491(x[491]), .x492(x[492]), .x493(x[493]), .x494(x[494]), .x495(x[495]), .x496(x[496]), .x497(x[497]), .x498(x[498]), .x499(x[499]), .x500(x[500]), .x501(x[501]), .x502(x[502]), .x503(x[503]), .x504(x[504]), .x505(x[505]), .x506(x[506]), .x507(x[507]), .x508(x[508]), .x509(x[509]), .x510(x[510]), .x511(x[511]), .x512(x[512]), .x513(x[513]), .x514(x[514]), .x515(x[515]), .x516(x[516]), .x517(x[517]), .x518(x[518]), .x519(x[519]), .x520(x[520]), .x521(x[521]), .x522(x[522]), .x523(x[523]), .x524(x[524]), .x525(x[525]), .x526(x[526]), .x527(x[527]), .x528(x[528]), .x529(x[529]), .x530(x[530]), .x531(x[531]), .x532(x[532]), .x533(x[533]), .x534(x[534]), .x535(x[535]), .x536(x[536]), .x537(x[537]), .x538(x[538]), .x539(x[539]), .x540(x[540]), .x541(x[541]), .x542(x[542]), .x543(x[543]), .x544(x[544]), .x545(x[545]), .x546(x[546]), .x547(x[547]), .x548(x[548]), .x549(x[549]), .x550(x[550]), .x551(x[551]), .x552(x[552]), .x553(x[553]), .x554(x[554]), .x555(x[555]), .x556(x[556]), .x557(x[557]), .x558(x[558]), .x559(x[559]), .x560(x[560]), .x561(x[561]), .x562(x[562]), .x563(x[563]), .x564(x[564]), .x565(x[565]), .x566(x[566]), .x567(x[567]), .x568(x[568]), .x569(x[569]), .x570(x[570]), .x571(x[571]), .x572(x[572]), .x573(x[573]), .x574(x[574]), .x575(x[575]), .x576(x[576]), .x577(x[577]), .x578(x[578]), .x579(x[579]), .x580(x[580]), .x581(x[581]), .x582(x[582]), .x583(x[583]), .x584(x[584]), .x585(x[585]), .x586(x[586]), .x587(x[587]), .x588(x[588]), .x589(x[589]), .x590(x[590]), .x591(x[591]), .x592(x[592]), .x593(x[593]), .x594(x[594]), .x595(x[595]), .x596(x[596]), .x597(x[597]), .x598(x[598]), .x599(x[599]), .x600(x[600]), .x601(x[601]), .x602(x[602]), .x603(x[603]), .x604(x[604]), .x605(x[605]), .x606(x[606]), .x607(x[607]), .x608(x[608]), .x609(x[609]), .x610(x[610]), .x611(x[611]), .x612(x[612]), .x613(x[613]), .x614(x[614]), .x615(x[615]), .x616(x[616]), .x617(x[617]), .x618(x[618]), .x619(x[619]), .x620(x[620]), .x621(x[621]), .x622(x[622]), .x623(x[623]), .x624(x[624]), .x625(x[625]), .x626(x[626]), .x627(x[627]), .x628(x[628]), .x629(x[629]), .x630(x[630]), .x631(x[631]), .x632(x[632]), .x633(x[633]), .x634(x[634]), .x635(x[635]), .x636(x[636]), .x637(x[637]), .x638(x[638]), .x639(x[639]), .x640(x[640]), .x641(x[641]), .x642(x[642]), .x643(x[643]), .x644(x[644]), .x645(x[645]), .x646(x[646]), .x647(x[647]), .x648(x[648]), .x649(x[649]), .x650(x[650]), .x651(x[651]), .x652(x[652]), .x653(x[653]), .x654(x[654]), .x655(x[655]), .x656(x[656]), .x657(x[657]), .x658(x[658]), .x659(x[659]), .x660(x[660]), .x661(x[661]), .x662(x[662]), .x663(x[663]), .x664(x[664]), .x665(x[665]), .x666(x[666]), .x667(x[667]), .x668(x[668]), .x669(x[669]), .x670(x[670]), .x671(x[671]), .x672(x[672]), .x673(x[673]), .x674(x[674]), .x675(x[675]), .x676(x[676]), .x677(x[677]), .x678(x[678]), .x679(x[679]), .x680(x[680]), .x681(x[681]), .x682(x[682]), .x683(x[683]), .x684(x[684]), .x685(x[685]), .x686(x[686]), .x687(x[687]), .x688(x[688]), .x689(x[689]), .x690(x[690]), .x691(x[691]), .x692(x[692]), .x693(x[693]), .x694(x[694]), .x695(x[695]), .x696(x[696]), .x697(x[697]), .x698(x[698]), .x699(x[699]), .x700(x[700]), .x701(x[701]), .x702(x[702]), .x703(x[703]), .x704(x[704]), .x705(x[705]), .x706(x[706]), .x707(x[707]), .x708(x[708]), .x709(x[709]), .x710(x[710]), .x711(x[711]), .x712(x[712]), .x713(x[713]), .x714(x[714]), .x715(x[715]), .x716(x[716]), .x717(x[717]), .x718(x[718]), .x719(x[719]), .x720(x[720]), .x721(x[721]), .x722(x[722]), .x723(x[723]), .x724(x[724]), .x725(x[725]), .x726(x[726]), .x727(x[727]), .x728(x[728]), .x729(x[729]), .x730(x[730]), .x731(x[731]), .x732(x[732]), .x733(x[733]), .x734(x[734]), .x735(x[735]), .x736(x[736]), .x737(x[737]), .x738(x[738]), .x739(x[739]), .x740(x[740]), .x741(x[741]), .x742(x[742]), .x743(x[743]), .x744(x[744]), .x745(x[745]), .x746(x[746]), .x747(x[747]), .x748(x[748]), .x749(x[749]), .x750(x[750]), .x751(x[751]), .x752(x[752]), .x753(x[753]), .x754(x[754]), .x755(x[755]), .x756(x[756]), .x757(x[757]), .x758(x[758]), .x759(x[759]), .x760(x[760]), .x761(x[761]), .x762(x[762]), .x763(x[763]), .x764(x[764]), .x765(x[765]), .x766(x[766]), .x767(x[767]), .x768(x[768]), .x769(x[769]), .x770(x[770]), .x771(x[771]), .x772(x[772]), .x773(x[773]), .x774(x[774]), .x775(x[775]), .x776(x[776]), .x777(x[777]), .x778(x[778]), .x779(x[779]), .x780(x[780]), .x781(x[781]), .x782(x[782]), .x783(x[783]), .x784(x[784]), .x785(x[785]), .x786(x[786]), .x787(x[787]), .x788(x[788]), .x789(x[789]), .x790(x[790]), .x791(x[791]), .x792(x[792]), .x793(x[793]), .x794(x[794]), .x795(x[795]), .x796(x[796]), .x797(x[797]), .x798(x[798]), .x799(x[799]), .x800(x[800]), .x801(x[801]), .x802(x[802]), .x803(x[803]), .x804(x[804]), .x805(x[805]), .x806(x[806]), .x807(x[807]), .x808(x[808]), .x809(x[809]), .x810(x[810]), .x811(x[811]), .x812(x[812]), .x813(x[813]), .x814(x[814]), .x815(x[815]), .x816(x[816]), .x817(x[817]), .x818(x[818]), .x819(x[819]), .x820(x[820]), .x821(x[821]), .x822(x[822]), .x823(x[823]), .x824(x[824]), .x825(x[825]), .x826(x[826]), .x827(x[827]), .x828(x[828]), .x829(x[829]), .x830(x[830]), .x831(x[831]), .x832(x[832]), .x833(x[833]), .x834(x[834]), .x835(x[835]), .x836(x[836]), .x837(x[837]), .x838(x[838]), .x839(x[839]), .x840(x[840]), .x841(x[841]), .x842(x[842]), .x843(x[843]), .x844(x[844]), .x845(x[845]), .x846(x[846]), .x847(x[847]), .x848(x[848]), .x849(x[849]), .x850(x[850]), .x851(x[851]), .x852(x[852]), .x853(x[853]), .x854(x[854]), .x855(x[855]), .x856(x[856]), .x857(x[857]), .x858(x[858]), .x859(x[859]), .x860(x[860]), .x861(x[861]), .x862(x[862]), .x863(x[863]), .x864(x[864]), .x865(x[865]), .x866(x[866]), .x867(x[867]), .x868(x[868]), .x869(x[869]), .x870(x[870]), .x871(x[871]), .x872(x[872]), .x873(x[873]), .x874(x[874]), .x875(x[875]), .x876(x[876]), .x877(x[877]), .x878(x[878]), .x879(x[879]), .x880(x[880]), .x881(x[881]), .x882(x[882]), .x883(x[883]), .x884(x[884]), .x885(x[885]), .x886(x[886]), .x887(x[887]), .x888(x[888]), .x889(x[889]), .x890(x[890]), .x891(x[891]), .x892(x[892]), .x893(x[893]), .x894(x[894]), .x895(x[895]), .x896(x[896]), .x897(x[897]), .x898(x[898]), .x899(x[899]), .x900(x[900]), .x901(x[901]), .x902(x[902]), .x903(x[903]), .x904(x[904]), .x905(x[905]), .x906(x[906]), .x907(x[907]), .x908(x[908]), .x909(x[909]), .x910(x[910]), .x911(x[911]), .x912(x[912]), .x913(x[913]), .x914(x[914]), .x915(x[915]), .x916(x[916]), .x917(x[917]), .x918(x[918]), .x919(x[919]), .x920(x[920]), .x921(x[921]), .x922(x[922]), .x923(x[923]), .x924(x[924]), .x925(x[925]), .x926(x[926]), .x927(x[927]), .x928(x[928]), .x929(x[929]), .x930(x[930]), .x931(x[931]), .x932(x[932]), .x933(x[933]), .x934(x[934]), .x935(x[935]), .x936(x[936]), .x937(x[937]), .x938(x[938]), .x939(x[939]), .x940(x[940]), .x941(x[941]), .x942(x[942]), .x943(x[943]), .x944(x[944]), .x945(x[945]), .x946(x[946]), .x947(x[947]), .x948(x[948]), .x949(x[949]), .x950(x[950]), .x951(x[951]), .x952(x[952]), .x953(x[953]), .x954(x[954]), .x955(x[955]), .x956(x[956]), .x957(x[957]), .x958(x[958]), .x959(x[959]), .x960(x[960]), .x961(x[961]), .x962(x[962]), .x963(x[963]), .x964(x[964]), .x965(x[965]), .x966(x[966]), .x967(x[967]), .x968(x[968]), .x969(x[969]), .x970(x[970]), .x971(x[971]), .x972(x[972]), .x973(x[973]), .x974(x[974]), .x975(x[975]), .x976(x[976]), .x977(x[977]), .x978(x[978]), .x979(x[979]), .x980(x[980]), .x981(x[981]), .x982(x[982]), .x983(x[983]), .x984(x[984]), .x985(x[985]), .x986(x[986]), .x987(x[987]), .x988(x[988]), .x989(x[989]), .x990(x[990]), .x991(x[991]), .x992(x[992]), .x993(x[993]), .x994(x[994]), .x995(x[995]), .x996(x[996]), .x997(x[997]), .x998(x[998]), .x999(x[999]), .x1000(x[1000]), .x1001(x[1001]), .x1002(x[1002]), .x1003(x[1003]), .x1004(x[1004]), .x1005(x[1005]), .x1006(x[1006]), .x1007(x[1007]), .x1008(x[1008]), .x1009(x[1009]), .x1010(x[1010]), .x1011(x[1011]), .x1012(x[1012]), .x1013(x[1013]), .x1014(x[1014]), .x1015(x[1015]), .x1016(x[1016]), .x1017(x[1017]), .x1018(x[1018]), .x1019(x[1019]), .x1020(x[1020]), .x1021(x[1021]), .x1022(x[1022]), .x1023(x[1023]), .x1024(x[1024]), .x1025(x[1025]), .x1026(x[1026]), .x1027(x[1027]), .x1028(x[1028]), .x1029(x[1029]), .x1030(x[1030]), .x1031(x[1031]), .x1032(x[1032]), .x1033(x[1033]), .x1034(x[1034]), .x1035(x[1035]), .x1036(x[1036]), .x1037(x[1037]), .x1038(x[1038]), .x1039(x[1039]), .x1040(x[1040]), .x1041(x[1041]), .x1042(x[1042]), .x1043(x[1043]), .x1044(x[1044]), .x1045(x[1045]), .x1046(x[1046]), .x1047(x[1047]), .x1048(x[1048]), .x1049(x[1049]), .x1050(x[1050]), .x1051(x[1051]), .x1052(x[1052]), .x1053(x[1053]), .x1054(x[1054]), .x1055(x[1055]), .x1056(x[1056]), .x1057(x[1057]), .x1058(x[1058]), .x1059(x[1059]), .x1060(x[1060]), .x1061(x[1061]), .x1062(x[1062]), .x1063(x[1063]), .x1064(x[1064]), .x1065(x[1065]), .x1066(x[1066]), .x1067(x[1067]), .x1068(x[1068]), .x1069(x[1069]), .x1070(x[1070]), .x1071(x[1071]), .x1072(x[1072]), .x1073(x[1073]), .x1074(x[1074]), .x1075(x[1075]), .x1076(x[1076]), .x1077(x[1077]), .x1078(x[1078]), .x1079(x[1079]), .x1080(x[1080]), .x1081(x[1081]), .x1082(x[1082]), .x1083(x[1083]), .x1084(x[1084]), .x1085(x[1085]), .x1086(x[1086]), .x1087(x[1087]), .x1088(x[1088]), .x1089(x[1089]), .x1090(x[1090]), .x1091(x[1091]), .x1092(x[1092]), .x1093(x[1093]), .x1094(x[1094]), .x1095(x[1095]), .x1096(x[1096]), .x1097(x[1097]), .x1098(x[1098]), .x1099(x[1099]), .x1100(x[1100]), .x1101(x[1101]), .x1102(x[1102]), .x1103(x[1103]), .x1104(x[1104]), .x1105(x[1105]), .x1106(x[1106]), .x1107(x[1107]), .x1108(x[1108]), .x1109(x[1109]), .x1110(x[1110]), .x1111(x[1111]), .x1112(x[1112]), .x1113(x[1113]), .x1114(x[1114]), .x1115(x[1115]), .x1116(x[1116]), .x1117(x[1117]), .x1118(x[1118]), .x1119(x[1119]), .x1120(x[1120]), .x1121(x[1121]), .x1122(x[1122]), .x1123(x[1123]), .x1124(x[1124]), .x1125(x[1125]), .x1126(x[1126]), .x1127(x[1127]), .x1128(x[1128]), .x1129(x[1129]), .x1130(x[1130]), .x1131(x[1131]), .x1132(x[1132]), .x1133(x[1133]), .x1134(x[1134]), .x1135(x[1135]), .x1136(x[1136]), .x1137(x[1137]), .x1138(x[1138]), .x1139(x[1139]), .x1140(x[1140]), .x1141(x[1141]), .x1142(x[1142]), .x1143(x[1143]), .x1144(x[1144]), .x1145(x[1145]), .x1146(x[1146]), .x1147(x[1147]), .x1148(x[1148]), .x1149(x[1149]), .x1150(x[1150]), .x1151(x[1151]), .x1152(x[1152]), .x1153(x[1153]), .x1154(x[1154]), .x1155(x[1155]), .x1156(x[1156]), .x1157(x[1157]), .x1158(x[1158]), .x1159(x[1159]), .x1160(x[1160]), .x1161(x[1161]), .x1162(x[1162]), .x1163(x[1163]), .x1164(x[1164]), .x1165(x[1165]), .x1166(x[1166]), .x1167(x[1167]), .x1168(x[1168]), .x1169(x[1169]), .x1170(x[1170]), .x1171(x[1171]), .x1172(x[1172]), .x1173(x[1173]), .x1174(x[1174]), .x1175(x[1175]), .x1176(x[1176]), .x1177(x[1177]), .x1178(x[1178]), .x1179(x[1179]), .x1180(x[1180]), .x1181(x[1181]), .x1182(x[1182]), .x1183(x[1183]), .x1184(x[1184]), .x1185(x[1185]), .x1186(x[1186]), .x1187(x[1187]), .x1188(x[1188]), .x1189(x[1189]), .x1190(x[1190]), .x1191(x[1191]), .x1192(x[1192]), .x1193(x[1193]), .x1194(x[1194]), .x1195(x[1195]), .x1196(x[1196]), .x1197(x[1197]), .x1198(x[1198]), .x1199(x[1199]), .x1200(x[1200]), .x1201(x[1201]), .x1202(x[1202]), .x1203(x[1203]), .x1204(x[1204]), .x1205(x[1205]), .x1206(x[1206]), .x1207(x[1207]), .x1208(x[1208]), .x1209(x[1209]), .x1210(x[1210]), .x1211(x[1211]), .x1212(x[1212]), .x1213(x[1213]), .x1214(x[1214]), .x1215(x[1215]), .x1216(x[1216]), .x1217(x[1217]), .x1218(x[1218]), .x1219(x[1219]), .x1220(x[1220]), .x1221(x[1221]), .x1222(x[1222]), .x1223(x[1223]), .x1224(x[1224]), .x1225(x[1225]), .x1226(x[1226]), .x1227(x[1227]), .x1228(x[1228]), .x1229(x[1229]), .x1230(x[1230]), .x1231(x[1231]), .x1232(x[1232]), .x1233(x[1233]), .x1234(x[1234]), .x1235(x[1235]), .x1236(x[1236]), .x1237(x[1237]), .x1238(x[1238]), .x1239(x[1239]), .x1240(x[1240]), .x1241(x[1241]), .x1242(x[1242]), .x1243(x[1243]), .x1244(x[1244]), .x1245(x[1245]), .x1246(x[1246]), .x1247(x[1247]), .x1248(x[1248]), .x1249(x[1249]), .x1250(x[1250]), .x1251(x[1251]), .x1252(x[1252]), .x1253(x[1253]), .x1254(x[1254]), .x1255(x[1255]), .x1256(x[1256]), .x1257(x[1257]), .x1258(x[1258]), .x1259(x[1259]), .x1260(x[1260]), .x1261(x[1261]), .x1262(x[1262]), .x1263(x[1263]), .x1264(x[1264]), .x1265(x[1265]), .x1266(x[1266]), .x1267(x[1267]), .x1268(x[1268]), .x1269(x[1269]), .x1270(x[1270]), .x1271(x[1271]), .x1272(x[1272]), .x1273(x[1273]), .x1274(x[1274]), .x1275(x[1275]), .x1276(x[1276]), .x1277(x[1277]), .x1278(x[1278]), .x1279(x[1279]), .x1280(x[1280]), .x1281(x[1281]), .x1282(x[1282]), .x1283(x[1283]), .x1284(x[1284]), .x1285(x[1285]), .x1286(x[1286]), .x1287(x[1287]), .x1288(x[1288]), .x1289(x[1289]), .x1290(x[1290]), .x1291(x[1291]), .x1292(x[1292]), .x1293(x[1293]), .x1294(x[1294]), .x1295(x[1295]), .x1296(x[1296]), .x1297(x[1297]), .x1298(x[1298]), .x1299(x[1299]), .x1300(x[1300]), .x1301(x[1301]), .x1302(x[1302]), .x1303(x[1303]), .x1304(x[1304]), .x1305(x[1305]), .x1306(x[1306]), .x1307(x[1307]), .x1308(x[1308]), .x1309(x[1309]), .x1310(x[1310]), .x1311(x[1311]), .x1312(x[1312]), .x1313(x[1313]), .x1314(x[1314]), .x1315(x[1315]), .x1316(x[1316]), .x1317(x[1317]), .x1318(x[1318]), .x1319(x[1319]), .x1320(x[1320]), .x1321(x[1321]), .x1322(x[1322]), .x1323(x[1323]), .x1324(x[1324]), .x1325(x[1325]), .x1326(x[1326]), .x1327(x[1327]), .x1328(x[1328]), .x1329(x[1329]), .x1330(x[1330]), .x1331(x[1331]), .x1332(x[1332]), .x1333(x[1333]), .x1334(x[1334]), .x1335(x[1335]), .x1336(x[1336]), .x1337(x[1337]), .x1338(x[1338]), .x1339(x[1339]), .x1340(x[1340]), .x1341(x[1341]), .x1342(x[1342]), .x1343(x[1343]), .x1344(x[1344]), .x1345(x[1345]), .x1346(x[1346]), .x1347(x[1347]), .x1348(x[1348]), .x1349(x[1349]), .x1350(x[1350]), .x1351(x[1351]), .x1352(x[1352]), .x1353(x[1353]), .x1354(x[1354]), .x1355(x[1355]), .x1356(x[1356]), .x1357(x[1357]), .x1358(x[1358]), .x1359(x[1359]), .x1360(x[1360]), .x1361(x[1361]), .x1362(x[1362]), .x1363(x[1363]), .x1364(x[1364]), .x1365(x[1365]), .x1366(x[1366]), .x1367(x[1367]), .x1368(x[1368]), .x1369(x[1369]), .x1370(x[1370]), .x1371(x[1371]), .x1372(x[1372]), .x1373(x[1373]), .x1374(x[1374]), .x1375(x[1375]), .x1376(x[1376]), .x1377(x[1377]), .x1378(x[1378]), .x1379(x[1379]), .x1380(x[1380]), .x1381(x[1381]), .x1382(x[1382]), .x1383(x[1383]), .x1384(x[1384]), .x1385(x[1385]), .x1386(x[1386]), .x1387(x[1387]), .x1388(x[1388]), .x1389(x[1389]), .x1390(x[1390]), .x1391(x[1391]), .x1392(x[1392]), .x1393(x[1393]), .x1394(x[1394]), .x1395(x[1395]), .x1396(x[1396]), .x1397(x[1397]), .x1398(x[1398]), .x1399(x[1399]), .x1400(x[1400]), .x1401(x[1401]), .x1402(x[1402]), .x1403(x[1403]), .x1404(x[1404]), .x1405(x[1405]), .x1406(x[1406]), .x1407(x[1407]), .x1408(x[1408]), .x1409(x[1409]), .x1410(x[1410]), .x1411(x[1411]), .x1412(x[1412]), .x1413(x[1413]), .x1414(x[1414]), .x1415(x[1415]), .x1416(x[1416]), .x1417(x[1417]), .x1418(x[1418]), .x1419(x[1419]), .x1420(x[1420]), .x1421(x[1421]), .x1422(x[1422]), .x1423(x[1423]), .x1424(x[1424]), .x1425(x[1425]), .x1426(x[1426]), .x1427(x[1427]), .x1428(x[1428]), .x1429(x[1429]), .x1430(x[1430]), .x1431(x[1431]), .x1432(x[1432]), .x1433(x[1433]), .x1434(x[1434]), .x1435(x[1435]), .x1436(x[1436]), .x1437(x[1437]), .x1438(x[1438]), .x1439(x[1439]), .x1440(x[1440]), .x1441(x[1441]), .x1442(x[1442]), .x1443(x[1443]), .x1444(x[1444]), .x1445(x[1445]), .x1446(x[1446]), .x1447(x[1447]), .x1448(x[1448]), .x1449(x[1449]), .x1450(x[1450]), .x1451(x[1451]), .x1452(x[1452]), .x1453(x[1453]), .x1454(x[1454]), .x1455(x[1455]), .x1456(x[1456]), .x1457(x[1457]), .x1458(x[1458]), .x1459(x[1459]), .x1460(x[1460]), .x1461(x[1461]), .x1462(x[1462]), .x1463(x[1463]), .x1464(x[1464]), .x1465(x[1465]), .x1466(x[1466]), .x1467(x[1467]), .x1468(x[1468]), .x1469(x[1469]), .x1470(x[1470]), .x1471(x[1471]), .x1472(x[1472]), .x1473(x[1473]), .x1474(x[1474]), .x1475(x[1475]), .x1476(x[1476]), .x1477(x[1477]), .x1478(x[1478]), .x1479(x[1479]), .x1480(x[1480]), .x1481(x[1481]), .x1482(x[1482]), .x1483(x[1483]), .x1484(x[1484]), .x1485(x[1485]), .x1486(x[1486]), .x1487(x[1487]), .x1488(x[1488]), .x1489(x[1489]), .x1490(x[1490]), .x1491(x[1491]), .x1492(x[1492]), .x1493(x[1493]), .x1494(x[1494]), .x1495(x[1495]), .x1496(x[1496]), .x1497(x[1497]), .x1498(x[1498]), .x1499(x[1499]), .x1500(x[1500]), .x1501(x[1501]), .x1502(x[1502]), .x1503(x[1503]), .x1504(x[1504]), .x1505(x[1505]), .x1506(x[1506]), .x1507(x[1507]), .x1508(x[1508]), .x1509(x[1509]), .x1510(x[1510]), .x1511(x[1511]), .x1512(x[1512]), .x1513(x[1513]), .x1514(x[1514]), .x1515(x[1515]), .x1516(x[1516]), .x1517(x[1517]), .x1518(x[1518]), .x1519(x[1519]), .x1520(x[1520]), .x1521(x[1521]), .x1522(x[1522]), .x1523(x[1523]), .x1524(x[1524]), .x1525(x[1525]), .x1526(x[1526]), .x1527(x[1527]), .x1528(x[1528]), .x1529(x[1529]), .x1530(x[1530]), .x1531(x[1531]), .x1532(x[1532]), .x1533(x[1533]), .x1534(x[1534]), .x1535(x[1535]), .x1536(x[1536]), .x1537(x[1537]), .x1538(x[1538]), .x1539(x[1539]), .x1540(x[1540]), .x1541(x[1541]), .x1542(x[1542]), .x1543(x[1543]), .x1544(x[1544]), .x1545(x[1545]), .x1546(x[1546]), .x1547(x[1547]), .x1548(x[1548]), .x1549(x[1549]), .x1550(x[1550]), .x1551(x[1551]), .x1552(x[1552]), .x1553(x[1553]), .x1554(x[1554]), .x1555(x[1555]), .x1556(x[1556]), .x1557(x[1557]), .x1558(x[1558]), .x1559(x[1559]), .x1560(x[1560]), .x1561(x[1561]), .x1562(x[1562]), .x1563(x[1563]), .x1564(x[1564]), .x1565(x[1565]), .x1566(x[1566]), .x1567(x[1567]), .x1568(x[1568]), .x1569(x[1569]), .x1570(x[1570]), .x1571(x[1571]), .x1572(x[1572]), .x1573(x[1573]), .x1574(x[1574]), .x1575(x[1575]), .x1576(x[1576]), .x1577(x[1577]), .x1578(x[1578]), .x1579(x[1579]), .x1580(x[1580]), .x1581(x[1581]), .x1582(x[1582]), .x1583(x[1583]), .x1584(x[1584]), .x1585(x[1585]), .x1586(x[1586]), .x1587(x[1587]), .x1588(x[1588]), .x1589(x[1589]), .x1590(x[1590]), .x1591(x[1591]), .x1592(x[1592]), .x1593(x[1593]), .x1594(x[1594]), .x1595(x[1595]), .x1596(x[1596]), .x1597(x[1597]), .x1598(x[1598]), .x1599(x[1599]), .x1600(x[1600]), .x1601(x[1601]), .x1602(x[1602]), .x1603(x[1603]), .x1604(x[1604]), .x1605(x[1605]), .x1606(x[1606]), .x1607(x[1607]), .x1608(x[1608]), .x1609(x[1609]), .x1610(x[1610]), .x1611(x[1611]), .x1612(x[1612]), .x1613(x[1613]), .x1614(x[1614]), .x1615(x[1615]), .x1616(x[1616]), .x1617(x[1617]), .x1618(x[1618]), .x1619(x[1619]), .x1620(x[1620]), .x1621(x[1621]), .x1622(x[1622]), .x1623(x[1623]), .x1624(x[1624]), .x1625(x[1625]), .x1626(x[1626]), .x1627(x[1627]), .x1628(x[1628]), .x1629(x[1629]), .x1630(x[1630]), .x1631(x[1631]), .x1632(x[1632]), .x1633(x[1633]), .x1634(x[1634]), .x1635(x[1635]), .x1636(x[1636]), .x1637(x[1637]), .x1638(x[1638]), .x1639(x[1639]), .x1640(x[1640]), .x1641(x[1641]), .x1642(x[1642]), .x1643(x[1643]), .x1644(x[1644]), .x1645(x[1645]), .x1646(x[1646]), .x1647(x[1647]), .x1648(x[1648]), .x1649(x[1649]), .x1650(x[1650]), .x1651(x[1651]), .x1652(x[1652]), .x1653(x[1653]), .x1654(x[1654]), .x1655(x[1655]), .x1656(x[1656]), .x1657(x[1657]), .x1658(x[1658]), .x1659(x[1659]), .x1660(x[1660]), .x1661(x[1661]), .x1662(x[1662]), .x1663(x[1663]), .x1664(x[1664]), .x1665(x[1665]), .x1666(x[1666]), .x1667(x[1667]), .x1668(x[1668]), .x1669(x[1669]), .x1670(x[1670]), .x1671(x[1671]), .x1672(x[1672]), .x1673(x[1673]), .x1674(x[1674]), .x1675(x[1675]), .x1676(x[1676]), .x1677(x[1677]), .x1678(x[1678]), .x1679(x[1679]), .x1680(x[1680]), .x1681(x[1681]), .x1682(x[1682]), .x1683(x[1683]), .x1684(x[1684]), .x1685(x[1685]), .x1686(x[1686]), .x1687(x[1687]), .x1688(x[1688]), .x1689(x[1689]), .x1690(x[1690]), .x1691(x[1691]), .x1692(x[1692]), .x1693(x[1693]), .x1694(x[1694]), .x1695(x[1695]), .x1696(x[1696]), .x1697(x[1697]), .x1698(x[1698]), .x1699(x[1699]), .x1700(x[1700]), .x1701(x[1701]), .x1702(x[1702]), .x1703(x[1703]), .x1704(x[1704]), .x1705(x[1705]), .x1706(x[1706]), .x1707(x[1707]), .x1708(x[1708]), .x1709(x[1709]), .x1710(x[1710]), .x1711(x[1711]), .x1712(x[1712]), .x1713(x[1713]), .x1714(x[1714]), .x1715(x[1715]), .x1716(x[1716]), .x1717(x[1717]), .x1718(x[1718]), .x1719(x[1719]), .x1720(x[1720]), .x1721(x[1721]), .x1722(x[1722]), .x1723(x[1723]), .x1724(x[1724]), .x1725(x[1725]), .x1726(x[1726]), .x1727(x[1727]), .x1728(x[1728]), .x1729(x[1729]), .x1730(x[1730]), .x1731(x[1731]), .x1732(x[1732]), .x1733(x[1733]), .x1734(x[1734]), .x1735(x[1735]), .x1736(x[1736]), .x1737(x[1737]), .x1738(x[1738]), .x1739(x[1739]), .x1740(x[1740]), .x1741(x[1741]), .x1742(x[1742]), .x1743(x[1743]), .x1744(x[1744]), .x1745(x[1745]), .x1746(x[1746]), .x1747(x[1747]), .x1748(x[1748]), .x1749(x[1749]), .x1750(x[1750]), .x1751(x[1751]), .x1752(x[1752]), .x1753(x[1753]), .x1754(x[1754]), .x1755(x[1755]), .x1756(x[1756]), .x1757(x[1757]), .x1758(x[1758]), .x1759(x[1759]), .x1760(x[1760]), .x1761(x[1761]), .x1762(x[1762]), .x1763(x[1763]), .x1764(x[1764]), .x1765(x[1765]), .x1766(x[1766]), .x1767(x[1767]), .x1768(x[1768]), .x1769(x[1769]), .x1770(x[1770]), .x1771(x[1771]), .x1772(x[1772]), .x1773(x[1773]), .x1774(x[1774]), .x1775(x[1775]), .x1776(x[1776]), .x1777(x[1777]), .x1778(x[1778]), .x1779(x[1779]), .x1780(x[1780]), .x1781(x[1781]), .x1782(x[1782]), .x1783(x[1783]), .x1784(x[1784]), .x1785(x[1785]), .x1786(x[1786]), .x1787(x[1787]), .x1788(x[1788]), .x1789(x[1789]), .x1790(x[1790]), .x1791(x[1791]), .x1792(x[1792]), .x1793(x[1793]), .x1794(x[1794]), .x1795(x[1795]), .x1796(x[1796]), .x1797(x[1797]), .x1798(x[1798]), .x1799(x[1799]), .x1800(x[1800]), .x1801(x[1801]), .x1802(x[1802]), .x1803(x[1803]), .x1804(x[1804]), .x1805(x[1805]), .x1806(x[1806]), .x1807(x[1807]), .x1808(x[1808]), .x1809(x[1809]), .x1810(x[1810]), .x1811(x[1811]), .x1812(x[1812]), .x1813(x[1813]), .x1814(x[1814]), .x1815(x[1815]), .x1816(x[1816]), .x1817(x[1817]), .x1818(x[1818]), .x1819(x[1819]), .x1820(x[1820]), .x1821(x[1821]), .x1822(x[1822]), .x1823(x[1823]), .x1824(x[1824]), .x1825(x[1825]), .x1826(x[1826]), .x1827(x[1827]), .x1828(x[1828]), .x1829(x[1829]), .x1830(x[1830]), .x1831(x[1831]), .x1832(x[1832]), .x1833(x[1833]), .x1834(x[1834]), .x1835(x[1835]), .x1836(x[1836]), .x1837(x[1837]), .x1838(x[1838]), .x1839(x[1839]), .x1840(x[1840]), .x1841(x[1841]), .x1842(x[1842]), .x1843(x[1843]), .x1844(x[1844]), .x1845(x[1845]), .x1846(x[1846]), .x1847(x[1847]), .x1848(x[1848]), .x1849(x[1849]), .x1850(x[1850]), .x1851(x[1851]), .x1852(x[1852]), .x1853(x[1853]), .x1854(x[1854]), .x1855(x[1855]), .x1856(x[1856]), .x1857(x[1857]), .x1858(x[1858]), .x1859(x[1859]), .x1860(x[1860]), .x1861(x[1861]), .x1862(x[1862]), .x1863(x[1863]), .x1864(x[1864]), .x1865(x[1865]), .x1866(x[1866]), .x1867(x[1867]), .x1868(x[1868]), .x1869(x[1869]), .x1870(x[1870]), .x1871(x[1871]), .x1872(x[1872]), .x1873(x[1873]), .x1874(x[1874]), .x1875(x[1875]), .x1876(x[1876]), .x1877(x[1877]), .x1878(x[1878]), .x1879(x[1879]), .x1880(x[1880]), .x1881(x[1881]), .x1882(x[1882]), .x1883(x[1883]), .x1884(x[1884]), .x1885(x[1885]), .x1886(x[1886]), .x1887(x[1887]), .x1888(x[1888]), .x1889(x[1889]), .x1890(x[1890]), .x1891(x[1891]), .x1892(x[1892]), .x1893(x[1893]), .x1894(x[1894]), .x1895(x[1895]), .x1896(x[1896]), .x1897(x[1897]), .x1898(x[1898]), .x1899(x[1899]), .x1900(x[1900]), .x1901(x[1901]), .x1902(x[1902]), .x1903(x[1903]), .x1904(x[1904]), .x1905(x[1905]), .x1906(x[1906]), .x1907(x[1907]), .x1908(x[1908]), .x1909(x[1909]), .x1910(x[1910]), .x1911(x[1911]), .x1912(x[1912]), .x1913(x[1913]), .x1914(x[1914]), .x1915(x[1915]), .x1916(x[1916]), .x1917(x[1917]), .x1918(x[1918]), .x1919(x[1919]), .x1920(x[1920]), .x1921(x[1921]), .x1922(x[1922]), .x1923(x[1923]), .x1924(x[1924]), .x1925(x[1925]), .x1926(x[1926]), .x1927(x[1927]), .x1928(x[1928]), .x1929(x[1929]), .x1930(x[1930]), .x1931(x[1931]), .x1932(x[1932]), .x1933(x[1933]), .x1934(x[1934]), .x1935(x[1935]), .x1936(x[1936]), .x1937(x[1937]), .x1938(x[1938]), .x1939(x[1939]), .x1940(x[1940]), .x1941(x[1941]), .x1942(x[1942]), .x1943(x[1943]), .x1944(x[1944]), .x1945(x[1945]), .x1946(x[1946]), .x1947(x[1947]), .x1948(x[1948]), .x1949(x[1949]), .x1950(x[1950]), .x1951(x[1951]), .x1952(x[1952]), .x1953(x[1953]), .x1954(x[1954]), .x1955(x[1955]), .x1956(x[1956]), .x1957(x[1957]), .x1958(x[1958]), .x1959(x[1959]), .x1960(x[1960]), .x1961(x[1961]), .x1962(x[1962]), .x1963(x[1963]), .x1964(x[1964]), .x1965(x[1965]), .x1966(x[1966]), .x1967(x[1967]), .x1968(x[1968]), .x1969(x[1969]), .x1970(x[1970]), .x1971(x[1971]), .x1972(x[1972]), .x1973(x[1973]), .x1974(x[1974]), .x1975(x[1975]), .x1976(x[1976]), .x1977(x[1977]), .x1978(x[1978]), .x1979(x[1979]), .x1980(x[1980]), .x1981(x[1981]), .x1982(x[1982]), .x1983(x[1983]), .x1984(x[1984]), .x1985(x[1985]), .x1986(x[1986]), .x1987(x[1987]), .x1988(x[1988]), .x1989(x[1989]), .x1990(x[1990]), .x1991(x[1991]), .x1992(x[1992]), .x1993(x[1993]), .x1994(x[1994]), .x1995(x[1995]), .x1996(x[1996]), .x1997(x[1997]), .x1998(x[1998]), .x1999(x[1999]), .x2000(x[2000]), .x2001(x[2001]), .x2002(x[2002]), .x2003(x[2003]), .x2004(x[2004]), .x2005(x[2005]), .x2006(x[2006]), .x2007(x[2007]), .x2008(x[2008]), .x2009(x[2009]), .x2010(x[2010]), .x2011(x[2011]), .x2012(x[2012]), .x2013(x[2013]), .x2014(x[2014]), .x2015(x[2015]), .x2016(x[2016]), .x2017(x[2017]), .x2018(x[2018]), .x2019(x[2019]), .x2020(x[2020]), .x2021(x[2021]), .x2022(x[2022]), .x2023(x[2023]), .x2024(x[2024]), .x2025(x[2025]), .x2026(x[2026]), .x2027(x[2027]), .x2028(x[2028]), .x2029(x[2029]), .x2030(x[2030]), .x2031(x[2031]), .x2032(x[2032]), .x2033(x[2033]), .x2034(x[2034]), .x2035(x[2035]), .x2036(x[2036]), .x2037(x[2037]), .x2038(x[2038]), .x2039(x[2039]), .x2040(x[2040]), .x2041(x[2041]), .x2042(x[2042]), .x2043(x[2043]), .x2044(x[2044]), .x2045(x[2045]), .x2046(x[2046]), .x2047(x[2047]), .x2048(x[2048]), .x2049(x[2049]), .x2050(x[2050]), .x2051(x[2051]), .x2052(x[2052]), .x2053(x[2053]), .x2054(x[2054]), .x2055(x[2055]), .x2056(x[2056]), .x2057(x[2057]), .x2058(x[2058]), .x2059(x[2059]), .x2060(x[2060]), .x2061(x[2061]), .x2062(x[2062]), .x2063(x[2063]), .x2064(x[2064]), .x2065(x[2065]), .x2066(x[2066]), .x2067(x[2067]), .x2068(x[2068]), .x2069(x[2069]), .x2070(x[2070]), .x2071(x[2071]), .x2072(x[2072]), .x2073(x[2073]), .x2074(x[2074]), .x2075(x[2075]), .x2076(x[2076]), .x2077(x[2077]), .x2078(x[2078]), .x2079(x[2079]), .x2080(x[2080]), .x2081(x[2081]), .x2082(x[2082]), .x2083(x[2083]), .x2084(x[2084]), .x2085(x[2085]), .x2086(x[2086]), .x2087(x[2087]), .x2088(x[2088]), .x2089(x[2089]), .x2090(x[2090]), .x2091(x[2091]), .x2092(x[2092]), .x2093(x[2093]), .x2094(x[2094]), .x2095(x[2095]), .x2096(x[2096]), .x2097(x[2097]), .x2098(x[2098]), .x2099(x[2099]), .x2100(x[2100]), .x2101(x[2101]), .x2102(x[2102]), .x2103(x[2103]), .x2104(x[2104]), .x2105(x[2105]), .x2106(x[2106]), .x2107(x[2107]), .x2108(x[2108]), .x2109(x[2109]), .x2110(x[2110]), .x2111(x[2111]), .x2112(x[2112]), .x2113(x[2113]), .x2114(x[2114]), .x2115(x[2115]), .x2116(x[2116]), .x2117(x[2117]), .x2118(x[2118]), .x2119(x[2119]), .x2120(x[2120]), .x2121(x[2121]), .x2122(x[2122]), .x2123(x[2123]), .x2124(x[2124]), .x2125(x[2125]), .x2126(x[2126]), .x2127(x[2127]), .x2128(x[2128]), .x2129(x[2129]), .x2130(x[2130]), .x2131(x[2131]), .x2132(x[2132]), .x2133(x[2133]), .x2134(x[2134]), .x2135(x[2135]), .x2136(x[2136]), .x2137(x[2137]), .x2138(x[2138]), .x2139(x[2139]), .x2140(x[2140]), .x2141(x[2141]), .x2142(x[2142]), .x2143(x[2143]), .x2144(x[2144]), .x2145(x[2145]), .x2146(x[2146]), .x2147(x[2147]), .x2148(x[2148]), .x2149(x[2149]), .x2150(x[2150]), .x2151(x[2151]), .x2152(x[2152]), .x2153(x[2153]), .x2154(x[2154]), .x2155(x[2155]), .x2156(x[2156]), .x2157(x[2157]), .x2158(x[2158]), .x2159(x[2159]), .x2160(x[2160]), .x2161(x[2161]), .x2162(x[2162]), .x2163(x[2163]), .x2164(x[2164]), .x2165(x[2165]), .x2166(x[2166]), .x2167(x[2167]), .x2168(x[2168]), .x2169(x[2169]), .x2170(x[2170]), .x2171(x[2171]), .x2172(x[2172]), .x2173(x[2173]), .x2174(x[2174]), .x2175(x[2175]), .x2176(x[2176]), .x2177(x[2177]), .x2178(x[2178]), .x2179(x[2179]), .x2180(x[2180]), .x2181(x[2181]), .x2182(x[2182]), .x2183(x[2183]), .x2184(x[2184]), .x2185(x[2185]), .x2186(x[2186]), .x2187(x[2187]), .x2188(x[2188]), .x2189(x[2189]), .x2190(x[2190]), .x2191(x[2191]), .x2192(x[2192]), .x2193(x[2193]), .x2194(x[2194]), .x2195(x[2195]), .x2196(x[2196]), .x2197(x[2197]), .x2198(x[2198]), .x2199(x[2199]), .x2200(x[2200]), .x2201(x[2201]), .x2202(x[2202]), .x2203(x[2203]), .x2204(x[2204]), .x2205(x[2205]), .x2206(x[2206]), .x2207(x[2207]), .x2208(x[2208]), .x2209(x[2209]), .x2210(x[2210]), .x2211(x[2211]), .x2212(x[2212]), .x2213(x[2213]), .x2214(x[2214]), .x2215(x[2215]), .x2216(x[2216]), .x2217(x[2217]), .x2218(x[2218]), .x2219(x[2219]), .x2220(x[2220]), .x2221(x[2221]), .x2222(x[2222]), .x2223(x[2223]), .x2224(x[2224]), .x2225(x[2225]), .x2226(x[2226]), .x2227(x[2227]), .x2228(x[2228]), .x2229(x[2229]), .x2230(x[2230]), .x2231(x[2231]), .x2232(x[2232]), .x2233(x[2233]), .x2234(x[2234]), .x2235(x[2235]), .x2236(x[2236]), .x2237(x[2237]), .x2238(x[2238]), .x2239(x[2239]), .x2240(x[2240]), .x2241(x[2241]), .x2242(x[2242]), .x2243(x[2243]), .x2244(x[2244]), .x2245(x[2245]), .x2246(x[2246]), .x2247(x[2247]), .x2248(x[2248]), .x2249(x[2249]), .x2250(x[2250]), .x2251(x[2251]), .x2252(x[2252]), .x2253(x[2253]), .x2254(x[2254]), .x2255(x[2255]), .x2256(x[2256]), .x2257(x[2257]), .x2258(x[2258]), .x2259(x[2259]), .x2260(x[2260]), .x2261(x[2261]), .x2262(x[2262]), .x2263(x[2263]), .x2264(x[2264]), .x2265(x[2265]), .x2266(x[2266]), .x2267(x[2267]), .x2268(x[2268]), .x2269(x[2269]), .x2270(x[2270]), .x2271(x[2271]), .x2272(x[2272]), .x2273(x[2273]), .x2274(x[2274]), .x2275(x[2275]), .x2276(x[2276]), .x2277(x[2277]), .x2278(x[2278]), .x2279(x[2279]), .x2280(x[2280]), .x2281(x[2281]), .x2282(x[2282]), .x2283(x[2283]), .x2284(x[2284]), .x2285(x[2285]), .x2286(x[2286]), .x2287(x[2287]), .x2288(x[2288]), .x2289(x[2289]), .x2290(x[2290]), .x2291(x[2291]), .x2292(x[2292]), .x2293(x[2293]), .x2294(x[2294]), .x2295(x[2295]), .x2296(x[2296]), .x2297(x[2297]), .x2298(x[2298]), .x2299(x[2299]), .x2300(x[2300]), .x2301(x[2301]), .x2302(x[2302]), .x2303(x[2303]), .x2304(x[2304]), .x2305(x[2305]), .x2306(x[2306]), .x2307(x[2307]), .x2308(x[2308]), .x2309(x[2309]), .x2310(x[2310]), .x2311(x[2311]), .x2312(x[2312]), .x2313(x[2313]), .x2314(x[2314]), .x2315(x[2315]), .x2316(x[2316]), .x2317(x[2317]), .x2318(x[2318]), .x2319(x[2319]), .x2320(x[2320]), .x2321(x[2321]), .x2322(x[2322]), .x2323(x[2323]), .x2324(x[2324]), .x2325(x[2325]), .x2326(x[2326]), .x2327(x[2327]), .x2328(x[2328]), .x2329(x[2329]), .x2330(x[2330]), .x2331(x[2331]), .x2332(x[2332]), .x2333(x[2333]), .x2334(x[2334]), .x2335(x[2335]), .x2336(x[2336]), .x2337(x[2337]), .x2338(x[2338]), .x2339(x[2339]), .x2340(x[2340]), .x2341(x[2341]), .x2342(x[2342]), .x2343(x[2343]), .x2344(x[2344]), .x2345(x[2345]), .x2346(x[2346]), .x2347(x[2347]), .x2348(x[2348]), .x2349(x[2349]), .x2350(x[2350]), .x2351(x[2351]), .x2352(x[2352]), .x2353(x[2353]), .x2354(x[2354]), .x2355(x[2355]), .x2356(x[2356]), .x2357(x[2357]), .x2358(x[2358]), .x2359(x[2359]), .x2360(x[2360]), .x2361(x[2361]), .x2362(x[2362]), .x2363(x[2363]), .x2364(x[2364]), .x2365(x[2365]), .x2366(x[2366]), .x2367(x[2367]), .x2368(x[2368]), .x2369(x[2369]), .x2370(x[2370]), .x2371(x[2371]), .x2372(x[2372]), .x2373(x[2373]), .x2374(x[2374]), .x2375(x[2375]), .x2376(x[2376]), .x2377(x[2377]), .x2378(x[2378]), .x2379(x[2379]), .x2380(x[2380]), .x2381(x[2381]), .x2382(x[2382]), .x2383(x[2383]), .x2384(x[2384]), .x2385(x[2385]), .x2386(x[2386]), .x2387(x[2387]), .x2388(x[2388]), .x2389(x[2389]), .x2390(x[2390]), .x2391(x[2391]), .x2392(x[2392]), .x2393(x[2393]), .x2394(x[2394]), .x2395(x[2395]), .x2396(x[2396]), .x2397(x[2397]), .x2398(x[2398]), .x2399(x[2399]), .x2400(x[2400]), .x2401(x[2401]), .x2402(x[2402]), .x2403(x[2403]), .x2404(x[2404]), .x2405(x[2405]), .x2406(x[2406]), .x2407(x[2407]), .x2408(x[2408]), .x2409(x[2409]), .x2410(x[2410]), .x2411(x[2411]), .x2412(x[2412]), .x2413(x[2413]), .x2414(x[2414]), .x2415(x[2415]), .x2416(x[2416]), .x2417(x[2417]), .x2418(x[2418]), .x2419(x[2419]), .x2420(x[2420]), .x2421(x[2421]), .x2422(x[2422]), .x2423(x[2423]), .x2424(x[2424]), .x2425(x[2425]), .x2426(x[2426]), .x2427(x[2427]), .x2428(x[2428]), .x2429(x[2429]), .x2430(x[2430]), .x2431(x[2431]), .x2432(x[2432]), .x2433(x[2433]), .x2434(x[2434]), .x2435(x[2435]), .x2436(x[2436]), .x2437(x[2437]), .x2438(x[2438]), .x2439(x[2439]), .x2440(x[2440]), .x2441(x[2441]), .x2442(x[2442]), .x2443(x[2443]), .x2444(x[2444]), .x2445(x[2445]), .x2446(x[2446]), .x2447(x[2447]), .x2448(x[2448]), .x2449(x[2449]), .x2450(x[2450]), .x2451(x[2451]), .x2452(x[2452]), .x2453(x[2453]), .x2454(x[2454]), .x2455(x[2455]), .x2456(x[2456]), .x2457(x[2457]), .x2458(x[2458]), .x2459(x[2459]), .x2460(x[2460]), .x2461(x[2461]), .x2462(x[2462]), .x2463(x[2463]), .x2464(x[2464]), .x2465(x[2465]), .x2466(x[2466]), .x2467(x[2467]), .x2468(x[2468]), .x2469(x[2469]), .x2470(x[2470]), .x2471(x[2471]), .x2472(x[2472]), .x2473(x[2473]), .x2474(x[2474]), .x2475(x[2475]), .x2476(x[2476]), .x2477(x[2477]), .x2478(x[2478]), .x2479(x[2479]), .x2480(x[2480]), .x2481(x[2481]), .x2482(x[2482]), .x2483(x[2483]), .x2484(x[2484]), .x2485(x[2485]), .x2486(x[2486]), .x2487(x[2487]), .x2488(x[2488]), .x2489(x[2489]), .x2490(x[2490]), .x2491(x[2491]), .x2492(x[2492]), .x2493(x[2493]), .x2494(x[2494]), .x2495(x[2495]), .x2496(x[2496]), .x2497(x[2497]), .x2498(x[2498]), .x2499(x[2499]), .x2500(x[2500]), .x2501(x[2501]), .x2502(x[2502]), .x2503(x[2503]), .x2504(x[2504]), .x2505(x[2505]), .x2506(x[2506]), .x2507(x[2507]), .x2508(x[2508]), .x2509(x[2509]), .x2510(x[2510]), .x2511(x[2511]), .x2512(x[2512]), .x2513(x[2513]), .x2514(x[2514]), .x2515(x[2515]), .x2516(x[2516]), .x2517(x[2517]), .x2518(x[2518]), .x2519(x[2519]), .x2520(x[2520]), .x2521(x[2521]), .x2522(x[2522]), .x2523(x[2523]), .x2524(x[2524]), .x2525(x[2525]), .x2526(x[2526]), .x2527(x[2527]), .x2528(x[2528]), .x2529(x[2529]), .x2530(x[2530]), .x2531(x[2531]), .x2532(x[2532]), .x2533(x[2533]), .x2534(x[2534]), .x2535(x[2535]), .x2536(x[2536]), .x2537(x[2537]), .x2538(x[2538]), .x2539(x[2539]), .x2540(x[2540]), .x2541(x[2541]), .x2542(x[2542]), .x2543(x[2543]), .x2544(x[2544]), .x2545(x[2545]), .x2546(x[2546]), .x2547(x[2547]), .x2548(x[2548]), .x2549(x[2549]), .x2550(x[2550]), .x2551(x[2551]), .x2552(x[2552]), .x2553(x[2553]), .x2554(x[2554]), .x2555(x[2555]), .x2556(x[2556]), .x2557(x[2557]), .x2558(x[2558]), .x2559(x[2559]), .x2560(x[2560]), .x2561(x[2561]), .x2562(x[2562]), .x2563(x[2563]), .x2564(x[2564]), .x2565(x[2565]), .x2566(x[2566]), .x2567(x[2567]), .x2568(x[2568]), .x2569(x[2569]), .x2570(x[2570]), .x2571(x[2571]), .x2572(x[2572]), .x2573(x[2573]), .x2574(x[2574]), .x2575(x[2575]), .x2576(x[2576]), .x2577(x[2577]), .x2578(x[2578]), .x2579(x[2579]), .x2580(x[2580]), .x2581(x[2581]), .x2582(x[2582]), .x2583(x[2583]), .x2584(x[2584]), .x2585(x[2585]), .x2586(x[2586]), .x2587(x[2587]), .x2588(x[2588]), .x2589(x[2589]), .x2590(x[2590]), .x2591(x[2591]), .x2592(x[2592]), .x2593(x[2593]), .x2594(x[2594]), .x2595(x[2595]), .x2596(x[2596]), .x2597(x[2597]), .x2598(x[2598]), .x2599(x[2599]), .x2600(x[2600]), .x2601(x[2601]), .x2602(x[2602]), .x2603(x[2603]), .x2604(x[2604]), .x2605(x[2605]), .x2606(x[2606]), .x2607(x[2607]), .x2608(x[2608]), .x2609(x[2609]), .x2610(x[2610]), .x2611(x[2611]), .x2612(x[2612]), .x2613(x[2613]), .x2614(x[2614]), .x2615(x[2615]), .x2616(x[2616]), .x2617(x[2617]), .x2618(x[2618]), .x2619(x[2619]), .x2620(x[2620]), .x2621(x[2621]), .x2622(x[2622]), .x2623(x[2623]), .x2624(x[2624]), .x2625(x[2625]), .x2626(x[2626]), .x2627(x[2627]), .x2628(x[2628]), .x2629(x[2629]), .x2630(x[2630]), .x2631(x[2631]), .x2632(x[2632]), .x2633(x[2633]), .x2634(x[2634]), .x2635(x[2635]), .x2636(x[2636]), .x2637(x[2637]), .x2638(x[2638]), .x2639(x[2639]), .x2640(x[2640]), .x2641(x[2641]), .x2642(x[2642]), .x2643(x[2643]), .x2644(x[2644]), .x2645(x[2645]), .x2646(x[2646]), .x2647(x[2647]), .x2648(x[2648]), .x2649(x[2649]), .x2650(x[2650]), .x2651(x[2651]), .x2652(x[2652]), .x2653(x[2653]), .x2654(x[2654]), .x2655(x[2655]), .x2656(x[2656]), .x2657(x[2657]), .x2658(x[2658]), .x2659(x[2659]), .x2660(x[2660]), .x2661(x[2661]), .x2662(x[2662]), .x2663(x[2663]), .x2664(x[2664]), .x2665(x[2665]), .x2666(x[2666]), .x2667(x[2667]), .x2668(x[2668]), .x2669(x[2669]), .x2670(x[2670]), .x2671(x[2671]), .x2672(x[2672]), .x2673(x[2673]), .x2674(x[2674]), .x2675(x[2675]), .x2676(x[2676]), .x2677(x[2677]), .x2678(x[2678]), .x2679(x[2679]), .x2680(x[2680]), .x2681(x[2681]), .x2682(x[2682]), .x2683(x[2683]), .x2684(x[2684]), .x2685(x[2685]), .x2686(x[2686]), .x2687(x[2687]), .x2688(x[2688]), .x2689(x[2689]), .x2690(x[2690]), .x2691(x[2691]), .x2692(x[2692]), .x2693(x[2693]), .x2694(x[2694]), .x2695(x[2695]), .x2696(x[2696]), .x2697(x[2697]), .x2698(x[2698]), .x2699(x[2699]), .x2700(x[2700]), .x2701(x[2701]), .x2702(x[2702]), .x2703(x[2703]), .x2704(x[2704]), .x2705(x[2705]), .x2706(x[2706]), .x2707(x[2707]), .x2708(x[2708]), .x2709(x[2709]), .x2710(x[2710]), .x2711(x[2711]), .x2712(x[2712]), .x2713(x[2713]), .x2714(x[2714]), .x2715(x[2715]), .x2716(x[2716]), .x2717(x[2717]), .x2718(x[2718]), .x2719(x[2719]), .x2720(x[2720]), .x2721(x[2721]), .x2722(x[2722]), .x2723(x[2723]), .x2724(x[2724]), .x2725(x[2725]), .x2726(x[2726]), .x2727(x[2727]), .x2728(x[2728]), .x2729(x[2729]), .x2730(x[2730]), .x2731(x[2731]), .x2732(x[2732]), .x2733(x[2733]), .x2734(x[2734]), .x2735(x[2735]), .x2736(x[2736]), .x2737(x[2737]), .x2738(x[2738]), .x2739(x[2739]), .x2740(x[2740]), .x2741(x[2741]), .x2742(x[2742]), .x2743(x[2743]), .x2744(x[2744]), .x2745(x[2745]), .x2746(x[2746]), .x2747(x[2747]), .x2748(x[2748]), .x2749(x[2749]), .x2750(x[2750]), .x2751(x[2751]), .x2752(x[2752]), .x2753(x[2753]), .x2754(x[2754]), .x2755(x[2755]), .x2756(x[2756]), .x2757(x[2757]), .x2758(x[2758]), .x2759(x[2759]), .x2760(x[2760]), .x2761(x[2761]), .x2762(x[2762]), .x2763(x[2763]), .x2764(x[2764]), .x2765(x[2765]), .x2766(x[2766]), .x2767(x[2767]), .x2768(x[2768]), .x2769(x[2769]), .x2770(x[2770]), .x2771(x[2771]), .x2772(x[2772]), .x2773(x[2773]), .x2774(x[2774]), .x2775(x[2775]), .x2776(x[2776]), .x2777(x[2777]), .x2778(x[2778]), .x2779(x[2779]), .x2780(x[2780]), .x2781(x[2781]), .x2782(x[2782]), .x2783(x[2783]), .x2784(x[2784]), .x2785(x[2785]), .x2786(x[2786]), .x2787(x[2787]), .x2788(x[2788]), .x2789(x[2789]), .x2790(x[2790]), .x2791(x[2791]), .x2792(x[2792]), .x2793(x[2793]), .x2794(x[2794]), .x2795(x[2795]), .x2796(x[2796]), .x2797(x[2797]), .x2798(x[2798]), .x2799(x[2799]), .x2800(x[2800]), .x2801(x[2801]), .x2802(x[2802]), .x2803(x[2803]), .x2804(x[2804]), .x2805(x[2805]), .x2806(x[2806]), .x2807(x[2807]), .x2808(x[2808]), .x2809(x[2809]), .x2810(x[2810]), .x2811(x[2811]), .x2812(x[2812]), .x2813(x[2813]), .x2814(x[2814]), .x2815(x[2815]), .x2816(x[2816]), .x2817(x[2817]), .x2818(x[2818]), .x2819(x[2819]), .x2820(x[2820]), .x2821(x[2821]), .x2822(x[2822]), .x2823(x[2823]), .x2824(x[2824]), .x2825(x[2825]), .x2826(x[2826]), .x2827(x[2827]), .x2828(x[2828]), .x2829(x[2829]), .x2830(x[2830]), .x2831(x[2831]), .x2832(x[2832]), .x2833(x[2833]), .x2834(x[2834]), .x2835(x[2835]), .x2836(x[2836]), .x2837(x[2837]), .x2838(x[2838]), .x2839(x[2839]), .x2840(x[2840]), .x2841(x[2841]), .x2842(x[2842]), .x2843(x[2843]), .x2844(x[2844]), .x2845(x[2845]), .x2846(x[2846]), .x2847(x[2847]), .x2848(x[2848]), .x2849(x[2849]), .x2850(x[2850]), .x2851(x[2851]), .x2852(x[2852]), .x2853(x[2853]), .x2854(x[2854]), .x2855(x[2855]), .x2856(x[2856]), .x2857(x[2857]), .x2858(x[2858]), .x2859(x[2859]), .x2860(x[2860]), .x2861(x[2861]), .x2862(x[2862]), .x2863(x[2863]), .x2864(x[2864]), .x2865(x[2865]), .x2866(x[2866]), .x2867(x[2867]), .x2868(x[2868]), .x2869(x[2869]), .x2870(x[2870]), .x2871(x[2871]), .x2872(x[2872]), .x2873(x[2873]), .x2874(x[2874]), .x2875(x[2875]), .x2876(x[2876]), .x2877(x[2877]), .x2878(x[2878]), .x2879(x[2879]), .x2880(x[2880]), .x2881(x[2881]), .x2882(x[2882]), .x2883(x[2883]), .x2884(x[2884]), .x2885(x[2885]), .x2886(x[2886]), .x2887(x[2887]), .x2888(x[2888]), .x2889(x[2889]), .x2890(x[2890]), .x2891(x[2891]), .x2892(x[2892]), .x2893(x[2893]), .x2894(x[2894]), .x2895(x[2895]), .x2896(x[2896]), .x2897(x[2897]), .x2898(x[2898]), .x2899(x[2899]), .x2900(x[2900]), .x2901(x[2901]), .x2902(x[2902]), .x2903(x[2903]), .x2904(x[2904]), .x2905(x[2905]), .x2906(x[2906]), .x2907(x[2907]), .x2908(x[2908]), .x2909(x[2909]), .x2910(x[2910]), .x2911(x[2911]), .x2912(x[2912]), .x2913(x[2913]), .x2914(x[2914]), .x2915(x[2915]), .x2916(x[2916]), .x2917(x[2917]), .x2918(x[2918]), .x2919(x[2919]), .x2920(x[2920]), .x2921(x[2921]), .x2922(x[2922]), .x2923(x[2923]), .x2924(x[2924]), .x2925(x[2925]), .x2926(x[2926]), .x2927(x[2927]), .x2928(x[2928]), .x2929(x[2929]), .x2930(x[2930]), .x2931(x[2931]), .x2932(x[2932]), .x2933(x[2933]), .x2934(x[2934]), .x2935(x[2935]), .x2936(x[2936]), .x2937(x[2937]), .x2938(x[2938]), .x2939(x[2939]), .x2940(x[2940]), .x2941(x[2941]), .x2942(x[2942]), .x2943(x[2943]), .x2944(x[2944]), .x2945(x[2945]), .x2946(x[2946]), .x2947(x[2947]), .x2948(x[2948]), .x2949(x[2949]), .x2950(x[2950]), .x2951(x[2951]), .x2952(x[2952]), .x2953(x[2953]), .x2954(x[2954]), .x2955(x[2955]), .x2956(x[2956]), .x2957(x[2957]), .x2958(x[2958]), .x2959(x[2959]), .x2960(x[2960]), .x2961(x[2961]), .x2962(x[2962]), .x2963(x[2963]), .x2964(x[2964]), .x2965(x[2965]), .x2966(x[2966]), .x2967(x[2967]), .x2968(x[2968]), .x2969(x[2969]), .x2970(x[2970]), .x2971(x[2971]), .x2972(x[2972]), .x2973(x[2973]), .x2974(x[2974]), .x2975(x[2975]), .x2976(x[2976]), .x2977(x[2977]), .x2978(x[2978]), .x2979(x[2979]), .x2980(x[2980]), .x2981(x[2981]), .x2982(x[2982]), .x2983(x[2983]), .x2984(x[2984]), .x2985(x[2985]), .x2986(x[2986]), .x2987(x[2987]), .x2988(x[2988]), .x2989(x[2989]), .x2990(x[2990]), .x2991(x[2991]), .x2992(x[2992]), .x2993(x[2993]), .x2994(x[2994]), .x2995(x[2995]), .x2996(x[2996]), .x2997(x[2997]), .x2998(x[2998]), .x2999(x[2999]), .x3000(x[3000]),
    .y0(y0)
  );

  // Optional reference function (majority reference for sanity check)
  function [11:0] popcount(input [3000:0] v);
    integer i; reg [11:0] c;
    begin
      c = 0;
      for (i = 0; i < 3001; i = i + 1)
        c = c + v[i];
      popcount = c;
    end
  endfunction

  // Reference majority: at least 1501 ones
  wire y_ref = (popcount(x) >= 1501);

  localparam [63:0] TOTAL_VECTORS = 64'd2460463844322234353863117626553505029281427791473667431532236058320117601229345897550720135677186919164859298508103609817025768361796473647170164964130696662469918700711690034826046640222721333845249456479513760832868956631387350026826181514417380753586593317621325883648986976903453010607425832010693495817247405346961838707873626211473240804705489553807680955767302200644818603966976727605861080964975819526968196507881457370264088817727469508542425184943557287898973377023442103123940865561494909647553616928361394206167723624368697131045480391593365244411023691024161104020620100511603178699291856002267490948441430027366827815085558127519667752202708470368490193340084321441258823163004742496016860894369684197220641160835984413324494657444244177027287367815340720418325307341282261873994004341001351002749447997532011655158601446506949781224500270343778349798159822583024799547744357038036459978752;

  initial begin
    $display("Time | x3000 x2999 x2998 x2997 x2996 x2995 x2994 x2993 x2992 x2991 x2990 x2989 x2988 x2987 x2986 x2985 x2984 x2983 x2982 x2981 x2980 x2979 x2978 x2977 x2976 x2975 x2974 x2973 x2972 x2971 x2970 x2969 x2968 x2967 x2966 x2965 x2964 x2963 x2962 x2961 x2960 x2959 x2958 x2957 x2956 x2955 x2954 x2953 x2952 x2951 x2950 x2949 x2948 x2947 x2946 x2945 x2944 x2943 x2942 x2941 x2940 x2939 x2938 x2937 x2936 x2935 x2934 x2933 x2932 x2931 x2930 x2929 x2928 x2927 x2926 x2925 x2924 x2923 x2922 x2921 x2920 x2919 x2918 x2917 x2916 x2915 x2914 x2913 x2912 x2911 x2910 x2909 x2908 x2907 x2906 x2905 x2904 x2903 x2902 x2901 x2900 x2899 x2898 x2897 x2896 x2895 x2894 x2893 x2892 x2891 x2890 x2889 x2888 x2887 x2886 x2885 x2884 x2883 x2882 x2881 x2880 x2879 x2878 x2877 x2876 x2875 x2874 x2873 x2872 x2871 x2870 x2869 x2868 x2867 x2866 x2865 x2864 x2863 x2862 x2861 x2860 x2859 x2858 x2857 x2856 x2855 x2854 x2853 x2852 x2851 x2850 x2849 x2848 x2847 x2846 x2845 x2844 x2843 x2842 x2841 x2840 x2839 x2838 x2837 x2836 x2835 x2834 x2833 x2832 x2831 x2830 x2829 x2828 x2827 x2826 x2825 x2824 x2823 x2822 x2821 x2820 x2819 x2818 x2817 x2816 x2815 x2814 x2813 x2812 x2811 x2810 x2809 x2808 x2807 x2806 x2805 x2804 x2803 x2802 x2801 x2800 x2799 x2798 x2797 x2796 x2795 x2794 x2793 x2792 x2791 x2790 x2789 x2788 x2787 x2786 x2785 x2784 x2783 x2782 x2781 x2780 x2779 x2778 x2777 x2776 x2775 x2774 x2773 x2772 x2771 x2770 x2769 x2768 x2767 x2766 x2765 x2764 x2763 x2762 x2761 x2760 x2759 x2758 x2757 x2756 x2755 x2754 x2753 x2752 x2751 x2750 x2749 x2748 x2747 x2746 x2745 x2744 x2743 x2742 x2741 x2740 x2739 x2738 x2737 x2736 x2735 x2734 x2733 x2732 x2731 x2730 x2729 x2728 x2727 x2726 x2725 x2724 x2723 x2722 x2721 x2720 x2719 x2718 x2717 x2716 x2715 x2714 x2713 x2712 x2711 x2710 x2709 x2708 x2707 x2706 x2705 x2704 x2703 x2702 x2701 x2700 x2699 x2698 x2697 x2696 x2695 x2694 x2693 x2692 x2691 x2690 x2689 x2688 x2687 x2686 x2685 x2684 x2683 x2682 x2681 x2680 x2679 x2678 x2677 x2676 x2675 x2674 x2673 x2672 x2671 x2670 x2669 x2668 x2667 x2666 x2665 x2664 x2663 x2662 x2661 x2660 x2659 x2658 x2657 x2656 x2655 x2654 x2653 x2652 x2651 x2650 x2649 x2648 x2647 x2646 x2645 x2644 x2643 x2642 x2641 x2640 x2639 x2638 x2637 x2636 x2635 x2634 x2633 x2632 x2631 x2630 x2629 x2628 x2627 x2626 x2625 x2624 x2623 x2622 x2621 x2620 x2619 x2618 x2617 x2616 x2615 x2614 x2613 x2612 x2611 x2610 x2609 x2608 x2607 x2606 x2605 x2604 x2603 x2602 x2601 x2600 x2599 x2598 x2597 x2596 x2595 x2594 x2593 x2592 x2591 x2590 x2589 x2588 x2587 x2586 x2585 x2584 x2583 x2582 x2581 x2580 x2579 x2578 x2577 x2576 x2575 x2574 x2573 x2572 x2571 x2570 x2569 x2568 x2567 x2566 x2565 x2564 x2563 x2562 x2561 x2560 x2559 x2558 x2557 x2556 x2555 x2554 x2553 x2552 x2551 x2550 x2549 x2548 x2547 x2546 x2545 x2544 x2543 x2542 x2541 x2540 x2539 x2538 x2537 x2536 x2535 x2534 x2533 x2532 x2531 x2530 x2529 x2528 x2527 x2526 x2525 x2524 x2523 x2522 x2521 x2520 x2519 x2518 x2517 x2516 x2515 x2514 x2513 x2512 x2511 x2510 x2509 x2508 x2507 x2506 x2505 x2504 x2503 x2502 x2501 x2500 x2499 x2498 x2497 x2496 x2495 x2494 x2493 x2492 x2491 x2490 x2489 x2488 x2487 x2486 x2485 x2484 x2483 x2482 x2481 x2480 x2479 x2478 x2477 x2476 x2475 x2474 x2473 x2472 x2471 x2470 x2469 x2468 x2467 x2466 x2465 x2464 x2463 x2462 x2461 x2460 x2459 x2458 x2457 x2456 x2455 x2454 x2453 x2452 x2451 x2450 x2449 x2448 x2447 x2446 x2445 x2444 x2443 x2442 x2441 x2440 x2439 x2438 x2437 x2436 x2435 x2434 x2433 x2432 x2431 x2430 x2429 x2428 x2427 x2426 x2425 x2424 x2423 x2422 x2421 x2420 x2419 x2418 x2417 x2416 x2415 x2414 x2413 x2412 x2411 x2410 x2409 x2408 x2407 x2406 x2405 x2404 x2403 x2402 x2401 x2400 x2399 x2398 x2397 x2396 x2395 x2394 x2393 x2392 x2391 x2390 x2389 x2388 x2387 x2386 x2385 x2384 x2383 x2382 x2381 x2380 x2379 x2378 x2377 x2376 x2375 x2374 x2373 x2372 x2371 x2370 x2369 x2368 x2367 x2366 x2365 x2364 x2363 x2362 x2361 x2360 x2359 x2358 x2357 x2356 x2355 x2354 x2353 x2352 x2351 x2350 x2349 x2348 x2347 x2346 x2345 x2344 x2343 x2342 x2341 x2340 x2339 x2338 x2337 x2336 x2335 x2334 x2333 x2332 x2331 x2330 x2329 x2328 x2327 x2326 x2325 x2324 x2323 x2322 x2321 x2320 x2319 x2318 x2317 x2316 x2315 x2314 x2313 x2312 x2311 x2310 x2309 x2308 x2307 x2306 x2305 x2304 x2303 x2302 x2301 x2300 x2299 x2298 x2297 x2296 x2295 x2294 x2293 x2292 x2291 x2290 x2289 x2288 x2287 x2286 x2285 x2284 x2283 x2282 x2281 x2280 x2279 x2278 x2277 x2276 x2275 x2274 x2273 x2272 x2271 x2270 x2269 x2268 x2267 x2266 x2265 x2264 x2263 x2262 x2261 x2260 x2259 x2258 x2257 x2256 x2255 x2254 x2253 x2252 x2251 x2250 x2249 x2248 x2247 x2246 x2245 x2244 x2243 x2242 x2241 x2240 x2239 x2238 x2237 x2236 x2235 x2234 x2233 x2232 x2231 x2230 x2229 x2228 x2227 x2226 x2225 x2224 x2223 x2222 x2221 x2220 x2219 x2218 x2217 x2216 x2215 x2214 x2213 x2212 x2211 x2210 x2209 x2208 x2207 x2206 x2205 x2204 x2203 x2202 x2201 x2200 x2199 x2198 x2197 x2196 x2195 x2194 x2193 x2192 x2191 x2190 x2189 x2188 x2187 x2186 x2185 x2184 x2183 x2182 x2181 x2180 x2179 x2178 x2177 x2176 x2175 x2174 x2173 x2172 x2171 x2170 x2169 x2168 x2167 x2166 x2165 x2164 x2163 x2162 x2161 x2160 x2159 x2158 x2157 x2156 x2155 x2154 x2153 x2152 x2151 x2150 x2149 x2148 x2147 x2146 x2145 x2144 x2143 x2142 x2141 x2140 x2139 x2138 x2137 x2136 x2135 x2134 x2133 x2132 x2131 x2130 x2129 x2128 x2127 x2126 x2125 x2124 x2123 x2122 x2121 x2120 x2119 x2118 x2117 x2116 x2115 x2114 x2113 x2112 x2111 x2110 x2109 x2108 x2107 x2106 x2105 x2104 x2103 x2102 x2101 x2100 x2099 x2098 x2097 x2096 x2095 x2094 x2093 x2092 x2091 x2090 x2089 x2088 x2087 x2086 x2085 x2084 x2083 x2082 x2081 x2080 x2079 x2078 x2077 x2076 x2075 x2074 x2073 x2072 x2071 x2070 x2069 x2068 x2067 x2066 x2065 x2064 x2063 x2062 x2061 x2060 x2059 x2058 x2057 x2056 x2055 x2054 x2053 x2052 x2051 x2050 x2049 x2048 x2047 x2046 x2045 x2044 x2043 x2042 x2041 x2040 x2039 x2038 x2037 x2036 x2035 x2034 x2033 x2032 x2031 x2030 x2029 x2028 x2027 x2026 x2025 x2024 x2023 x2022 x2021 x2020 x2019 x2018 x2017 x2016 x2015 x2014 x2013 x2012 x2011 x2010 x2009 x2008 x2007 x2006 x2005 x2004 x2003 x2002 x2001 x2000 x1999 x1998 x1997 x1996 x1995 x1994 x1993 x1992 x1991 x1990 x1989 x1988 x1987 x1986 x1985 x1984 x1983 x1982 x1981 x1980 x1979 x1978 x1977 x1976 x1975 x1974 x1973 x1972 x1971 x1970 x1969 x1968 x1967 x1966 x1965 x1964 x1963 x1962 x1961 x1960 x1959 x1958 x1957 x1956 x1955 x1954 x1953 x1952 x1951 x1950 x1949 x1948 x1947 x1946 x1945 x1944 x1943 x1942 x1941 x1940 x1939 x1938 x1937 x1936 x1935 x1934 x1933 x1932 x1931 x1930 x1929 x1928 x1927 x1926 x1925 x1924 x1923 x1922 x1921 x1920 x1919 x1918 x1917 x1916 x1915 x1914 x1913 x1912 x1911 x1910 x1909 x1908 x1907 x1906 x1905 x1904 x1903 x1902 x1901 x1900 x1899 x1898 x1897 x1896 x1895 x1894 x1893 x1892 x1891 x1890 x1889 x1888 x1887 x1886 x1885 x1884 x1883 x1882 x1881 x1880 x1879 x1878 x1877 x1876 x1875 x1874 x1873 x1872 x1871 x1870 x1869 x1868 x1867 x1866 x1865 x1864 x1863 x1862 x1861 x1860 x1859 x1858 x1857 x1856 x1855 x1854 x1853 x1852 x1851 x1850 x1849 x1848 x1847 x1846 x1845 x1844 x1843 x1842 x1841 x1840 x1839 x1838 x1837 x1836 x1835 x1834 x1833 x1832 x1831 x1830 x1829 x1828 x1827 x1826 x1825 x1824 x1823 x1822 x1821 x1820 x1819 x1818 x1817 x1816 x1815 x1814 x1813 x1812 x1811 x1810 x1809 x1808 x1807 x1806 x1805 x1804 x1803 x1802 x1801 x1800 x1799 x1798 x1797 x1796 x1795 x1794 x1793 x1792 x1791 x1790 x1789 x1788 x1787 x1786 x1785 x1784 x1783 x1782 x1781 x1780 x1779 x1778 x1777 x1776 x1775 x1774 x1773 x1772 x1771 x1770 x1769 x1768 x1767 x1766 x1765 x1764 x1763 x1762 x1761 x1760 x1759 x1758 x1757 x1756 x1755 x1754 x1753 x1752 x1751 x1750 x1749 x1748 x1747 x1746 x1745 x1744 x1743 x1742 x1741 x1740 x1739 x1738 x1737 x1736 x1735 x1734 x1733 x1732 x1731 x1730 x1729 x1728 x1727 x1726 x1725 x1724 x1723 x1722 x1721 x1720 x1719 x1718 x1717 x1716 x1715 x1714 x1713 x1712 x1711 x1710 x1709 x1708 x1707 x1706 x1705 x1704 x1703 x1702 x1701 x1700 x1699 x1698 x1697 x1696 x1695 x1694 x1693 x1692 x1691 x1690 x1689 x1688 x1687 x1686 x1685 x1684 x1683 x1682 x1681 x1680 x1679 x1678 x1677 x1676 x1675 x1674 x1673 x1672 x1671 x1670 x1669 x1668 x1667 x1666 x1665 x1664 x1663 x1662 x1661 x1660 x1659 x1658 x1657 x1656 x1655 x1654 x1653 x1652 x1651 x1650 x1649 x1648 x1647 x1646 x1645 x1644 x1643 x1642 x1641 x1640 x1639 x1638 x1637 x1636 x1635 x1634 x1633 x1632 x1631 x1630 x1629 x1628 x1627 x1626 x1625 x1624 x1623 x1622 x1621 x1620 x1619 x1618 x1617 x1616 x1615 x1614 x1613 x1612 x1611 x1610 x1609 x1608 x1607 x1606 x1605 x1604 x1603 x1602 x1601 x1600 x1599 x1598 x1597 x1596 x1595 x1594 x1593 x1592 x1591 x1590 x1589 x1588 x1587 x1586 x1585 x1584 x1583 x1582 x1581 x1580 x1579 x1578 x1577 x1576 x1575 x1574 x1573 x1572 x1571 x1570 x1569 x1568 x1567 x1566 x1565 x1564 x1563 x1562 x1561 x1560 x1559 x1558 x1557 x1556 x1555 x1554 x1553 x1552 x1551 x1550 x1549 x1548 x1547 x1546 x1545 x1544 x1543 x1542 x1541 x1540 x1539 x1538 x1537 x1536 x1535 x1534 x1533 x1532 x1531 x1530 x1529 x1528 x1527 x1526 x1525 x1524 x1523 x1522 x1521 x1520 x1519 x1518 x1517 x1516 x1515 x1514 x1513 x1512 x1511 x1510 x1509 x1508 x1507 x1506 x1505 x1504 x1503 x1502 x1501 x1500 x1499 x1498 x1497 x1496 x1495 x1494 x1493 x1492 x1491 x1490 x1489 x1488 x1487 x1486 x1485 x1484 x1483 x1482 x1481 x1480 x1479 x1478 x1477 x1476 x1475 x1474 x1473 x1472 x1471 x1470 x1469 x1468 x1467 x1466 x1465 x1464 x1463 x1462 x1461 x1460 x1459 x1458 x1457 x1456 x1455 x1454 x1453 x1452 x1451 x1450 x1449 x1448 x1447 x1446 x1445 x1444 x1443 x1442 x1441 x1440 x1439 x1438 x1437 x1436 x1435 x1434 x1433 x1432 x1431 x1430 x1429 x1428 x1427 x1426 x1425 x1424 x1423 x1422 x1421 x1420 x1419 x1418 x1417 x1416 x1415 x1414 x1413 x1412 x1411 x1410 x1409 x1408 x1407 x1406 x1405 x1404 x1403 x1402 x1401 x1400 x1399 x1398 x1397 x1396 x1395 x1394 x1393 x1392 x1391 x1390 x1389 x1388 x1387 x1386 x1385 x1384 x1383 x1382 x1381 x1380 x1379 x1378 x1377 x1376 x1375 x1374 x1373 x1372 x1371 x1370 x1369 x1368 x1367 x1366 x1365 x1364 x1363 x1362 x1361 x1360 x1359 x1358 x1357 x1356 x1355 x1354 x1353 x1352 x1351 x1350 x1349 x1348 x1347 x1346 x1345 x1344 x1343 x1342 x1341 x1340 x1339 x1338 x1337 x1336 x1335 x1334 x1333 x1332 x1331 x1330 x1329 x1328 x1327 x1326 x1325 x1324 x1323 x1322 x1321 x1320 x1319 x1318 x1317 x1316 x1315 x1314 x1313 x1312 x1311 x1310 x1309 x1308 x1307 x1306 x1305 x1304 x1303 x1302 x1301 x1300 x1299 x1298 x1297 x1296 x1295 x1294 x1293 x1292 x1291 x1290 x1289 x1288 x1287 x1286 x1285 x1284 x1283 x1282 x1281 x1280 x1279 x1278 x1277 x1276 x1275 x1274 x1273 x1272 x1271 x1270 x1269 x1268 x1267 x1266 x1265 x1264 x1263 x1262 x1261 x1260 x1259 x1258 x1257 x1256 x1255 x1254 x1253 x1252 x1251 x1250 x1249 x1248 x1247 x1246 x1245 x1244 x1243 x1242 x1241 x1240 x1239 x1238 x1237 x1236 x1235 x1234 x1233 x1232 x1231 x1230 x1229 x1228 x1227 x1226 x1225 x1224 x1223 x1222 x1221 x1220 x1219 x1218 x1217 x1216 x1215 x1214 x1213 x1212 x1211 x1210 x1209 x1208 x1207 x1206 x1205 x1204 x1203 x1202 x1201 x1200 x1199 x1198 x1197 x1196 x1195 x1194 x1193 x1192 x1191 x1190 x1189 x1188 x1187 x1186 x1185 x1184 x1183 x1182 x1181 x1180 x1179 x1178 x1177 x1176 x1175 x1174 x1173 x1172 x1171 x1170 x1169 x1168 x1167 x1166 x1165 x1164 x1163 x1162 x1161 x1160 x1159 x1158 x1157 x1156 x1155 x1154 x1153 x1152 x1151 x1150 x1149 x1148 x1147 x1146 x1145 x1144 x1143 x1142 x1141 x1140 x1139 x1138 x1137 x1136 x1135 x1134 x1133 x1132 x1131 x1130 x1129 x1128 x1127 x1126 x1125 x1124 x1123 x1122 x1121 x1120 x1119 x1118 x1117 x1116 x1115 x1114 x1113 x1112 x1111 x1110 x1109 x1108 x1107 x1106 x1105 x1104 x1103 x1102 x1101 x1100 x1099 x1098 x1097 x1096 x1095 x1094 x1093 x1092 x1091 x1090 x1089 x1088 x1087 x1086 x1085 x1084 x1083 x1082 x1081 x1080 x1079 x1078 x1077 x1076 x1075 x1074 x1073 x1072 x1071 x1070 x1069 x1068 x1067 x1066 x1065 x1064 x1063 x1062 x1061 x1060 x1059 x1058 x1057 x1056 x1055 x1054 x1053 x1052 x1051 x1050 x1049 x1048 x1047 x1046 x1045 x1044 x1043 x1042 x1041 x1040 x1039 x1038 x1037 x1036 x1035 x1034 x1033 x1032 x1031 x1030 x1029 x1028 x1027 x1026 x1025 x1024 x1023 x1022 x1021 x1020 x1019 x1018 x1017 x1016 x1015 x1014 x1013 x1012 x1011 x1010 x1009 x1008 x1007 x1006 x1005 x1004 x1003 x1002 x1001 x1000 x999 x998 x997 x996 x995 x994 x993 x992 x991 x990 x989 x988 x987 x986 x985 x984 x983 x982 x981 x980 x979 x978 x977 x976 x975 x974 x973 x972 x971 x970 x969 x968 x967 x966 x965 x964 x963 x962 x961 x960 x959 x958 x957 x956 x955 x954 x953 x952 x951 x950 x949 x948 x947 x946 x945 x944 x943 x942 x941 x940 x939 x938 x937 x936 x935 x934 x933 x932 x931 x930 x929 x928 x927 x926 x925 x924 x923 x922 x921 x920 x919 x918 x917 x916 x915 x914 x913 x912 x911 x910 x909 x908 x907 x906 x905 x904 x903 x902 x901 x900 x899 x898 x897 x896 x895 x894 x893 x892 x891 x890 x889 x888 x887 x886 x885 x884 x883 x882 x881 x880 x879 x878 x877 x876 x875 x874 x873 x872 x871 x870 x869 x868 x867 x866 x865 x864 x863 x862 x861 x860 x859 x858 x857 x856 x855 x854 x853 x852 x851 x850 x849 x848 x847 x846 x845 x844 x843 x842 x841 x840 x839 x838 x837 x836 x835 x834 x833 x832 x831 x830 x829 x828 x827 x826 x825 x824 x823 x822 x821 x820 x819 x818 x817 x816 x815 x814 x813 x812 x811 x810 x809 x808 x807 x806 x805 x804 x803 x802 x801 x800 x799 x798 x797 x796 x795 x794 x793 x792 x791 x790 x789 x788 x787 x786 x785 x784 x783 x782 x781 x780 x779 x778 x777 x776 x775 x774 x773 x772 x771 x770 x769 x768 x767 x766 x765 x764 x763 x762 x761 x760 x759 x758 x757 x756 x755 x754 x753 x752 x751 x750 x749 x748 x747 x746 x745 x744 x743 x742 x741 x740 x739 x738 x737 x736 x735 x734 x733 x732 x731 x730 x729 x728 x727 x726 x725 x724 x723 x722 x721 x720 x719 x718 x717 x716 x715 x714 x713 x712 x711 x710 x709 x708 x707 x706 x705 x704 x703 x702 x701 x700 x699 x698 x697 x696 x695 x694 x693 x692 x691 x690 x689 x688 x687 x686 x685 x684 x683 x682 x681 x680 x679 x678 x677 x676 x675 x674 x673 x672 x671 x670 x669 x668 x667 x666 x665 x664 x663 x662 x661 x660 x659 x658 x657 x656 x655 x654 x653 x652 x651 x650 x649 x648 x647 x646 x645 x644 x643 x642 x641 x640 x639 x638 x637 x636 x635 x634 x633 x632 x631 x630 x629 x628 x627 x626 x625 x624 x623 x622 x621 x620 x619 x618 x617 x616 x615 x614 x613 x612 x611 x610 x609 x608 x607 x606 x605 x604 x603 x602 x601 x600 x599 x598 x597 x596 x595 x594 x593 x592 x591 x590 x589 x588 x587 x586 x585 x584 x583 x582 x581 x580 x579 x578 x577 x576 x575 x574 x573 x572 x571 x570 x569 x568 x567 x566 x565 x564 x563 x562 x561 x560 x559 x558 x557 x556 x555 x554 x553 x552 x551 x550 x549 x548 x547 x546 x545 x544 x543 x542 x541 x540 x539 x538 x537 x536 x535 x534 x533 x532 x531 x530 x529 x528 x527 x526 x525 x524 x523 x522 x521 x520 x519 x518 x517 x516 x515 x514 x513 x512 x511 x510 x509 x508 x507 x506 x505 x504 x503 x502 x501 x500 x499 x498 x497 x496 x495 x494 x493 x492 x491 x490 x489 x488 x487 x486 x485 x484 x483 x482 x481 x480 x479 x478 x477 x476 x475 x474 x473 x472 x471 x470 x469 x468 x467 x466 x465 x464 x463 x462 x461 x460 x459 x458 x457 x456 x455 x454 x453 x452 x451 x450 x449 x448 x447 x446 x445 x444 x443 x442 x441 x440 x439 x438 x437 x436 x435 x434 x433 x432 x431 x430 x429 x428 x427 x426 x425 x424 x423 x422 x421 x420 x419 x418 x417 x416 x415 x414 x413 x412 x411 x410 x409 x408 x407 x406 x405 x404 x403 x402 x401 x400 x399 x398 x397 x396 x395 x394 x393 x392 x391 x390 x389 x388 x387 x386 x385 x384 x383 x382 x381 x380 x379 x378 x377 x376 x375 x374 x373 x372 x371 x370 x369 x368 x367 x366 x365 x364 x363 x362 x361 x360 x359 x358 x357 x356 x355 x354 x353 x352 x351 x350 x349 x348 x347 x346 x345 x344 x343 x342 x341 x340 x339 x338 x337 x336 x335 x334 x333 x332 x331 x330 x329 x328 x327 x326 x325 x324 x323 x322 x321 x320 x319 x318 x317 x316 x315 x314 x313 x312 x311 x310 x309 x308 x307 x306 x305 x304 x303 x302 x301 x300 x299 x298 x297 x296 x295 x294 x293 x292 x291 x290 x289 x288 x287 x286 x285 x284 x283 x282 x281 x280 x279 x278 x277 x276 x275 x274 x273 x272 x271 x270 x269 x268 x267 x266 x265 x264 x263 x262 x261 x260 x259 x258 x257 x256 x255 x254 x253 x252 x251 x250 x249 x248 x247 x246 x245 x244 x243 x242 x241 x240 x239 x238 x237 x236 x235 x234 x233 x232 x231 x230 x229 x228 x227 x226 x225 x224 x223 x222 x221 x220 x219 x218 x217 x216 x215 x214 x213 x212 x211 x210 x209 x208 x207 x206 x205 x204 x203 x202 x201 x200 x199 x198 x197 x196 x195 x194 x193 x192 x191 x190 x189 x188 x187 x186 x185 x184 x183 x182 x181 x180 x179 x178 x177 x176 x175 x174 x173 x172 x171 x170 x169 x168 x167 x166 x165 x164 x163 x162 x161 x160 x159 x158 x157 x156 x155 x154 x153 x152 x151 x150 x149 x148 x147 x146 x145 x144 x143 x142 x141 x140 x139 x138 x137 x136 x135 x134 x133 x132 x131 x130 x129 x128 x127 x126 x125 x124 x123 x122 x121 x120 x119 x118 x117 x116 x115 x114 x113 x112 x111 x110 x109 x108 x107 x106 x105 x104 x103 x102 x101 x100 x99 x98 x97 x96 x95 x94 x93 x92 x91 x90 x89 x88 x87 x86 x85 x84 x83 x82 x81 x80 x79 x78 x77 x76 x75 x74 x73 x72 x71 x70 x69 x68 x67 x66 x65 x64 x63 x62 x61 x60 x59 x58 x57 x56 x55 x54 x53 x52 x51 x50 x49 x48 x47 x46 x45 x44 x43 x42 x41 x40 x39 x38 x37 x36 x35 x34 x33 x32 x31 x30 x29 x28 x27 x26 x25 x24 x23 x22 x21 x20 x19 x18 x17 x16 x15 x14 x13 x12 x11 x10 x9 x8 x7 x6 x5 x4 x3 x2 x1 x0 | y0 (DUT) y_ref (Maj3001)");
    $display("---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------");
    // Loop through all 2460463844322234353863117626553505029281427791473667431532236058320117601229345897550720135677186919164859298508103609817025768361796473647170164964130696662469918700711690034826046640222721333845249456479513760832868956631387350026826181514417380753586593317621325883648986976903453010607425832010693495817247405346961838707873626211473240804705489553807680955767302200644818603966976727605861080964975819526968196507881457370264088817727469508542425184943557287898973377023442103123940865561494909647553616928361394206167723624368697131045480391593365244411023691024161104020620100511603178699291856002267490948441430027366827815085558127519667752202708470368490193340084321441258823163004742496016860894369684197220641160835984413324494657444244177027287367815340720418325307341282261873994004341001351002749447997532011655158601446506949781224500270343778349798159822583024799547744357038036459978752 combinations
    for (idx = 0; idx < TOTAL_VECTORS; idx = idx + 1) begin
      x = idx[3000:0];
      #10 $display("%4t |  %b  |   %b       %b",
                   $time, x, y0, y_ref);
    end
    #10 $finish;
  end

  // Optional mismatch check
  always #1 if (^x !== 1'bx && y0 !== y_ref)
    $display("Mismatch at t=%0t x=%b HW=%0d y0=%0b ref=%0b",
             $time, x, popcount(x), y0, y_ref);

endmodule

`default_nettype wire
