module top (x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, y0);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58;
  output y0;
  wire n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n136, n137, n135, n138, n139, n140, n141;
  LUT3 #(.INIT(8'hE8)) lut_n61 (.I0(x0), .I1(x1), .I2(x2), .O(n61));
  LUT3 #(.INIT(8'hE8)) lut_n62 (.I0(x6), .I1(x7), .I2(x8), .O(n62));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n63 (.I0(x3), .I1(x4), .I2(x5), .I3(n61), .I4(n62), .O(n63));
  LUT3 #(.INIT(8'hE8)) lut_n64 (.I0(x12), .I1(x13), .I2(x14), .O(n64));
  LUT5 #(.INIT(32'hE81717E8)) lut_n65 (.I0(x3), .I1(x4), .I2(x5), .I3(n61), .I4(n62), .O(n65));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n66 (.I0(x9), .I1(x10), .I2(x11), .I3(n64), .I4(n65), .O(n66));
  LUT3 #(.INIT(8'hE8)) lut_n67 (.I0(x18), .I1(x19), .I2(x20), .O(n67));
  LUT5 #(.INIT(32'hE81717E8)) lut_n68 (.I0(x9), .I1(x10), .I2(x11), .I3(n64), .I4(n65), .O(n68));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n69 (.I0(x15), .I1(x16), .I2(x17), .I3(n67), .I4(n68), .O(n69));
  LUT3 #(.INIT(8'hE8)) lut_n70 (.I0(n63), .I1(n66), .I2(n69), .O(n70));
  LUT3 #(.INIT(8'hE8)) lut_n71 (.I0(x24), .I1(x25), .I2(x26), .O(n71));
  LUT5 #(.INIT(32'hE81717E8)) lut_n72 (.I0(x15), .I1(x16), .I2(x17), .I3(n67), .I4(n68), .O(n72));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n73 (.I0(x21), .I1(x22), .I2(x23), .I3(n71), .I4(n72), .O(n73));
  LUT3 #(.INIT(8'hE8)) lut_n74 (.I0(x27), .I1(x28), .I2(x29), .O(n74));
  LUT5 #(.INIT(32'hE81717E8)) lut_n75 (.I0(x21), .I1(x22), .I2(x23), .I3(n71), .I4(n72), .O(n75));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n76 (.I0(x30), .I1(x31), .I2(x32), .I3(n74), .I4(n75), .O(n76));
  LUT3 #(.INIT(8'h96)) lut_n77 (.I0(n63), .I1(n66), .I2(n69), .O(n77));
  LUT3 #(.INIT(8'hE8)) lut_n78 (.I0(n73), .I1(n76), .I2(n77), .O(n78));
  LUT3 #(.INIT(8'hE8)) lut_n79 (.I0(x36), .I1(x37), .I2(x38), .O(n79));
  LUT5 #(.INIT(32'hE81717E8)) lut_n80 (.I0(x30), .I1(x31), .I2(x32), .I3(n74), .I4(n75), .O(n80));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n81 (.I0(x33), .I1(x34), .I2(x35), .I3(n79), .I4(n80), .O(n81));
  LUT3 #(.INIT(8'hE8)) lut_n82 (.I0(x42), .I1(x43), .I2(x44), .O(n82));
  LUT5 #(.INIT(32'hE81717E8)) lut_n83 (.I0(x33), .I1(x34), .I2(x35), .I3(n79), .I4(n80), .O(n83));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n84 (.I0(x39), .I1(x40), .I2(x41), .I3(n82), .I4(n83), .O(n84));
  LUT3 #(.INIT(8'h96)) lut_n85 (.I0(n73), .I1(n76), .I2(n77), .O(n85));
  LUT3 #(.INIT(8'hE8)) lut_n86 (.I0(n81), .I1(n84), .I2(n85), .O(n86));
  LUT3 #(.INIT(8'hE8)) lut_n87 (.I0(n70), .I1(n78), .I2(n86), .O(n87));
  LUT3 #(.INIT(8'hE8)) lut_n88 (.I0(x48), .I1(x49), .I2(x50), .O(n88));
  LUT5 #(.INIT(32'hE81717E8)) lut_n89 (.I0(x39), .I1(x40), .I2(x41), .I3(n82), .I4(n83), .O(n89));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n90 (.I0(x45), .I1(x46), .I2(x47), .I3(n88), .I4(n89), .O(n90));
  LUT3 #(.INIT(8'hE8)) lut_n91 (.I0(x54), .I1(x55), .I2(x56), .O(n91));
  LUT5 #(.INIT(32'hE81717E8)) lut_n92 (.I0(x45), .I1(x46), .I2(x47), .I3(n88), .I4(n89), .O(n92));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n93 (.I0(x51), .I1(x52), .I2(x53), .I3(n91), .I4(n92), .O(n93));
  LUT3 #(.INIT(8'h96)) lut_n94 (.I0(n81), .I1(n84), .I2(n85), .O(n94));
  LUT3 #(.INIT(8'hE8)) lut_n95 (.I0(n90), .I1(n93), .I2(n94), .O(n95));
  LUT5 #(.INIT(32'hE81717E8)) lut_n96 (.I0(x51), .I1(x52), .I2(x53), .I3(n91), .I4(n92), .O(n96));
  LUT3 #(.INIT(8'hE0)) lut_n97 (.I0(x57), .I1(x58), .I2(n96), .O(n97));
  LUT3 #(.INIT(8'h96)) lut_n98 (.I0(x0), .I1(x1), .I2(x2), .O(n98));
  LUT3 #(.INIT(8'h96)) lut_n99 (.I0(x6), .I1(x7), .I2(x8), .O(n99));
  LUT5 #(.INIT(32'hFF969600)) lut_n100 (.I0(x3), .I1(x4), .I2(x5), .I3(n98), .I4(n99), .O(n100));
  LUT3 #(.INIT(8'h96)) lut_n101 (.I0(x12), .I1(x13), .I2(x14), .O(n101));
  LUT5 #(.INIT(32'h96696996)) lut_n102 (.I0(x3), .I1(x4), .I2(x5), .I3(n98), .I4(n99), .O(n102));
  LUT5 #(.INIT(32'hFF969600)) lut_n103 (.I0(x9), .I1(x10), .I2(x11), .I3(n101), .I4(n102), .O(n103));
  LUT3 #(.INIT(8'h1E)) lut_n104 (.I0(x57), .I1(x58), .I2(n96), .O(n104));
  LUT3 #(.INIT(8'hE8)) lut_n105 (.I0(n100), .I1(n103), .I2(n104), .O(n105));
  LUT3 #(.INIT(8'h96)) lut_n106 (.I0(n90), .I1(n93), .I2(n94), .O(n106));
  LUT3 #(.INIT(8'hE8)) lut_n107 (.I0(n97), .I1(n105), .I2(n106), .O(n107));
  LUT3 #(.INIT(8'h96)) lut_n108 (.I0(n70), .I1(n78), .I2(n86), .O(n108));
  LUT3 #(.INIT(8'h96)) lut_n109 (.I0(x18), .I1(x19), .I2(x20), .O(n109));
  LUT5 #(.INIT(32'h96696996)) lut_n110 (.I0(x9), .I1(x10), .I2(x11), .I3(n101), .I4(n102), .O(n110));
  LUT5 #(.INIT(32'hFF969600)) lut_n111 (.I0(x15), .I1(x16), .I2(x17), .I3(n109), .I4(n110), .O(n111));
  LUT3 #(.INIT(8'h96)) lut_n112 (.I0(x24), .I1(x25), .I2(x26), .O(n112));
  LUT5 #(.INIT(32'h96696996)) lut_n113 (.I0(x15), .I1(x16), .I2(x17), .I3(n109), .I4(n110), .O(n113));
  LUT5 #(.INIT(32'hFF969600)) lut_n114 (.I0(x21), .I1(x22), .I2(x23), .I3(n112), .I4(n113), .O(n114));
  LUT3 #(.INIT(8'h96)) lut_n115 (.I0(n100), .I1(n103), .I2(n104), .O(n115));
  LUT3 #(.INIT(8'hE8)) lut_n116 (.I0(n111), .I1(n114), .I2(n115), .O(n116));
  LUT3 #(.INIT(8'h96)) lut_n117 (.I0(x27), .I1(x28), .I2(x29), .O(n117));
  LUT5 #(.INIT(32'h96696996)) lut_n118 (.I0(x21), .I1(x22), .I2(x23), .I3(n112), .I4(n113), .O(n118));
  LUT5 #(.INIT(32'hFF969600)) lut_n119 (.I0(x30), .I1(x31), .I2(x32), .I3(n117), .I4(n118), .O(n119));
  LUT3 #(.INIT(8'h96)) lut_n120 (.I0(x36), .I1(x37), .I2(x38), .O(n120));
  LUT5 #(.INIT(32'h96696996)) lut_n121 (.I0(x30), .I1(x31), .I2(x32), .I3(n117), .I4(n118), .O(n121));
  LUT5 #(.INIT(32'hFF969600)) lut_n122 (.I0(x33), .I1(x34), .I2(x35), .I3(n120), .I4(n121), .O(n122));
  LUT3 #(.INIT(8'h96)) lut_n123 (.I0(n111), .I1(n114), .I2(n115), .O(n123));
  LUT3 #(.INIT(8'hE8)) lut_n124 (.I0(n119), .I1(n122), .I2(n123), .O(n124));
  LUT3 #(.INIT(8'h96)) lut_n125 (.I0(n97), .I1(n105), .I2(n106), .O(n125));
  LUT3 #(.INIT(8'hE8)) lut_n126 (.I0(n116), .I1(n124), .I2(n125), .O(n126));
  LUT3 #(.INIT(8'h96)) lut_n127 (.I0(x42), .I1(x43), .I2(x44), .O(n127));
  LUT5 #(.INIT(32'h96696996)) lut_n128 (.I0(x33), .I1(x34), .I2(x35), .I3(n120), .I4(n121), .O(n128));
  LUT5 #(.INIT(32'hFF969600)) lut_n129 (.I0(x39), .I1(x40), .I2(x41), .I3(n127), .I4(n128), .O(n129));
  LUT3 #(.INIT(8'h96)) lut_n130 (.I0(x48), .I1(x49), .I2(x50), .O(n130));
  LUT5 #(.INIT(32'h96696996)) lut_n131 (.I0(x39), .I1(x40), .I2(x41), .I3(n127), .I4(n128), .O(n131));
  LUT5 #(.INIT(32'hFF969600)) lut_n132 (.I0(x45), .I1(x46), .I2(x47), .I3(n130), .I4(n131), .O(n132));
  LUT3 #(.INIT(8'h96)) lut_n133 (.I0(n119), .I1(n122), .I2(n123), .O(n133));
  LUT3 #(.INIT(8'h96)) lut_n134 (.I0(x51), .I1(x52), .I2(x53), .O(n134));
  LUT5 #(.INIT(32'h96696996)) lut_n136 (.I0(x45), .I1(x46), .I2(x47), .I3(n130), .I4(n131), .O(n136));
  LUT5 #(.INIT(32'hFF969600)) lut_n137 (.I0(x54), .I1(x55), .I2(x56), .I3(n134), .I4(n136), .O(n137));
  LUT3 #(.INIT(8'h96)) lut_n135 (.I0(x54), .I1(x55), .I2(x56), .O(n135));
  LUT5 #(.INIT(32'h06606006)) lut_n138 (.I0(x57), .I1(x58), .I2(n134), .I3(n135), .I4(n136), .O(n138));
  LUT3 #(.INIT(8'h96)) lut_n139 (.I0(n116), .I1(n124), .I2(n125), .O(n139));
  LUT6 #(.INIT(64'hFEE8FFFE8000E880)) lut_n140 (.I0(n129), .I1(n132), .I2(n133), .I3(n137), .I4(n138), .I5(n139), .O(n140));
  LUT6 #(.INIT(64'hFEEAEAA8EAA8A880)) lut_n141 (.I0(n87), .I1(n95), .I2(n107), .I3(n108), .I4(n126), .I5(n140), .O(n141));
  assign y0 = n141;
endmodule
