module top (x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255, x256, x257, x258, x259, x260, x261, x262, x263, x264, x265, x266, x267, x268, x269, x270, x271, x272, x273, x274, x275, x276, x277, x278, x279, x280, x281, x282, x283, x284, x285, x286, x287, x288, x289, x290, x291, x292, x293, x294, x295, x296, x297, x298, x299, x300, x301, x302, x303, x304, x305, x306, x307, x308, x309, x310, x311, x312, x313, x314, x315, x316, x317, x318, x319, x320, x321, x322, x323, x324, x325, x326, x327, x328, x329, x330, x331, x332, x333, x334, x335, x336, x337, x338, x339, x340, x341, x342, x343, x344, x345, x346, x347, x348, x349, x350, x351, x352, x353, x354, x355, x356, x357, x358, x359, x360, x361, x362, x363, x364, x365, x366, x367, x368, x369, x370, x371, x372, x373, x374, x375, x376, x377, x378, x379, x380, x381, x382, x383, x384, x385, x386, x387, x388, x389, x390, x391, x392, x393, x394, x395, x396, x397, x398, x399, x400, x401, x402, x403, x404, x405, x406, x407, x408, x409, x410, x411, x412, x413, x414, x415, x416, x417, x418, x419, x420, x421, x422, x423, x424, x425, x426, x427, x428, x429, x430, x431, x432, x433, x434, x435, x436, x437, x438, x439, x440, x441, x442, x443, x444, x445, x446, x447, x448, x449, x450, x451, x452, x453, x454, x455, x456, x457, x458, x459, x460, x461, x462, x463, x464, x465, x466, x467, x468, x469, x470, x471, x472, x473, x474, x475, x476, x477, x478, x479, x480, x481, x482, x483, x484, x485, x486, x487, x488, x489, x490, x491, x492, x493, x494, x495, x496, x497, x498, x499, x500, x501, x502, x503, x504, x505, x506, x507, x508, x509, x510, x511, x512, x513, x514, x515, x516, x517, x518, x519, x520, x521, x522, x523, x524, x525, x526, x527, x528, x529, x530, x531, x532, x533, x534, x535, x536, x537, x538, x539, x540, x541, x542, x543, x544, x545, x546, x547, x548, x549, x550, x551, x552, x553, x554, x555, x556, x557, x558, x559, x560, x561, x562, x563, x564, x565, x566, x567, x568, x569, x570, x571, x572, x573, x574, x575, x576, x577, x578, x579, x580, x581, x582, x583, x584, x585, x586, x587, x588, x589, x590, x591, x592, x593, x594, x595, x596, x597, x598, x599, x600, x601, x602, x603, x604, x605, x606, x607, x608, x609, x610, x611, x612, x613, x614, x615, x616, x617, x618, x619, x620, x621, x622, x623, x624, x625, x626, x627, x628, x629, x630, x631, x632, x633, x634, x635, x636, x637, x638, x639, x640, x641, x642, x643, x644, x645, x646, x647, x648, x649, x650, x651, x652, x653, x654, x655, x656, x657, x658, x659, x660, x661, x662, x663, x664, x665, x666, x667, x668, x669, x670, x671, x672, x673, x674, x675, x676, x677, x678, x679, x680, x681, x682, x683, x684, x685, x686, x687, x688, x689, x690, x691, x692, x693, x694, x695, x696, x697, x698, x699, x700, x701, x702, x703, x704, x705, x706, x707, x708, x709, x710, x711, x712, x713, x714, x715, x716, x717, x718, x719, x720, x721, x722, x723, x724, x725, x726, x727, x728, x729, x730, x731, x732, x733, x734, x735, x736, x737, x738, x739, x740, x741, x742, x743, x744, x745, x746, x747, x748, x749, x750, x751, x752, x753, x754, x755, x756, x757, x758, x759, x760, x761, x762, x763, x764, x765, x766, x767, x768, x769, x770, x771, x772, x773, x774, x775, x776, x777, x778, x779, x780, x781, x782, x783, x784, x785, x786, x787, x788, x789, x790, x791, x792, x793, x794, x795, x796, x797, x798, x799, x800, x801, x802, x803, x804, x805, x806, x807, x808, x809, x810, x811, x812, x813, x814, x815, x816, x817, x818, x819, x820, x821, x822, x823, x824, x825, x826, x827, x828, x829, x830, x831, x832, x833, x834, x835, x836, x837, x838, x839, x840, x841, x842, x843, x844, x845, x846, x847, x848, x849, x850, x851, x852, x853, x854, x855, x856, x857, x858, x859, x860, x861, x862, x863, x864, x865, x866, x867, x868, x869, x870, x871, x872, x873, x874, x875, x876, x877, x878, x879, x880, x881, x882, x883, x884, x885, x886, x887, x888, x889, x890, x891, x892, x893, x894, x895, x896, x897, x898, x899, x900, x901, x902, x903, x904, x905, x906, x907, x908, x909, x910, x911, x912, x913, x914, x915, x916, x917, x918, x919, x920, x921, x922, x923, x924, x925, x926, x927, x928, x929, x930, x931, x932, x933, x934, x935, x936, x937, x938, x939, x940, x941, x942, x943, x944, x945, x946, x947, x948, x949, x950, x951, x952, x953, x954, x955, x956, x957, x958, x959, x960, x961, x962, x963, x964, x965, x966, x967, x968, x969, x970, x971, x972, x973, x974, x975, x976, x977, x978, x979, x980, x981, x982, x983, x984, x985, x986, x987, x988, x989, x990, x991, x992, x993, x994, x995, x996, x997, x998, x999, x1000, x1001, x1002, x1003, x1004, x1005, x1006, x1007, x1008, x1009, x1010, x1011, x1012, x1013, x1014, x1015, x1016, x1017, x1018, x1019, x1020, x1021, x1022, x1023, x1024, x1025, x1026, x1027, x1028, x1029, x1030, x1031, x1032, x1033, x1034, x1035, x1036, x1037, x1038, x1039, x1040, x1041, x1042, x1043, x1044, x1045, x1046, x1047, x1048, x1049, x1050, x1051, x1052, x1053, x1054, x1055, x1056, x1057, x1058, x1059, x1060, x1061, x1062, x1063, x1064, x1065, x1066, x1067, x1068, x1069, x1070, x1071, x1072, x1073, x1074, x1075, x1076, x1077, x1078, x1079, x1080, x1081, x1082, x1083, x1084, x1085, x1086, x1087, x1088, x1089, x1090, x1091, x1092, x1093, x1094, x1095, x1096, x1097, x1098, x1099, x1100, x1101, x1102, x1103, x1104, x1105, x1106, x1107, x1108, x1109, x1110, x1111, x1112, x1113, x1114, x1115, x1116, x1117, x1118, x1119, x1120, x1121, x1122, x1123, x1124, x1125, x1126, x1127, x1128, x1129, x1130, x1131, x1132, x1133, x1134, x1135, x1136, x1137, x1138, x1139, x1140, x1141, x1142, x1143, x1144, x1145, x1146, x1147, x1148, x1149, x1150, x1151, x1152, x1153, x1154, x1155, x1156, x1157, x1158, x1159, x1160, x1161, x1162, x1163, x1164, x1165, x1166, x1167, x1168, x1169, x1170, x1171, x1172, x1173, x1174, x1175, x1176, x1177, x1178, x1179, x1180, x1181, x1182, x1183, x1184, x1185, x1186, x1187, x1188, x1189, x1190, x1191, x1192, x1193, x1194, x1195, x1196, x1197, x1198, x1199, x1200, x1201, x1202, x1203, x1204, x1205, x1206, x1207, x1208, x1209, x1210, x1211, x1212, x1213, x1214, x1215, x1216, x1217, x1218, x1219, x1220, x1221, x1222, x1223, x1224, x1225, x1226, x1227, x1228, x1229, x1230, x1231, x1232, x1233, x1234, x1235, x1236, x1237, x1238, x1239, x1240, x1241, x1242, x1243, x1244, x1245, x1246, x1247, x1248, x1249, x1250, x1251, x1252, x1253, x1254, x1255, x1256, x1257, x1258, x1259, x1260, x1261, x1262, x1263, x1264, x1265, x1266, x1267, x1268, x1269, x1270, x1271, x1272, x1273, x1274, x1275, x1276, x1277, x1278, x1279, x1280, x1281, x1282, x1283, x1284, x1285, x1286, x1287, x1288, x1289, x1290, x1291, x1292, x1293, x1294, x1295, x1296, x1297, x1298, x1299, x1300, x1301, x1302, x1303, x1304, x1305, x1306, x1307, x1308, x1309, x1310, x1311, x1312, x1313, x1314, x1315, x1316, x1317, x1318, x1319, x1320, x1321, x1322, x1323, x1324, x1325, x1326, x1327, x1328, x1329, x1330, x1331, x1332, x1333, x1334, x1335, x1336, x1337, x1338, x1339, x1340, x1341, x1342, x1343, x1344, x1345, x1346, x1347, x1348, x1349, x1350, x1351, x1352, x1353, x1354, x1355, x1356, x1357, x1358, x1359, x1360, x1361, x1362, x1363, x1364, x1365, x1366, x1367, x1368, x1369, x1370, x1371, x1372, x1373, x1374, x1375, x1376, x1377, x1378, x1379, x1380, x1381, x1382, x1383, x1384, x1385, x1386, x1387, x1388, x1389, x1390, x1391, x1392, x1393, x1394, x1395, x1396, x1397, x1398, x1399, x1400, x1401, x1402, x1403, x1404, x1405, x1406, x1407, x1408, x1409, x1410, x1411, x1412, x1413, x1414, x1415, x1416, x1417, x1418, x1419, x1420, x1421, x1422, x1423, x1424, x1425, x1426, x1427, x1428, x1429, x1430, x1431, x1432, x1433, x1434, x1435, x1436, x1437, x1438, x1439, x1440, x1441, x1442, x1443, x1444, x1445, x1446, x1447, x1448, x1449, x1450, x1451, x1452, x1453, x1454, x1455, x1456, x1457, x1458, x1459, x1460, x1461, x1462, x1463, x1464, x1465, x1466, x1467, x1468, x1469, x1470, x1471, x1472, x1473, x1474, x1475, x1476, x1477, x1478, x1479, x1480, x1481, x1482, x1483, x1484, x1485, x1486, x1487, x1488, x1489, x1490, x1491, x1492, x1493, x1494, x1495, x1496, x1497, x1498, x1499, x1500, x1501, x1502, x1503, x1504, x1505, x1506, x1507, x1508, x1509, x1510, x1511, x1512, x1513, x1514, x1515, x1516, x1517, x1518, x1519, x1520, x1521, x1522, x1523, x1524, x1525, x1526, x1527, x1528, x1529, x1530, x1531, x1532, x1533, x1534, x1535, x1536, x1537, x1538, x1539, x1540, x1541, x1542, x1543, x1544, x1545, x1546, x1547, x1548, x1549, x1550, x1551, x1552, x1553, x1554, x1555, x1556, x1557, x1558, x1559, x1560, x1561, x1562, x1563, x1564, x1565, x1566, x1567, x1568, x1569, x1570, x1571, x1572, x1573, x1574, x1575, x1576, x1577, x1578, x1579, x1580, x1581, x1582, x1583, x1584, x1585, x1586, x1587, x1588, x1589, x1590, x1591, x1592, x1593, x1594, x1595, x1596, x1597, x1598, x1599, x1600, x1601, x1602, x1603, x1604, x1605, x1606, x1607, x1608, x1609, x1610, x1611, x1612, x1613, x1614, x1615, x1616, x1617, x1618, x1619, x1620, x1621, x1622, x1623, x1624, x1625, x1626, x1627, x1628, x1629, x1630, x1631, x1632, x1633, x1634, x1635, x1636, x1637, x1638, x1639, x1640, x1641, x1642, x1643, x1644, x1645, x1646, x1647, x1648, x1649, x1650, x1651, x1652, x1653, x1654, x1655, x1656, x1657, x1658, x1659, x1660, x1661, x1662, x1663, x1664, x1665, x1666, x1667, x1668, x1669, x1670, x1671, x1672, x1673, x1674, x1675, x1676, x1677, x1678, x1679, x1680, x1681, x1682, x1683, x1684, x1685, x1686, x1687, x1688, x1689, x1690, x1691, x1692, x1693, x1694, x1695, x1696, x1697, x1698, x1699, x1700, x1701, x1702, x1703, x1704, x1705, x1706, x1707, x1708, x1709, x1710, x1711, x1712, x1713, x1714, x1715, x1716, x1717, x1718, x1719, x1720, x1721, x1722, x1723, x1724, x1725, x1726, x1727, x1728, x1729, x1730, x1731, x1732, x1733, x1734, x1735, x1736, x1737, x1738, x1739, x1740, x1741, x1742, x1743, x1744, x1745, x1746, x1747, x1748, x1749, x1750, x1751, x1752, x1753, x1754, x1755, x1756, x1757, x1758, x1759, x1760, x1761, x1762, x1763, x1764, x1765, x1766, x1767, x1768, x1769, x1770, x1771, x1772, x1773, x1774, x1775, x1776, x1777, x1778, x1779, x1780, x1781, x1782, x1783, x1784, x1785, x1786, x1787, x1788, x1789, x1790, x1791, x1792, x1793, x1794, x1795, x1796, x1797, x1798, x1799, x1800, x1801, x1802, x1803, x1804, x1805, x1806, x1807, x1808, x1809, x1810, x1811, x1812, x1813, x1814, x1815, x1816, x1817, x1818, x1819, x1820, x1821, x1822, x1823, x1824, x1825, x1826, x1827, x1828, x1829, x1830, x1831, x1832, x1833, x1834, x1835, x1836, x1837, x1838, x1839, x1840, x1841, x1842, x1843, x1844, x1845, x1846, x1847, x1848, x1849, x1850, x1851, x1852, x1853, x1854, x1855, x1856, x1857, x1858, x1859, x1860, x1861, x1862, x1863, x1864, x1865, x1866, x1867, x1868, x1869, x1870, x1871, x1872, x1873, x1874, x1875, x1876, x1877, x1878, x1879, x1880, x1881, x1882, x1883, x1884, x1885, x1886, x1887, x1888, x1889, x1890, x1891, x1892, x1893, x1894, x1895, x1896, x1897, x1898, x1899, x1900, x1901, x1902, x1903, x1904, x1905, x1906, x1907, x1908, x1909, x1910, x1911, x1912, x1913, x1914, x1915, x1916, x1917, x1918, x1919, x1920, x1921, x1922, x1923, x1924, x1925, x1926, x1927, x1928, x1929, x1930, x1931, x1932, x1933, x1934, x1935, x1936, x1937, x1938, x1939, x1940, x1941, x1942, x1943, x1944, x1945, x1946, x1947, x1948, x1949, x1950, x1951, x1952, x1953, x1954, x1955, x1956, x1957, x1958, x1959, x1960, x1961, x1962, x1963, x1964, x1965, x1966, x1967, x1968, x1969, x1970, x1971, x1972, x1973, x1974, x1975, x1976, x1977, x1978, x1979, x1980, x1981, x1982, x1983, x1984, x1985, x1986, x1987, x1988, x1989, x1990, x1991, x1992, x1993, x1994, x1995, x1996, x1997, x1998, x1999, x2000, x2001, x2002, x2003, x2004, x2005, x2006, x2007, x2008, x2009, x2010, x2011, x2012, x2013, x2014, x2015, x2016, x2017, x2018, x2019, x2020, x2021, x2022, x2023, x2024, y0);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255, x256, x257, x258, x259, x260, x261, x262, x263, x264, x265, x266, x267, x268, x269, x270, x271, x272, x273, x274, x275, x276, x277, x278, x279, x280, x281, x282, x283, x284, x285, x286, x287, x288, x289, x290, x291, x292, x293, x294, x295, x296, x297, x298, x299, x300, x301, x302, x303, x304, x305, x306, x307, x308, x309, x310, x311, x312, x313, x314, x315, x316, x317, x318, x319, x320, x321, x322, x323, x324, x325, x326, x327, x328, x329, x330, x331, x332, x333, x334, x335, x336, x337, x338, x339, x340, x341, x342, x343, x344, x345, x346, x347, x348, x349, x350, x351, x352, x353, x354, x355, x356, x357, x358, x359, x360, x361, x362, x363, x364, x365, x366, x367, x368, x369, x370, x371, x372, x373, x374, x375, x376, x377, x378, x379, x380, x381, x382, x383, x384, x385, x386, x387, x388, x389, x390, x391, x392, x393, x394, x395, x396, x397, x398, x399, x400, x401, x402, x403, x404, x405, x406, x407, x408, x409, x410, x411, x412, x413, x414, x415, x416, x417, x418, x419, x420, x421, x422, x423, x424, x425, x426, x427, x428, x429, x430, x431, x432, x433, x434, x435, x436, x437, x438, x439, x440, x441, x442, x443, x444, x445, x446, x447, x448, x449, x450, x451, x452, x453, x454, x455, x456, x457, x458, x459, x460, x461, x462, x463, x464, x465, x466, x467, x468, x469, x470, x471, x472, x473, x474, x475, x476, x477, x478, x479, x480, x481, x482, x483, x484, x485, x486, x487, x488, x489, x490, x491, x492, x493, x494, x495, x496, x497, x498, x499, x500, x501, x502, x503, x504, x505, x506, x507, x508, x509, x510, x511, x512, x513, x514, x515, x516, x517, x518, x519, x520, x521, x522, x523, x524, x525, x526, x527, x528, x529, x530, x531, x532, x533, x534, x535, x536, x537, x538, x539, x540, x541, x542, x543, x544, x545, x546, x547, x548, x549, x550, x551, x552, x553, x554, x555, x556, x557, x558, x559, x560, x561, x562, x563, x564, x565, x566, x567, x568, x569, x570, x571, x572, x573, x574, x575, x576, x577, x578, x579, x580, x581, x582, x583, x584, x585, x586, x587, x588, x589, x590, x591, x592, x593, x594, x595, x596, x597, x598, x599, x600, x601, x602, x603, x604, x605, x606, x607, x608, x609, x610, x611, x612, x613, x614, x615, x616, x617, x618, x619, x620, x621, x622, x623, x624, x625, x626, x627, x628, x629, x630, x631, x632, x633, x634, x635, x636, x637, x638, x639, x640, x641, x642, x643, x644, x645, x646, x647, x648, x649, x650, x651, x652, x653, x654, x655, x656, x657, x658, x659, x660, x661, x662, x663, x664, x665, x666, x667, x668, x669, x670, x671, x672, x673, x674, x675, x676, x677, x678, x679, x680, x681, x682, x683, x684, x685, x686, x687, x688, x689, x690, x691, x692, x693, x694, x695, x696, x697, x698, x699, x700, x701, x702, x703, x704, x705, x706, x707, x708, x709, x710, x711, x712, x713, x714, x715, x716, x717, x718, x719, x720, x721, x722, x723, x724, x725, x726, x727, x728, x729, x730, x731, x732, x733, x734, x735, x736, x737, x738, x739, x740, x741, x742, x743, x744, x745, x746, x747, x748, x749, x750, x751, x752, x753, x754, x755, x756, x757, x758, x759, x760, x761, x762, x763, x764, x765, x766, x767, x768, x769, x770, x771, x772, x773, x774, x775, x776, x777, x778, x779, x780, x781, x782, x783, x784, x785, x786, x787, x788, x789, x790, x791, x792, x793, x794, x795, x796, x797, x798, x799, x800, x801, x802, x803, x804, x805, x806, x807, x808, x809, x810, x811, x812, x813, x814, x815, x816, x817, x818, x819, x820, x821, x822, x823, x824, x825, x826, x827, x828, x829, x830, x831, x832, x833, x834, x835, x836, x837, x838, x839, x840, x841, x842, x843, x844, x845, x846, x847, x848, x849, x850, x851, x852, x853, x854, x855, x856, x857, x858, x859, x860, x861, x862, x863, x864, x865, x866, x867, x868, x869, x870, x871, x872, x873, x874, x875, x876, x877, x878, x879, x880, x881, x882, x883, x884, x885, x886, x887, x888, x889, x890, x891, x892, x893, x894, x895, x896, x897, x898, x899, x900, x901, x902, x903, x904, x905, x906, x907, x908, x909, x910, x911, x912, x913, x914, x915, x916, x917, x918, x919, x920, x921, x922, x923, x924, x925, x926, x927, x928, x929, x930, x931, x932, x933, x934, x935, x936, x937, x938, x939, x940, x941, x942, x943, x944, x945, x946, x947, x948, x949, x950, x951, x952, x953, x954, x955, x956, x957, x958, x959, x960, x961, x962, x963, x964, x965, x966, x967, x968, x969, x970, x971, x972, x973, x974, x975, x976, x977, x978, x979, x980, x981, x982, x983, x984, x985, x986, x987, x988, x989, x990, x991, x992, x993, x994, x995, x996, x997, x998, x999, x1000, x1001, x1002, x1003, x1004, x1005, x1006, x1007, x1008, x1009, x1010, x1011, x1012, x1013, x1014, x1015, x1016, x1017, x1018, x1019, x1020, x1021, x1022, x1023, x1024, x1025, x1026, x1027, x1028, x1029, x1030, x1031, x1032, x1033, x1034, x1035, x1036, x1037, x1038, x1039, x1040, x1041, x1042, x1043, x1044, x1045, x1046, x1047, x1048, x1049, x1050, x1051, x1052, x1053, x1054, x1055, x1056, x1057, x1058, x1059, x1060, x1061, x1062, x1063, x1064, x1065, x1066, x1067, x1068, x1069, x1070, x1071, x1072, x1073, x1074, x1075, x1076, x1077, x1078, x1079, x1080, x1081, x1082, x1083, x1084, x1085, x1086, x1087, x1088, x1089, x1090, x1091, x1092, x1093, x1094, x1095, x1096, x1097, x1098, x1099, x1100, x1101, x1102, x1103, x1104, x1105, x1106, x1107, x1108, x1109, x1110, x1111, x1112, x1113, x1114, x1115, x1116, x1117, x1118, x1119, x1120, x1121, x1122, x1123, x1124, x1125, x1126, x1127, x1128, x1129, x1130, x1131, x1132, x1133, x1134, x1135, x1136, x1137, x1138, x1139, x1140, x1141, x1142, x1143, x1144, x1145, x1146, x1147, x1148, x1149, x1150, x1151, x1152, x1153, x1154, x1155, x1156, x1157, x1158, x1159, x1160, x1161, x1162, x1163, x1164, x1165, x1166, x1167, x1168, x1169, x1170, x1171, x1172, x1173, x1174, x1175, x1176, x1177, x1178, x1179, x1180, x1181, x1182, x1183, x1184, x1185, x1186, x1187, x1188, x1189, x1190, x1191, x1192, x1193, x1194, x1195, x1196, x1197, x1198, x1199, x1200, x1201, x1202, x1203, x1204, x1205, x1206, x1207, x1208, x1209, x1210, x1211, x1212, x1213, x1214, x1215, x1216, x1217, x1218, x1219, x1220, x1221, x1222, x1223, x1224, x1225, x1226, x1227, x1228, x1229, x1230, x1231, x1232, x1233, x1234, x1235, x1236, x1237, x1238, x1239, x1240, x1241, x1242, x1243, x1244, x1245, x1246, x1247, x1248, x1249, x1250, x1251, x1252, x1253, x1254, x1255, x1256, x1257, x1258, x1259, x1260, x1261, x1262, x1263, x1264, x1265, x1266, x1267, x1268, x1269, x1270, x1271, x1272, x1273, x1274, x1275, x1276, x1277, x1278, x1279, x1280, x1281, x1282, x1283, x1284, x1285, x1286, x1287, x1288, x1289, x1290, x1291, x1292, x1293, x1294, x1295, x1296, x1297, x1298, x1299, x1300, x1301, x1302, x1303, x1304, x1305, x1306, x1307, x1308, x1309, x1310, x1311, x1312, x1313, x1314, x1315, x1316, x1317, x1318, x1319, x1320, x1321, x1322, x1323, x1324, x1325, x1326, x1327, x1328, x1329, x1330, x1331, x1332, x1333, x1334, x1335, x1336, x1337, x1338, x1339, x1340, x1341, x1342, x1343, x1344, x1345, x1346, x1347, x1348, x1349, x1350, x1351, x1352, x1353, x1354, x1355, x1356, x1357, x1358, x1359, x1360, x1361, x1362, x1363, x1364, x1365, x1366, x1367, x1368, x1369, x1370, x1371, x1372, x1373, x1374, x1375, x1376, x1377, x1378, x1379, x1380, x1381, x1382, x1383, x1384, x1385, x1386, x1387, x1388, x1389, x1390, x1391, x1392, x1393, x1394, x1395, x1396, x1397, x1398, x1399, x1400, x1401, x1402, x1403, x1404, x1405, x1406, x1407, x1408, x1409, x1410, x1411, x1412, x1413, x1414, x1415, x1416, x1417, x1418, x1419, x1420, x1421, x1422, x1423, x1424, x1425, x1426, x1427, x1428, x1429, x1430, x1431, x1432, x1433, x1434, x1435, x1436, x1437, x1438, x1439, x1440, x1441, x1442, x1443, x1444, x1445, x1446, x1447, x1448, x1449, x1450, x1451, x1452, x1453, x1454, x1455, x1456, x1457, x1458, x1459, x1460, x1461, x1462, x1463, x1464, x1465, x1466, x1467, x1468, x1469, x1470, x1471, x1472, x1473, x1474, x1475, x1476, x1477, x1478, x1479, x1480, x1481, x1482, x1483, x1484, x1485, x1486, x1487, x1488, x1489, x1490, x1491, x1492, x1493, x1494, x1495, x1496, x1497, x1498, x1499, x1500, x1501, x1502, x1503, x1504, x1505, x1506, x1507, x1508, x1509, x1510, x1511, x1512, x1513, x1514, x1515, x1516, x1517, x1518, x1519, x1520, x1521, x1522, x1523, x1524, x1525, x1526, x1527, x1528, x1529, x1530, x1531, x1532, x1533, x1534, x1535, x1536, x1537, x1538, x1539, x1540, x1541, x1542, x1543, x1544, x1545, x1546, x1547, x1548, x1549, x1550, x1551, x1552, x1553, x1554, x1555, x1556, x1557, x1558, x1559, x1560, x1561, x1562, x1563, x1564, x1565, x1566, x1567, x1568, x1569, x1570, x1571, x1572, x1573, x1574, x1575, x1576, x1577, x1578, x1579, x1580, x1581, x1582, x1583, x1584, x1585, x1586, x1587, x1588, x1589, x1590, x1591, x1592, x1593, x1594, x1595, x1596, x1597, x1598, x1599, x1600, x1601, x1602, x1603, x1604, x1605, x1606, x1607, x1608, x1609, x1610, x1611, x1612, x1613, x1614, x1615, x1616, x1617, x1618, x1619, x1620, x1621, x1622, x1623, x1624, x1625, x1626, x1627, x1628, x1629, x1630, x1631, x1632, x1633, x1634, x1635, x1636, x1637, x1638, x1639, x1640, x1641, x1642, x1643, x1644, x1645, x1646, x1647, x1648, x1649, x1650, x1651, x1652, x1653, x1654, x1655, x1656, x1657, x1658, x1659, x1660, x1661, x1662, x1663, x1664, x1665, x1666, x1667, x1668, x1669, x1670, x1671, x1672, x1673, x1674, x1675, x1676, x1677, x1678, x1679, x1680, x1681, x1682, x1683, x1684, x1685, x1686, x1687, x1688, x1689, x1690, x1691, x1692, x1693, x1694, x1695, x1696, x1697, x1698, x1699, x1700, x1701, x1702, x1703, x1704, x1705, x1706, x1707, x1708, x1709, x1710, x1711, x1712, x1713, x1714, x1715, x1716, x1717, x1718, x1719, x1720, x1721, x1722, x1723, x1724, x1725, x1726, x1727, x1728, x1729, x1730, x1731, x1732, x1733, x1734, x1735, x1736, x1737, x1738, x1739, x1740, x1741, x1742, x1743, x1744, x1745, x1746, x1747, x1748, x1749, x1750, x1751, x1752, x1753, x1754, x1755, x1756, x1757, x1758, x1759, x1760, x1761, x1762, x1763, x1764, x1765, x1766, x1767, x1768, x1769, x1770, x1771, x1772, x1773, x1774, x1775, x1776, x1777, x1778, x1779, x1780, x1781, x1782, x1783, x1784, x1785, x1786, x1787, x1788, x1789, x1790, x1791, x1792, x1793, x1794, x1795, x1796, x1797, x1798, x1799, x1800, x1801, x1802, x1803, x1804, x1805, x1806, x1807, x1808, x1809, x1810, x1811, x1812, x1813, x1814, x1815, x1816, x1817, x1818, x1819, x1820, x1821, x1822, x1823, x1824, x1825, x1826, x1827, x1828, x1829, x1830, x1831, x1832, x1833, x1834, x1835, x1836, x1837, x1838, x1839, x1840, x1841, x1842, x1843, x1844, x1845, x1846, x1847, x1848, x1849, x1850, x1851, x1852, x1853, x1854, x1855, x1856, x1857, x1858, x1859, x1860, x1861, x1862, x1863, x1864, x1865, x1866, x1867, x1868, x1869, x1870, x1871, x1872, x1873, x1874, x1875, x1876, x1877, x1878, x1879, x1880, x1881, x1882, x1883, x1884, x1885, x1886, x1887, x1888, x1889, x1890, x1891, x1892, x1893, x1894, x1895, x1896, x1897, x1898, x1899, x1900, x1901, x1902, x1903, x1904, x1905, x1906, x1907, x1908, x1909, x1910, x1911, x1912, x1913, x1914, x1915, x1916, x1917, x1918, x1919, x1920, x1921, x1922, x1923, x1924, x1925, x1926, x1927, x1928, x1929, x1930, x1931, x1932, x1933, x1934, x1935, x1936, x1937, x1938, x1939, x1940, x1941, x1942, x1943, x1944, x1945, x1946, x1947, x1948, x1949, x1950, x1951, x1952, x1953, x1954, x1955, x1956, x1957, x1958, x1959, x1960, x1961, x1962, x1963, x1964, x1965, x1966, x1967, x1968, x1969, x1970, x1971, x1972, x1973, x1974, x1975, x1976, x1977, x1978, x1979, x1980, x1981, x1982, x1983, x1984, x1985, x1986, x1987, x1988, x1989, x1990, x1991, x1992, x1993, x1994, x1995, x1996, x1997, x1998, x1999, x2000, x2001, x2002, x2003, x2004, x2005, x2006, x2007, x2008, x2009, x2010, x2011, x2012, x2013, x2014, x2015, x2016, x2017, x2018, x2019, x2020, x2021, x2022, x2023, x2024;
  output y0;
  wire n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368;
  LUT3 #(.INIT(8'hE8)) lut_n2027 (.I0(x0), .I1(x1), .I2(x2), .O(n2027));
  LUT3 #(.INIT(8'hE8)) lut_n2028 (.I0(x6), .I1(x7), .I2(x8), .O(n2028));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2029 (.I0(x3), .I1(x4), .I2(x5), .I3(n2027), .I4(n2028), .O(n2029));
  LUT3 #(.INIT(8'hE8)) lut_n2030 (.I0(x12), .I1(x13), .I2(x14), .O(n2030));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2031 (.I0(x3), .I1(x4), .I2(x5), .I3(n2027), .I4(n2028), .O(n2031));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2032 (.I0(x9), .I1(x10), .I2(x11), .I3(n2030), .I4(n2031), .O(n2032));
  LUT3 #(.INIT(8'hE8)) lut_n2033 (.I0(x18), .I1(x19), .I2(x20), .O(n2033));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2034 (.I0(x9), .I1(x10), .I2(x11), .I3(n2030), .I4(n2031), .O(n2034));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2035 (.I0(x15), .I1(x16), .I2(x17), .I3(n2033), .I4(n2034), .O(n2035));
  LUT3 #(.INIT(8'hE8)) lut_n2036 (.I0(n2029), .I1(n2032), .I2(n2035), .O(n2036));
  LUT3 #(.INIT(8'hE8)) lut_n2037 (.I0(x24), .I1(x25), .I2(x26), .O(n2037));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2038 (.I0(x15), .I1(x16), .I2(x17), .I3(n2033), .I4(n2034), .O(n2038));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2039 (.I0(x21), .I1(x22), .I2(x23), .I3(n2037), .I4(n2038), .O(n2039));
  LUT3 #(.INIT(8'hE8)) lut_n2040 (.I0(x27), .I1(x28), .I2(x29), .O(n2040));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2041 (.I0(x21), .I1(x22), .I2(x23), .I3(n2037), .I4(n2038), .O(n2041));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2042 (.I0(x30), .I1(x31), .I2(x32), .I3(n2040), .I4(n2041), .O(n2042));
  LUT3 #(.INIT(8'h96)) lut_n2043 (.I0(n2029), .I1(n2032), .I2(n2035), .O(n2043));
  LUT3 #(.INIT(8'hE8)) lut_n2044 (.I0(n2039), .I1(n2042), .I2(n2043), .O(n2044));
  LUT3 #(.INIT(8'hE8)) lut_n2045 (.I0(x36), .I1(x37), .I2(x38), .O(n2045));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2046 (.I0(x30), .I1(x31), .I2(x32), .I3(n2040), .I4(n2041), .O(n2046));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2047 (.I0(x33), .I1(x34), .I2(x35), .I3(n2045), .I4(n2046), .O(n2047));
  LUT3 #(.INIT(8'hE8)) lut_n2048 (.I0(x42), .I1(x43), .I2(x44), .O(n2048));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2049 (.I0(x33), .I1(x34), .I2(x35), .I3(n2045), .I4(n2046), .O(n2049));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2050 (.I0(x39), .I1(x40), .I2(x41), .I3(n2048), .I4(n2049), .O(n2050));
  LUT3 #(.INIT(8'h96)) lut_n2051 (.I0(n2039), .I1(n2042), .I2(n2043), .O(n2051));
  LUT3 #(.INIT(8'hE8)) lut_n2052 (.I0(n2047), .I1(n2050), .I2(n2051), .O(n2052));
  LUT3 #(.INIT(8'hE8)) lut_n2053 (.I0(n2036), .I1(n2044), .I2(n2052), .O(n2053));
  LUT3 #(.INIT(8'hE8)) lut_n2054 (.I0(x48), .I1(x49), .I2(x50), .O(n2054));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2055 (.I0(x39), .I1(x40), .I2(x41), .I3(n2048), .I4(n2049), .O(n2055));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2056 (.I0(x45), .I1(x46), .I2(x47), .I3(n2054), .I4(n2055), .O(n2056));
  LUT3 #(.INIT(8'hE8)) lut_n2057 (.I0(x54), .I1(x55), .I2(x56), .O(n2057));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2058 (.I0(x45), .I1(x46), .I2(x47), .I3(n2054), .I4(n2055), .O(n2058));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2059 (.I0(x51), .I1(x52), .I2(x53), .I3(n2057), .I4(n2058), .O(n2059));
  LUT3 #(.INIT(8'h96)) lut_n2060 (.I0(n2047), .I1(n2050), .I2(n2051), .O(n2060));
  LUT3 #(.INIT(8'hE8)) lut_n2061 (.I0(n2056), .I1(n2059), .I2(n2060), .O(n2061));
  LUT3 #(.INIT(8'hE8)) lut_n2062 (.I0(x60), .I1(x61), .I2(x62), .O(n2062));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2063 (.I0(x51), .I1(x52), .I2(x53), .I3(n2057), .I4(n2058), .O(n2063));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2064 (.I0(x57), .I1(x58), .I2(x59), .I3(n2062), .I4(n2063), .O(n2064));
  LUT3 #(.INIT(8'hE8)) lut_n2065 (.I0(x66), .I1(x67), .I2(x68), .O(n2065));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2066 (.I0(x57), .I1(x58), .I2(x59), .I3(n2062), .I4(n2063), .O(n2066));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2067 (.I0(x63), .I1(x64), .I2(x65), .I3(n2065), .I4(n2066), .O(n2067));
  LUT3 #(.INIT(8'h96)) lut_n2068 (.I0(n2056), .I1(n2059), .I2(n2060), .O(n2068));
  LUT3 #(.INIT(8'hE8)) lut_n2069 (.I0(n2064), .I1(n2067), .I2(n2068), .O(n2069));
  LUT3 #(.INIT(8'h96)) lut_n2070 (.I0(n2036), .I1(n2044), .I2(n2052), .O(n2070));
  LUT3 #(.INIT(8'hE8)) lut_n2071 (.I0(n2061), .I1(n2069), .I2(n2070), .O(n2071));
  LUT3 #(.INIT(8'hE8)) lut_n2072 (.I0(x72), .I1(x73), .I2(x74), .O(n2072));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2073 (.I0(x63), .I1(x64), .I2(x65), .I3(n2065), .I4(n2066), .O(n2073));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2074 (.I0(x69), .I1(x70), .I2(x71), .I3(n2072), .I4(n2073), .O(n2074));
  LUT3 #(.INIT(8'hE8)) lut_n2075 (.I0(x78), .I1(x79), .I2(x80), .O(n2075));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2076 (.I0(x69), .I1(x70), .I2(x71), .I3(n2072), .I4(n2073), .O(n2076));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2077 (.I0(x75), .I1(x76), .I2(x77), .I3(n2075), .I4(n2076), .O(n2077));
  LUT3 #(.INIT(8'h96)) lut_n2078 (.I0(n2064), .I1(n2067), .I2(n2068), .O(n2078));
  LUT3 #(.INIT(8'hE8)) lut_n2079 (.I0(n2074), .I1(n2077), .I2(n2078), .O(n2079));
  LUT3 #(.INIT(8'hE8)) lut_n2080 (.I0(x84), .I1(x85), .I2(x86), .O(n2080));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2081 (.I0(x75), .I1(x76), .I2(x77), .I3(n2075), .I4(n2076), .O(n2081));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2082 (.I0(x81), .I1(x82), .I2(x83), .I3(n2080), .I4(n2081), .O(n2082));
  LUT3 #(.INIT(8'hE8)) lut_n2083 (.I0(x90), .I1(x91), .I2(x92), .O(n2083));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2084 (.I0(x81), .I1(x82), .I2(x83), .I3(n2080), .I4(n2081), .O(n2084));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2085 (.I0(x87), .I1(x88), .I2(x89), .I3(n2083), .I4(n2084), .O(n2085));
  LUT3 #(.INIT(8'h96)) lut_n2086 (.I0(n2074), .I1(n2077), .I2(n2078), .O(n2086));
  LUT3 #(.INIT(8'hE8)) lut_n2087 (.I0(n2082), .I1(n2085), .I2(n2086), .O(n2087));
  LUT3 #(.INIT(8'h96)) lut_n2088 (.I0(n2061), .I1(n2069), .I2(n2070), .O(n2088));
  LUT3 #(.INIT(8'hE8)) lut_n2089 (.I0(n2079), .I1(n2087), .I2(n2088), .O(n2089));
  LUT3 #(.INIT(8'hE8)) lut_n2090 (.I0(n2053), .I1(n2071), .I2(n2089), .O(n2090));
  LUT3 #(.INIT(8'hE8)) lut_n2091 (.I0(x96), .I1(x97), .I2(x98), .O(n2091));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2092 (.I0(x87), .I1(x88), .I2(x89), .I3(n2083), .I4(n2084), .O(n2092));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2093 (.I0(x93), .I1(x94), .I2(x95), .I3(n2091), .I4(n2092), .O(n2093));
  LUT3 #(.INIT(8'hE8)) lut_n2094 (.I0(x102), .I1(x103), .I2(x104), .O(n2094));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2095 (.I0(x93), .I1(x94), .I2(x95), .I3(n2091), .I4(n2092), .O(n2095));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2096 (.I0(x99), .I1(x100), .I2(x101), .I3(n2094), .I4(n2095), .O(n2096));
  LUT3 #(.INIT(8'h96)) lut_n2097 (.I0(n2082), .I1(n2085), .I2(n2086), .O(n2097));
  LUT3 #(.INIT(8'hE8)) lut_n2098 (.I0(n2093), .I1(n2096), .I2(n2097), .O(n2098));
  LUT3 #(.INIT(8'hE8)) lut_n2099 (.I0(x108), .I1(x109), .I2(x110), .O(n2099));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2100 (.I0(x99), .I1(x100), .I2(x101), .I3(n2094), .I4(n2095), .O(n2100));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2101 (.I0(x105), .I1(x106), .I2(x107), .I3(n2099), .I4(n2100), .O(n2101));
  LUT3 #(.INIT(8'hE8)) lut_n2102 (.I0(x114), .I1(x115), .I2(x116), .O(n2102));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2103 (.I0(x105), .I1(x106), .I2(x107), .I3(n2099), .I4(n2100), .O(n2103));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2104 (.I0(x111), .I1(x112), .I2(x113), .I3(n2102), .I4(n2103), .O(n2104));
  LUT3 #(.INIT(8'h96)) lut_n2105 (.I0(n2093), .I1(n2096), .I2(n2097), .O(n2105));
  LUT3 #(.INIT(8'hE8)) lut_n2106 (.I0(n2101), .I1(n2104), .I2(n2105), .O(n2106));
  LUT3 #(.INIT(8'h96)) lut_n2107 (.I0(n2079), .I1(n2087), .I2(n2088), .O(n2107));
  LUT3 #(.INIT(8'hE8)) lut_n2108 (.I0(n2098), .I1(n2106), .I2(n2107), .O(n2108));
  LUT3 #(.INIT(8'hE8)) lut_n2109 (.I0(x120), .I1(x121), .I2(x122), .O(n2109));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2110 (.I0(x111), .I1(x112), .I2(x113), .I3(n2102), .I4(n2103), .O(n2110));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2111 (.I0(x117), .I1(x118), .I2(x119), .I3(n2109), .I4(n2110), .O(n2111));
  LUT3 #(.INIT(8'hE8)) lut_n2112 (.I0(x126), .I1(x127), .I2(x128), .O(n2112));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2113 (.I0(x117), .I1(x118), .I2(x119), .I3(n2109), .I4(n2110), .O(n2113));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2114 (.I0(x123), .I1(x124), .I2(x125), .I3(n2112), .I4(n2113), .O(n2114));
  LUT3 #(.INIT(8'h96)) lut_n2115 (.I0(n2101), .I1(n2104), .I2(n2105), .O(n2115));
  LUT3 #(.INIT(8'hE8)) lut_n2116 (.I0(n2111), .I1(n2114), .I2(n2115), .O(n2116));
  LUT3 #(.INIT(8'hE8)) lut_n2117 (.I0(x132), .I1(x133), .I2(x134), .O(n2117));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2118 (.I0(x123), .I1(x124), .I2(x125), .I3(n2112), .I4(n2113), .O(n2118));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2119 (.I0(x129), .I1(x130), .I2(x131), .I3(n2117), .I4(n2118), .O(n2119));
  LUT3 #(.INIT(8'hE8)) lut_n2120 (.I0(x138), .I1(x139), .I2(x140), .O(n2120));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2121 (.I0(x129), .I1(x130), .I2(x131), .I3(n2117), .I4(n2118), .O(n2121));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2122 (.I0(x135), .I1(x136), .I2(x137), .I3(n2120), .I4(n2121), .O(n2122));
  LUT3 #(.INIT(8'h96)) lut_n2123 (.I0(n2111), .I1(n2114), .I2(n2115), .O(n2123));
  LUT3 #(.INIT(8'hE8)) lut_n2124 (.I0(n2119), .I1(n2122), .I2(n2123), .O(n2124));
  LUT3 #(.INIT(8'h96)) lut_n2125 (.I0(n2098), .I1(n2106), .I2(n2107), .O(n2125));
  LUT3 #(.INIT(8'hE8)) lut_n2126 (.I0(n2116), .I1(n2124), .I2(n2125), .O(n2126));
  LUT3 #(.INIT(8'h96)) lut_n2127 (.I0(n2053), .I1(n2071), .I2(n2089), .O(n2127));
  LUT3 #(.INIT(8'hE8)) lut_n2128 (.I0(n2108), .I1(n2126), .I2(n2127), .O(n2128));
  LUT3 #(.INIT(8'hE8)) lut_n2129 (.I0(x144), .I1(x145), .I2(x146), .O(n2129));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2130 (.I0(x135), .I1(x136), .I2(x137), .I3(n2120), .I4(n2121), .O(n2130));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2131 (.I0(x141), .I1(x142), .I2(x143), .I3(n2129), .I4(n2130), .O(n2131));
  LUT3 #(.INIT(8'hE8)) lut_n2132 (.I0(x150), .I1(x151), .I2(x152), .O(n2132));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2133 (.I0(x141), .I1(x142), .I2(x143), .I3(n2129), .I4(n2130), .O(n2133));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2134 (.I0(x147), .I1(x148), .I2(x149), .I3(n2132), .I4(n2133), .O(n2134));
  LUT3 #(.INIT(8'h96)) lut_n2135 (.I0(n2119), .I1(n2122), .I2(n2123), .O(n2135));
  LUT3 #(.INIT(8'hE8)) lut_n2136 (.I0(n2131), .I1(n2134), .I2(n2135), .O(n2136));
  LUT3 #(.INIT(8'hE8)) lut_n2137 (.I0(x156), .I1(x157), .I2(x158), .O(n2137));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2138 (.I0(x147), .I1(x148), .I2(x149), .I3(n2132), .I4(n2133), .O(n2138));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2139 (.I0(x153), .I1(x154), .I2(x155), .I3(n2137), .I4(n2138), .O(n2139));
  LUT3 #(.INIT(8'hE8)) lut_n2140 (.I0(x162), .I1(x163), .I2(x164), .O(n2140));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2141 (.I0(x153), .I1(x154), .I2(x155), .I3(n2137), .I4(n2138), .O(n2141));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2142 (.I0(x159), .I1(x160), .I2(x161), .I3(n2140), .I4(n2141), .O(n2142));
  LUT3 #(.INIT(8'h96)) lut_n2143 (.I0(n2131), .I1(n2134), .I2(n2135), .O(n2143));
  LUT3 #(.INIT(8'hE8)) lut_n2144 (.I0(n2139), .I1(n2142), .I2(n2143), .O(n2144));
  LUT3 #(.INIT(8'h96)) lut_n2145 (.I0(n2116), .I1(n2124), .I2(n2125), .O(n2145));
  LUT3 #(.INIT(8'hE8)) lut_n2146 (.I0(n2136), .I1(n2144), .I2(n2145), .O(n2146));
  LUT3 #(.INIT(8'hE8)) lut_n2147 (.I0(x168), .I1(x169), .I2(x170), .O(n2147));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2148 (.I0(x159), .I1(x160), .I2(x161), .I3(n2140), .I4(n2141), .O(n2148));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2149 (.I0(x165), .I1(x166), .I2(x167), .I3(n2147), .I4(n2148), .O(n2149));
  LUT3 #(.INIT(8'hE8)) lut_n2150 (.I0(x174), .I1(x175), .I2(x176), .O(n2150));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2151 (.I0(x165), .I1(x166), .I2(x167), .I3(n2147), .I4(n2148), .O(n2151));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2152 (.I0(x171), .I1(x172), .I2(x173), .I3(n2150), .I4(n2151), .O(n2152));
  LUT3 #(.INIT(8'h96)) lut_n2153 (.I0(n2139), .I1(n2142), .I2(n2143), .O(n2153));
  LUT3 #(.INIT(8'hE8)) lut_n2154 (.I0(n2149), .I1(n2152), .I2(n2153), .O(n2154));
  LUT3 #(.INIT(8'hE8)) lut_n2155 (.I0(x180), .I1(x181), .I2(x182), .O(n2155));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2156 (.I0(x171), .I1(x172), .I2(x173), .I3(n2150), .I4(n2151), .O(n2156));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2157 (.I0(x177), .I1(x178), .I2(x179), .I3(n2155), .I4(n2156), .O(n2157));
  LUT3 #(.INIT(8'hE8)) lut_n2158 (.I0(x186), .I1(x187), .I2(x188), .O(n2158));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2159 (.I0(x177), .I1(x178), .I2(x179), .I3(n2155), .I4(n2156), .O(n2159));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2160 (.I0(x183), .I1(x184), .I2(x185), .I3(n2158), .I4(n2159), .O(n2160));
  LUT3 #(.INIT(8'h96)) lut_n2161 (.I0(n2149), .I1(n2152), .I2(n2153), .O(n2161));
  LUT3 #(.INIT(8'hE8)) lut_n2162 (.I0(n2157), .I1(n2160), .I2(n2161), .O(n2162));
  LUT3 #(.INIT(8'h96)) lut_n2163 (.I0(n2136), .I1(n2144), .I2(n2145), .O(n2163));
  LUT3 #(.INIT(8'hE8)) lut_n2164 (.I0(n2154), .I1(n2162), .I2(n2163), .O(n2164));
  LUT3 #(.INIT(8'h96)) lut_n2165 (.I0(n2108), .I1(n2126), .I2(n2127), .O(n2165));
  LUT3 #(.INIT(8'hE8)) lut_n2166 (.I0(n2146), .I1(n2164), .I2(n2165), .O(n2166));
  LUT3 #(.INIT(8'hE8)) lut_n2167 (.I0(n2090), .I1(n2128), .I2(n2166), .O(n2167));
  LUT3 #(.INIT(8'hE8)) lut_n2168 (.I0(x192), .I1(x193), .I2(x194), .O(n2168));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2169 (.I0(x183), .I1(x184), .I2(x185), .I3(n2158), .I4(n2159), .O(n2169));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2170 (.I0(x189), .I1(x190), .I2(x191), .I3(n2168), .I4(n2169), .O(n2170));
  LUT3 #(.INIT(8'hE8)) lut_n2171 (.I0(x198), .I1(x199), .I2(x200), .O(n2171));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2172 (.I0(x189), .I1(x190), .I2(x191), .I3(n2168), .I4(n2169), .O(n2172));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2173 (.I0(x195), .I1(x196), .I2(x197), .I3(n2171), .I4(n2172), .O(n2173));
  LUT3 #(.INIT(8'h96)) lut_n2174 (.I0(n2157), .I1(n2160), .I2(n2161), .O(n2174));
  LUT3 #(.INIT(8'hE8)) lut_n2175 (.I0(n2170), .I1(n2173), .I2(n2174), .O(n2175));
  LUT3 #(.INIT(8'hE8)) lut_n2176 (.I0(x204), .I1(x205), .I2(x206), .O(n2176));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2177 (.I0(x195), .I1(x196), .I2(x197), .I3(n2171), .I4(n2172), .O(n2177));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2178 (.I0(x201), .I1(x202), .I2(x203), .I3(n2176), .I4(n2177), .O(n2178));
  LUT3 #(.INIT(8'hE8)) lut_n2179 (.I0(x210), .I1(x211), .I2(x212), .O(n2179));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2180 (.I0(x201), .I1(x202), .I2(x203), .I3(n2176), .I4(n2177), .O(n2180));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2181 (.I0(x207), .I1(x208), .I2(x209), .I3(n2179), .I4(n2180), .O(n2181));
  LUT3 #(.INIT(8'h96)) lut_n2182 (.I0(n2170), .I1(n2173), .I2(n2174), .O(n2182));
  LUT3 #(.INIT(8'hE8)) lut_n2183 (.I0(n2178), .I1(n2181), .I2(n2182), .O(n2183));
  LUT3 #(.INIT(8'h96)) lut_n2184 (.I0(n2154), .I1(n2162), .I2(n2163), .O(n2184));
  LUT3 #(.INIT(8'hE8)) lut_n2185 (.I0(n2175), .I1(n2183), .I2(n2184), .O(n2185));
  LUT3 #(.INIT(8'hE8)) lut_n2186 (.I0(x216), .I1(x217), .I2(x218), .O(n2186));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2187 (.I0(x207), .I1(x208), .I2(x209), .I3(n2179), .I4(n2180), .O(n2187));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2188 (.I0(x213), .I1(x214), .I2(x215), .I3(n2186), .I4(n2187), .O(n2188));
  LUT3 #(.INIT(8'hE8)) lut_n2189 (.I0(x222), .I1(x223), .I2(x224), .O(n2189));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2190 (.I0(x213), .I1(x214), .I2(x215), .I3(n2186), .I4(n2187), .O(n2190));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2191 (.I0(x219), .I1(x220), .I2(x221), .I3(n2189), .I4(n2190), .O(n2191));
  LUT3 #(.INIT(8'h96)) lut_n2192 (.I0(n2178), .I1(n2181), .I2(n2182), .O(n2192));
  LUT3 #(.INIT(8'hE8)) lut_n2193 (.I0(n2188), .I1(n2191), .I2(n2192), .O(n2193));
  LUT3 #(.INIT(8'hE8)) lut_n2194 (.I0(x228), .I1(x229), .I2(x230), .O(n2194));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2195 (.I0(x219), .I1(x220), .I2(x221), .I3(n2189), .I4(n2190), .O(n2195));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2196 (.I0(x225), .I1(x226), .I2(x227), .I3(n2194), .I4(n2195), .O(n2196));
  LUT3 #(.INIT(8'hE8)) lut_n2197 (.I0(x234), .I1(x235), .I2(x236), .O(n2197));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2198 (.I0(x225), .I1(x226), .I2(x227), .I3(n2194), .I4(n2195), .O(n2198));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2199 (.I0(x231), .I1(x232), .I2(x233), .I3(n2197), .I4(n2198), .O(n2199));
  LUT3 #(.INIT(8'h96)) lut_n2200 (.I0(n2188), .I1(n2191), .I2(n2192), .O(n2200));
  LUT3 #(.INIT(8'hE8)) lut_n2201 (.I0(n2196), .I1(n2199), .I2(n2200), .O(n2201));
  LUT3 #(.INIT(8'h96)) lut_n2202 (.I0(n2175), .I1(n2183), .I2(n2184), .O(n2202));
  LUT3 #(.INIT(8'hE8)) lut_n2203 (.I0(n2193), .I1(n2201), .I2(n2202), .O(n2203));
  LUT3 #(.INIT(8'h96)) lut_n2204 (.I0(n2146), .I1(n2164), .I2(n2165), .O(n2204));
  LUT3 #(.INIT(8'hE8)) lut_n2205 (.I0(n2185), .I1(n2203), .I2(n2204), .O(n2205));
  LUT3 #(.INIT(8'hE8)) lut_n2206 (.I0(x240), .I1(x241), .I2(x242), .O(n2206));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2207 (.I0(x231), .I1(x232), .I2(x233), .I3(n2197), .I4(n2198), .O(n2207));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2208 (.I0(x237), .I1(x238), .I2(x239), .I3(n2206), .I4(n2207), .O(n2208));
  LUT3 #(.INIT(8'hE8)) lut_n2209 (.I0(x246), .I1(x247), .I2(x248), .O(n2209));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2210 (.I0(x237), .I1(x238), .I2(x239), .I3(n2206), .I4(n2207), .O(n2210));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2211 (.I0(x243), .I1(x244), .I2(x245), .I3(n2209), .I4(n2210), .O(n2211));
  LUT3 #(.INIT(8'h96)) lut_n2212 (.I0(n2196), .I1(n2199), .I2(n2200), .O(n2212));
  LUT3 #(.INIT(8'hE8)) lut_n2213 (.I0(n2208), .I1(n2211), .I2(n2212), .O(n2213));
  LUT3 #(.INIT(8'hE8)) lut_n2214 (.I0(x252), .I1(x253), .I2(x254), .O(n2214));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2215 (.I0(x243), .I1(x244), .I2(x245), .I3(n2209), .I4(n2210), .O(n2215));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2216 (.I0(x249), .I1(x250), .I2(x251), .I3(n2214), .I4(n2215), .O(n2216));
  LUT3 #(.INIT(8'hE8)) lut_n2217 (.I0(x258), .I1(x259), .I2(x260), .O(n2217));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2218 (.I0(x249), .I1(x250), .I2(x251), .I3(n2214), .I4(n2215), .O(n2218));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2219 (.I0(x255), .I1(x256), .I2(x257), .I3(n2217), .I4(n2218), .O(n2219));
  LUT3 #(.INIT(8'h96)) lut_n2220 (.I0(n2208), .I1(n2211), .I2(n2212), .O(n2220));
  LUT3 #(.INIT(8'hE8)) lut_n2221 (.I0(n2216), .I1(n2219), .I2(n2220), .O(n2221));
  LUT3 #(.INIT(8'h96)) lut_n2222 (.I0(n2193), .I1(n2201), .I2(n2202), .O(n2222));
  LUT3 #(.INIT(8'hE8)) lut_n2223 (.I0(n2213), .I1(n2221), .I2(n2222), .O(n2223));
  LUT3 #(.INIT(8'hE8)) lut_n2224 (.I0(x264), .I1(x265), .I2(x266), .O(n2224));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2225 (.I0(x255), .I1(x256), .I2(x257), .I3(n2217), .I4(n2218), .O(n2225));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2226 (.I0(x261), .I1(x262), .I2(x263), .I3(n2224), .I4(n2225), .O(n2226));
  LUT3 #(.INIT(8'hE8)) lut_n2227 (.I0(x270), .I1(x271), .I2(x272), .O(n2227));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2228 (.I0(x261), .I1(x262), .I2(x263), .I3(n2224), .I4(n2225), .O(n2228));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2229 (.I0(x267), .I1(x268), .I2(x269), .I3(n2227), .I4(n2228), .O(n2229));
  LUT3 #(.INIT(8'h96)) lut_n2230 (.I0(n2216), .I1(n2219), .I2(n2220), .O(n2230));
  LUT3 #(.INIT(8'hE8)) lut_n2231 (.I0(n2226), .I1(n2229), .I2(n2230), .O(n2231));
  LUT3 #(.INIT(8'hE8)) lut_n2232 (.I0(x276), .I1(x277), .I2(x278), .O(n2232));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2233 (.I0(x267), .I1(x268), .I2(x269), .I3(n2227), .I4(n2228), .O(n2233));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2234 (.I0(x273), .I1(x274), .I2(x275), .I3(n2232), .I4(n2233), .O(n2234));
  LUT3 #(.INIT(8'hE8)) lut_n2235 (.I0(x282), .I1(x283), .I2(x284), .O(n2235));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2236 (.I0(x273), .I1(x274), .I2(x275), .I3(n2232), .I4(n2233), .O(n2236));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2237 (.I0(x279), .I1(x280), .I2(x281), .I3(n2235), .I4(n2236), .O(n2237));
  LUT3 #(.INIT(8'h96)) lut_n2238 (.I0(n2226), .I1(n2229), .I2(n2230), .O(n2238));
  LUT3 #(.INIT(8'hE8)) lut_n2239 (.I0(n2234), .I1(n2237), .I2(n2238), .O(n2239));
  LUT3 #(.INIT(8'h96)) lut_n2240 (.I0(n2213), .I1(n2221), .I2(n2222), .O(n2240));
  LUT3 #(.INIT(8'hE8)) lut_n2241 (.I0(n2231), .I1(n2239), .I2(n2240), .O(n2241));
  LUT3 #(.INIT(8'h96)) lut_n2242 (.I0(n2185), .I1(n2203), .I2(n2204), .O(n2242));
  LUT3 #(.INIT(8'hE8)) lut_n2243 (.I0(n2223), .I1(n2241), .I2(n2242), .O(n2243));
  LUT3 #(.INIT(8'h96)) lut_n2244 (.I0(n2090), .I1(n2128), .I2(n2166), .O(n2244));
  LUT3 #(.INIT(8'hE8)) lut_n2245 (.I0(n2205), .I1(n2243), .I2(n2244), .O(n2245));
  LUT3 #(.INIT(8'hE8)) lut_n2246 (.I0(x288), .I1(x289), .I2(x290), .O(n2246));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2247 (.I0(x279), .I1(x280), .I2(x281), .I3(n2235), .I4(n2236), .O(n2247));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2248 (.I0(x285), .I1(x286), .I2(x287), .I3(n2246), .I4(n2247), .O(n2248));
  LUT3 #(.INIT(8'hE8)) lut_n2249 (.I0(x294), .I1(x295), .I2(x296), .O(n2249));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2250 (.I0(x285), .I1(x286), .I2(x287), .I3(n2246), .I4(n2247), .O(n2250));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2251 (.I0(x291), .I1(x292), .I2(x293), .I3(n2249), .I4(n2250), .O(n2251));
  LUT3 #(.INIT(8'h96)) lut_n2252 (.I0(n2234), .I1(n2237), .I2(n2238), .O(n2252));
  LUT3 #(.INIT(8'hE8)) lut_n2253 (.I0(n2248), .I1(n2251), .I2(n2252), .O(n2253));
  LUT3 #(.INIT(8'hE8)) lut_n2254 (.I0(x297), .I1(x298), .I2(x299), .O(n2254));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2255 (.I0(x291), .I1(x292), .I2(x293), .I3(n2249), .I4(n2250), .O(n2255));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2256 (.I0(x300), .I1(x301), .I2(x302), .I3(n2254), .I4(n2255), .O(n2256));
  LUT3 #(.INIT(8'hE8)) lut_n2257 (.I0(x306), .I1(x307), .I2(x308), .O(n2257));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2258 (.I0(x300), .I1(x301), .I2(x302), .I3(n2254), .I4(n2255), .O(n2258));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2259 (.I0(x303), .I1(x304), .I2(x305), .I3(n2257), .I4(n2258), .O(n2259));
  LUT3 #(.INIT(8'h96)) lut_n2260 (.I0(n2248), .I1(n2251), .I2(n2252), .O(n2260));
  LUT3 #(.INIT(8'hE8)) lut_n2261 (.I0(n2256), .I1(n2259), .I2(n2260), .O(n2261));
  LUT3 #(.INIT(8'h96)) lut_n2262 (.I0(n2231), .I1(n2239), .I2(n2240), .O(n2262));
  LUT3 #(.INIT(8'hE8)) lut_n2263 (.I0(n2253), .I1(n2261), .I2(n2262), .O(n2263));
  LUT3 #(.INIT(8'hE8)) lut_n2264 (.I0(x312), .I1(x313), .I2(x314), .O(n2264));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2265 (.I0(x303), .I1(x304), .I2(x305), .I3(n2257), .I4(n2258), .O(n2265));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2266 (.I0(x309), .I1(x310), .I2(x311), .I3(n2264), .I4(n2265), .O(n2266));
  LUT3 #(.INIT(8'hE8)) lut_n2267 (.I0(x318), .I1(x319), .I2(x320), .O(n2267));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2268 (.I0(x309), .I1(x310), .I2(x311), .I3(n2264), .I4(n2265), .O(n2268));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2269 (.I0(x315), .I1(x316), .I2(x317), .I3(n2267), .I4(n2268), .O(n2269));
  LUT3 #(.INIT(8'h96)) lut_n2270 (.I0(n2256), .I1(n2259), .I2(n2260), .O(n2270));
  LUT3 #(.INIT(8'hE8)) lut_n2271 (.I0(n2266), .I1(n2269), .I2(n2270), .O(n2271));
  LUT3 #(.INIT(8'hE8)) lut_n2272 (.I0(x324), .I1(x325), .I2(x326), .O(n2272));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2273 (.I0(x315), .I1(x316), .I2(x317), .I3(n2267), .I4(n2268), .O(n2273));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2274 (.I0(x321), .I1(x322), .I2(x323), .I3(n2272), .I4(n2273), .O(n2274));
  LUT3 #(.INIT(8'hE8)) lut_n2275 (.I0(x330), .I1(x331), .I2(x332), .O(n2275));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2276 (.I0(x321), .I1(x322), .I2(x323), .I3(n2272), .I4(n2273), .O(n2276));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2277 (.I0(x327), .I1(x328), .I2(x329), .I3(n2275), .I4(n2276), .O(n2277));
  LUT3 #(.INIT(8'h96)) lut_n2278 (.I0(n2266), .I1(n2269), .I2(n2270), .O(n2278));
  LUT3 #(.INIT(8'hE8)) lut_n2279 (.I0(n2274), .I1(n2277), .I2(n2278), .O(n2279));
  LUT3 #(.INIT(8'h96)) lut_n2280 (.I0(n2253), .I1(n2261), .I2(n2262), .O(n2280));
  LUT3 #(.INIT(8'hE8)) lut_n2281 (.I0(n2271), .I1(n2279), .I2(n2280), .O(n2281));
  LUT3 #(.INIT(8'h96)) lut_n2282 (.I0(n2223), .I1(n2241), .I2(n2242), .O(n2282));
  LUT3 #(.INIT(8'hE8)) lut_n2283 (.I0(n2263), .I1(n2281), .I2(n2282), .O(n2283));
  LUT3 #(.INIT(8'hE8)) lut_n2284 (.I0(x336), .I1(x337), .I2(x338), .O(n2284));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2285 (.I0(x327), .I1(x328), .I2(x329), .I3(n2275), .I4(n2276), .O(n2285));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2286 (.I0(x333), .I1(x334), .I2(x335), .I3(n2284), .I4(n2285), .O(n2286));
  LUT3 #(.INIT(8'hE8)) lut_n2287 (.I0(x342), .I1(x343), .I2(x344), .O(n2287));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2288 (.I0(x333), .I1(x334), .I2(x335), .I3(n2284), .I4(n2285), .O(n2288));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2289 (.I0(x339), .I1(x340), .I2(x341), .I3(n2287), .I4(n2288), .O(n2289));
  LUT3 #(.INIT(8'h96)) lut_n2290 (.I0(n2274), .I1(n2277), .I2(n2278), .O(n2290));
  LUT3 #(.INIT(8'hE8)) lut_n2291 (.I0(n2286), .I1(n2289), .I2(n2290), .O(n2291));
  LUT3 #(.INIT(8'hE8)) lut_n2292 (.I0(x348), .I1(x349), .I2(x350), .O(n2292));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2293 (.I0(x339), .I1(x340), .I2(x341), .I3(n2287), .I4(n2288), .O(n2293));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2294 (.I0(x345), .I1(x346), .I2(x347), .I3(n2292), .I4(n2293), .O(n2294));
  LUT3 #(.INIT(8'hE8)) lut_n2295 (.I0(x354), .I1(x355), .I2(x356), .O(n2295));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2296 (.I0(x345), .I1(x346), .I2(x347), .I3(n2292), .I4(n2293), .O(n2296));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2297 (.I0(x351), .I1(x352), .I2(x353), .I3(n2295), .I4(n2296), .O(n2297));
  LUT3 #(.INIT(8'h96)) lut_n2298 (.I0(n2286), .I1(n2289), .I2(n2290), .O(n2298));
  LUT3 #(.INIT(8'hE8)) lut_n2299 (.I0(n2294), .I1(n2297), .I2(n2298), .O(n2299));
  LUT3 #(.INIT(8'h96)) lut_n2300 (.I0(n2271), .I1(n2279), .I2(n2280), .O(n2300));
  LUT3 #(.INIT(8'hE8)) lut_n2301 (.I0(n2291), .I1(n2299), .I2(n2300), .O(n2301));
  LUT3 #(.INIT(8'hE8)) lut_n2302 (.I0(x360), .I1(x361), .I2(x362), .O(n2302));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2303 (.I0(x351), .I1(x352), .I2(x353), .I3(n2295), .I4(n2296), .O(n2303));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2304 (.I0(x357), .I1(x358), .I2(x359), .I3(n2302), .I4(n2303), .O(n2304));
  LUT3 #(.INIT(8'hE8)) lut_n2305 (.I0(x366), .I1(x367), .I2(x368), .O(n2305));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2306 (.I0(x357), .I1(x358), .I2(x359), .I3(n2302), .I4(n2303), .O(n2306));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2307 (.I0(x363), .I1(x364), .I2(x365), .I3(n2305), .I4(n2306), .O(n2307));
  LUT3 #(.INIT(8'h96)) lut_n2308 (.I0(n2294), .I1(n2297), .I2(n2298), .O(n2308));
  LUT3 #(.INIT(8'hE8)) lut_n2309 (.I0(n2304), .I1(n2307), .I2(n2308), .O(n2309));
  LUT3 #(.INIT(8'hE8)) lut_n2310 (.I0(x372), .I1(x373), .I2(x374), .O(n2310));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2311 (.I0(x363), .I1(x364), .I2(x365), .I3(n2305), .I4(n2306), .O(n2311));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2312 (.I0(x369), .I1(x370), .I2(x371), .I3(n2310), .I4(n2311), .O(n2312));
  LUT3 #(.INIT(8'hE8)) lut_n2313 (.I0(x378), .I1(x379), .I2(x380), .O(n2313));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2314 (.I0(x369), .I1(x370), .I2(x371), .I3(n2310), .I4(n2311), .O(n2314));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2315 (.I0(x375), .I1(x376), .I2(x377), .I3(n2313), .I4(n2314), .O(n2315));
  LUT3 #(.INIT(8'h96)) lut_n2316 (.I0(n2304), .I1(n2307), .I2(n2308), .O(n2316));
  LUT3 #(.INIT(8'hE8)) lut_n2317 (.I0(n2312), .I1(n2315), .I2(n2316), .O(n2317));
  LUT3 #(.INIT(8'h96)) lut_n2318 (.I0(n2291), .I1(n2299), .I2(n2300), .O(n2318));
  LUT3 #(.INIT(8'hE8)) lut_n2319 (.I0(n2309), .I1(n2317), .I2(n2318), .O(n2319));
  LUT3 #(.INIT(8'h96)) lut_n2320 (.I0(n2263), .I1(n2281), .I2(n2282), .O(n2320));
  LUT3 #(.INIT(8'hE8)) lut_n2321 (.I0(n2301), .I1(n2319), .I2(n2320), .O(n2321));
  LUT3 #(.INIT(8'h96)) lut_n2322 (.I0(n2205), .I1(n2243), .I2(n2244), .O(n2322));
  LUT3 #(.INIT(8'hE8)) lut_n2323 (.I0(n2283), .I1(n2321), .I2(n2322), .O(n2323));
  LUT3 #(.INIT(8'hE8)) lut_n2324 (.I0(n2167), .I1(n2245), .I2(n2323), .O(n2324));
  LUT3 #(.INIT(8'hE8)) lut_n2325 (.I0(x384), .I1(x385), .I2(x386), .O(n2325));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2326 (.I0(x375), .I1(x376), .I2(x377), .I3(n2313), .I4(n2314), .O(n2326));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2327 (.I0(x381), .I1(x382), .I2(x383), .I3(n2325), .I4(n2326), .O(n2327));
  LUT3 #(.INIT(8'hE8)) lut_n2328 (.I0(x390), .I1(x391), .I2(x392), .O(n2328));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2329 (.I0(x381), .I1(x382), .I2(x383), .I3(n2325), .I4(n2326), .O(n2329));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2330 (.I0(x387), .I1(x388), .I2(x389), .I3(n2328), .I4(n2329), .O(n2330));
  LUT3 #(.INIT(8'h96)) lut_n2331 (.I0(n2312), .I1(n2315), .I2(n2316), .O(n2331));
  LUT3 #(.INIT(8'hE8)) lut_n2332 (.I0(n2327), .I1(n2330), .I2(n2331), .O(n2332));
  LUT3 #(.INIT(8'hE8)) lut_n2333 (.I0(x396), .I1(x397), .I2(x398), .O(n2333));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2334 (.I0(x387), .I1(x388), .I2(x389), .I3(n2328), .I4(n2329), .O(n2334));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2335 (.I0(x393), .I1(x394), .I2(x395), .I3(n2333), .I4(n2334), .O(n2335));
  LUT3 #(.INIT(8'hE8)) lut_n2336 (.I0(x402), .I1(x403), .I2(x404), .O(n2336));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2337 (.I0(x393), .I1(x394), .I2(x395), .I3(n2333), .I4(n2334), .O(n2337));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2338 (.I0(x399), .I1(x400), .I2(x401), .I3(n2336), .I4(n2337), .O(n2338));
  LUT3 #(.INIT(8'h96)) lut_n2339 (.I0(n2327), .I1(n2330), .I2(n2331), .O(n2339));
  LUT3 #(.INIT(8'hE8)) lut_n2340 (.I0(n2335), .I1(n2338), .I2(n2339), .O(n2340));
  LUT3 #(.INIT(8'h96)) lut_n2341 (.I0(n2309), .I1(n2317), .I2(n2318), .O(n2341));
  LUT3 #(.INIT(8'hE8)) lut_n2342 (.I0(n2332), .I1(n2340), .I2(n2341), .O(n2342));
  LUT3 #(.INIT(8'hE8)) lut_n2343 (.I0(x408), .I1(x409), .I2(x410), .O(n2343));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2344 (.I0(x399), .I1(x400), .I2(x401), .I3(n2336), .I4(n2337), .O(n2344));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2345 (.I0(x405), .I1(x406), .I2(x407), .I3(n2343), .I4(n2344), .O(n2345));
  LUT3 #(.INIT(8'hE8)) lut_n2346 (.I0(x414), .I1(x415), .I2(x416), .O(n2346));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2347 (.I0(x405), .I1(x406), .I2(x407), .I3(n2343), .I4(n2344), .O(n2347));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2348 (.I0(x411), .I1(x412), .I2(x413), .I3(n2346), .I4(n2347), .O(n2348));
  LUT3 #(.INIT(8'h96)) lut_n2349 (.I0(n2335), .I1(n2338), .I2(n2339), .O(n2349));
  LUT3 #(.INIT(8'hE8)) lut_n2350 (.I0(n2345), .I1(n2348), .I2(n2349), .O(n2350));
  LUT3 #(.INIT(8'hE8)) lut_n2351 (.I0(x420), .I1(x421), .I2(x422), .O(n2351));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2352 (.I0(x411), .I1(x412), .I2(x413), .I3(n2346), .I4(n2347), .O(n2352));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2353 (.I0(x417), .I1(x418), .I2(x419), .I3(n2351), .I4(n2352), .O(n2353));
  LUT3 #(.INIT(8'hE8)) lut_n2354 (.I0(x426), .I1(x427), .I2(x428), .O(n2354));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2355 (.I0(x417), .I1(x418), .I2(x419), .I3(n2351), .I4(n2352), .O(n2355));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2356 (.I0(x423), .I1(x424), .I2(x425), .I3(n2354), .I4(n2355), .O(n2356));
  LUT3 #(.INIT(8'h96)) lut_n2357 (.I0(n2345), .I1(n2348), .I2(n2349), .O(n2357));
  LUT3 #(.INIT(8'hE8)) lut_n2358 (.I0(n2353), .I1(n2356), .I2(n2357), .O(n2358));
  LUT3 #(.INIT(8'h96)) lut_n2359 (.I0(n2332), .I1(n2340), .I2(n2341), .O(n2359));
  LUT3 #(.INIT(8'hE8)) lut_n2360 (.I0(n2350), .I1(n2358), .I2(n2359), .O(n2360));
  LUT3 #(.INIT(8'h96)) lut_n2361 (.I0(n2301), .I1(n2319), .I2(n2320), .O(n2361));
  LUT3 #(.INIT(8'hE8)) lut_n2362 (.I0(n2342), .I1(n2360), .I2(n2361), .O(n2362));
  LUT3 #(.INIT(8'hE8)) lut_n2363 (.I0(x432), .I1(x433), .I2(x434), .O(n2363));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2364 (.I0(x423), .I1(x424), .I2(x425), .I3(n2354), .I4(n2355), .O(n2364));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2365 (.I0(x429), .I1(x430), .I2(x431), .I3(n2363), .I4(n2364), .O(n2365));
  LUT3 #(.INIT(8'hE8)) lut_n2366 (.I0(x438), .I1(x439), .I2(x440), .O(n2366));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2367 (.I0(x429), .I1(x430), .I2(x431), .I3(n2363), .I4(n2364), .O(n2367));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2368 (.I0(x435), .I1(x436), .I2(x437), .I3(n2366), .I4(n2367), .O(n2368));
  LUT3 #(.INIT(8'h96)) lut_n2369 (.I0(n2353), .I1(n2356), .I2(n2357), .O(n2369));
  LUT3 #(.INIT(8'hE8)) lut_n2370 (.I0(n2365), .I1(n2368), .I2(n2369), .O(n2370));
  LUT3 #(.INIT(8'hE8)) lut_n2371 (.I0(x444), .I1(x445), .I2(x446), .O(n2371));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2372 (.I0(x435), .I1(x436), .I2(x437), .I3(n2366), .I4(n2367), .O(n2372));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2373 (.I0(x441), .I1(x442), .I2(x443), .I3(n2371), .I4(n2372), .O(n2373));
  LUT3 #(.INIT(8'hE8)) lut_n2374 (.I0(x450), .I1(x451), .I2(x452), .O(n2374));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2375 (.I0(x441), .I1(x442), .I2(x443), .I3(n2371), .I4(n2372), .O(n2375));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2376 (.I0(x447), .I1(x448), .I2(x449), .I3(n2374), .I4(n2375), .O(n2376));
  LUT3 #(.INIT(8'h96)) lut_n2377 (.I0(n2365), .I1(n2368), .I2(n2369), .O(n2377));
  LUT3 #(.INIT(8'hE8)) lut_n2378 (.I0(n2373), .I1(n2376), .I2(n2377), .O(n2378));
  LUT3 #(.INIT(8'h96)) lut_n2379 (.I0(n2350), .I1(n2358), .I2(n2359), .O(n2379));
  LUT3 #(.INIT(8'hE8)) lut_n2380 (.I0(n2370), .I1(n2378), .I2(n2379), .O(n2380));
  LUT3 #(.INIT(8'hE8)) lut_n2381 (.I0(x456), .I1(x457), .I2(x458), .O(n2381));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2382 (.I0(x447), .I1(x448), .I2(x449), .I3(n2374), .I4(n2375), .O(n2382));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2383 (.I0(x453), .I1(x454), .I2(x455), .I3(n2381), .I4(n2382), .O(n2383));
  LUT3 #(.INIT(8'hE8)) lut_n2384 (.I0(x462), .I1(x463), .I2(x464), .O(n2384));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2385 (.I0(x453), .I1(x454), .I2(x455), .I3(n2381), .I4(n2382), .O(n2385));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2386 (.I0(x459), .I1(x460), .I2(x461), .I3(n2384), .I4(n2385), .O(n2386));
  LUT3 #(.INIT(8'h96)) lut_n2387 (.I0(n2373), .I1(n2376), .I2(n2377), .O(n2387));
  LUT3 #(.INIT(8'hE8)) lut_n2388 (.I0(n2383), .I1(n2386), .I2(n2387), .O(n2388));
  LUT3 #(.INIT(8'hE8)) lut_n2389 (.I0(x468), .I1(x469), .I2(x470), .O(n2389));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2390 (.I0(x459), .I1(x460), .I2(x461), .I3(n2384), .I4(n2385), .O(n2390));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2391 (.I0(x465), .I1(x466), .I2(x467), .I3(n2389), .I4(n2390), .O(n2391));
  LUT3 #(.INIT(8'hE8)) lut_n2392 (.I0(x474), .I1(x475), .I2(x476), .O(n2392));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2393 (.I0(x465), .I1(x466), .I2(x467), .I3(n2389), .I4(n2390), .O(n2393));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2394 (.I0(x471), .I1(x472), .I2(x473), .I3(n2392), .I4(n2393), .O(n2394));
  LUT3 #(.INIT(8'h96)) lut_n2395 (.I0(n2383), .I1(n2386), .I2(n2387), .O(n2395));
  LUT3 #(.INIT(8'hE8)) lut_n2396 (.I0(n2391), .I1(n2394), .I2(n2395), .O(n2396));
  LUT3 #(.INIT(8'h96)) lut_n2397 (.I0(n2370), .I1(n2378), .I2(n2379), .O(n2397));
  LUT3 #(.INIT(8'hE8)) lut_n2398 (.I0(n2388), .I1(n2396), .I2(n2397), .O(n2398));
  LUT3 #(.INIT(8'h96)) lut_n2399 (.I0(n2342), .I1(n2360), .I2(n2361), .O(n2399));
  LUT3 #(.INIT(8'hE8)) lut_n2400 (.I0(n2380), .I1(n2398), .I2(n2399), .O(n2400));
  LUT3 #(.INIT(8'h96)) lut_n2401 (.I0(n2283), .I1(n2321), .I2(n2322), .O(n2401));
  LUT3 #(.INIT(8'hE8)) lut_n2402 (.I0(n2362), .I1(n2400), .I2(n2401), .O(n2402));
  LUT3 #(.INIT(8'hE8)) lut_n2403 (.I0(x480), .I1(x481), .I2(x482), .O(n2403));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2404 (.I0(x471), .I1(x472), .I2(x473), .I3(n2392), .I4(n2393), .O(n2404));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2405 (.I0(x477), .I1(x478), .I2(x479), .I3(n2403), .I4(n2404), .O(n2405));
  LUT3 #(.INIT(8'hE8)) lut_n2406 (.I0(x486), .I1(x487), .I2(x488), .O(n2406));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2407 (.I0(x477), .I1(x478), .I2(x479), .I3(n2403), .I4(n2404), .O(n2407));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2408 (.I0(x483), .I1(x484), .I2(x485), .I3(n2406), .I4(n2407), .O(n2408));
  LUT3 #(.INIT(8'h96)) lut_n2409 (.I0(n2391), .I1(n2394), .I2(n2395), .O(n2409));
  LUT3 #(.INIT(8'hE8)) lut_n2410 (.I0(n2405), .I1(n2408), .I2(n2409), .O(n2410));
  LUT3 #(.INIT(8'hE8)) lut_n2411 (.I0(x492), .I1(x493), .I2(x494), .O(n2411));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2412 (.I0(x483), .I1(x484), .I2(x485), .I3(n2406), .I4(n2407), .O(n2412));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2413 (.I0(x489), .I1(x490), .I2(x491), .I3(n2411), .I4(n2412), .O(n2413));
  LUT3 #(.INIT(8'hE8)) lut_n2414 (.I0(x498), .I1(x499), .I2(x500), .O(n2414));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2415 (.I0(x489), .I1(x490), .I2(x491), .I3(n2411), .I4(n2412), .O(n2415));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2416 (.I0(x495), .I1(x496), .I2(x497), .I3(n2414), .I4(n2415), .O(n2416));
  LUT3 #(.INIT(8'h96)) lut_n2417 (.I0(n2405), .I1(n2408), .I2(n2409), .O(n2417));
  LUT3 #(.INIT(8'hE8)) lut_n2418 (.I0(n2413), .I1(n2416), .I2(n2417), .O(n2418));
  LUT3 #(.INIT(8'h96)) lut_n2419 (.I0(n2388), .I1(n2396), .I2(n2397), .O(n2419));
  LUT3 #(.INIT(8'hE8)) lut_n2420 (.I0(n2410), .I1(n2418), .I2(n2419), .O(n2420));
  LUT3 #(.INIT(8'hE8)) lut_n2421 (.I0(x504), .I1(x505), .I2(x506), .O(n2421));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2422 (.I0(x495), .I1(x496), .I2(x497), .I3(n2414), .I4(n2415), .O(n2422));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2423 (.I0(x501), .I1(x502), .I2(x503), .I3(n2421), .I4(n2422), .O(n2423));
  LUT3 #(.INIT(8'hE8)) lut_n2424 (.I0(x510), .I1(x511), .I2(x512), .O(n2424));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2425 (.I0(x501), .I1(x502), .I2(x503), .I3(n2421), .I4(n2422), .O(n2425));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2426 (.I0(x507), .I1(x508), .I2(x509), .I3(n2424), .I4(n2425), .O(n2426));
  LUT3 #(.INIT(8'h96)) lut_n2427 (.I0(n2413), .I1(n2416), .I2(n2417), .O(n2427));
  LUT3 #(.INIT(8'hE8)) lut_n2428 (.I0(n2423), .I1(n2426), .I2(n2427), .O(n2428));
  LUT3 #(.INIT(8'hE8)) lut_n2429 (.I0(x516), .I1(x517), .I2(x518), .O(n2429));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2430 (.I0(x507), .I1(x508), .I2(x509), .I3(n2424), .I4(n2425), .O(n2430));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2431 (.I0(x513), .I1(x514), .I2(x515), .I3(n2429), .I4(n2430), .O(n2431));
  LUT3 #(.INIT(8'hE8)) lut_n2432 (.I0(x522), .I1(x523), .I2(x524), .O(n2432));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2433 (.I0(x513), .I1(x514), .I2(x515), .I3(n2429), .I4(n2430), .O(n2433));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2434 (.I0(x519), .I1(x520), .I2(x521), .I3(n2432), .I4(n2433), .O(n2434));
  LUT3 #(.INIT(8'h96)) lut_n2435 (.I0(n2423), .I1(n2426), .I2(n2427), .O(n2435));
  LUT3 #(.INIT(8'hE8)) lut_n2436 (.I0(n2431), .I1(n2434), .I2(n2435), .O(n2436));
  LUT3 #(.INIT(8'h96)) lut_n2437 (.I0(n2410), .I1(n2418), .I2(n2419), .O(n2437));
  LUT3 #(.INIT(8'hE8)) lut_n2438 (.I0(n2428), .I1(n2436), .I2(n2437), .O(n2438));
  LUT3 #(.INIT(8'h96)) lut_n2439 (.I0(n2380), .I1(n2398), .I2(n2399), .O(n2439));
  LUT3 #(.INIT(8'hE8)) lut_n2440 (.I0(n2420), .I1(n2438), .I2(n2439), .O(n2440));
  LUT3 #(.INIT(8'hE8)) lut_n2441 (.I0(x528), .I1(x529), .I2(x530), .O(n2441));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2442 (.I0(x519), .I1(x520), .I2(x521), .I3(n2432), .I4(n2433), .O(n2442));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2443 (.I0(x525), .I1(x526), .I2(x527), .I3(n2441), .I4(n2442), .O(n2443));
  LUT3 #(.INIT(8'hE8)) lut_n2444 (.I0(x534), .I1(x535), .I2(x536), .O(n2444));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2445 (.I0(x525), .I1(x526), .I2(x527), .I3(n2441), .I4(n2442), .O(n2445));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2446 (.I0(x531), .I1(x532), .I2(x533), .I3(n2444), .I4(n2445), .O(n2446));
  LUT3 #(.INIT(8'h96)) lut_n2447 (.I0(n2431), .I1(n2434), .I2(n2435), .O(n2447));
  LUT3 #(.INIT(8'hE8)) lut_n2448 (.I0(n2443), .I1(n2446), .I2(n2447), .O(n2448));
  LUT3 #(.INIT(8'hE8)) lut_n2449 (.I0(x540), .I1(x541), .I2(x542), .O(n2449));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2450 (.I0(x531), .I1(x532), .I2(x533), .I3(n2444), .I4(n2445), .O(n2450));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2451 (.I0(x537), .I1(x538), .I2(x539), .I3(n2449), .I4(n2450), .O(n2451));
  LUT3 #(.INIT(8'hE8)) lut_n2452 (.I0(x546), .I1(x547), .I2(x548), .O(n2452));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2453 (.I0(x537), .I1(x538), .I2(x539), .I3(n2449), .I4(n2450), .O(n2453));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2454 (.I0(x543), .I1(x544), .I2(x545), .I3(n2452), .I4(n2453), .O(n2454));
  LUT3 #(.INIT(8'h96)) lut_n2455 (.I0(n2443), .I1(n2446), .I2(n2447), .O(n2455));
  LUT3 #(.INIT(8'hE8)) lut_n2456 (.I0(n2451), .I1(n2454), .I2(n2455), .O(n2456));
  LUT3 #(.INIT(8'h96)) lut_n2457 (.I0(n2428), .I1(n2436), .I2(n2437), .O(n2457));
  LUT3 #(.INIT(8'hE8)) lut_n2458 (.I0(n2448), .I1(n2456), .I2(n2457), .O(n2458));
  LUT3 #(.INIT(8'hE8)) lut_n2459 (.I0(x552), .I1(x553), .I2(x554), .O(n2459));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2460 (.I0(x543), .I1(x544), .I2(x545), .I3(n2452), .I4(n2453), .O(n2460));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2461 (.I0(x549), .I1(x550), .I2(x551), .I3(n2459), .I4(n2460), .O(n2461));
  LUT3 #(.INIT(8'hE8)) lut_n2462 (.I0(x558), .I1(x559), .I2(x560), .O(n2462));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2463 (.I0(x549), .I1(x550), .I2(x551), .I3(n2459), .I4(n2460), .O(n2463));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2464 (.I0(x555), .I1(x556), .I2(x557), .I3(n2462), .I4(n2463), .O(n2464));
  LUT3 #(.INIT(8'h96)) lut_n2465 (.I0(n2451), .I1(n2454), .I2(n2455), .O(n2465));
  LUT3 #(.INIT(8'hE8)) lut_n2466 (.I0(n2461), .I1(n2464), .I2(n2465), .O(n2466));
  LUT3 #(.INIT(8'hE8)) lut_n2467 (.I0(x564), .I1(x565), .I2(x566), .O(n2467));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2468 (.I0(x555), .I1(x556), .I2(x557), .I3(n2462), .I4(n2463), .O(n2468));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2469 (.I0(x561), .I1(x562), .I2(x563), .I3(n2467), .I4(n2468), .O(n2469));
  LUT3 #(.INIT(8'hE8)) lut_n2470 (.I0(x570), .I1(x571), .I2(x572), .O(n2470));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2471 (.I0(x561), .I1(x562), .I2(x563), .I3(n2467), .I4(n2468), .O(n2471));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2472 (.I0(x567), .I1(x568), .I2(x569), .I3(n2470), .I4(n2471), .O(n2472));
  LUT3 #(.INIT(8'h96)) lut_n2473 (.I0(n2461), .I1(n2464), .I2(n2465), .O(n2473));
  LUT3 #(.INIT(8'hE8)) lut_n2474 (.I0(n2469), .I1(n2472), .I2(n2473), .O(n2474));
  LUT3 #(.INIT(8'h96)) lut_n2475 (.I0(n2448), .I1(n2456), .I2(n2457), .O(n2475));
  LUT3 #(.INIT(8'hE8)) lut_n2476 (.I0(n2466), .I1(n2474), .I2(n2475), .O(n2476));
  LUT3 #(.INIT(8'h96)) lut_n2477 (.I0(n2420), .I1(n2438), .I2(n2439), .O(n2477));
  LUT3 #(.INIT(8'hE8)) lut_n2478 (.I0(n2458), .I1(n2476), .I2(n2477), .O(n2478));
  LUT3 #(.INIT(8'h96)) lut_n2479 (.I0(n2362), .I1(n2400), .I2(n2401), .O(n2479));
  LUT3 #(.INIT(8'hE8)) lut_n2480 (.I0(n2440), .I1(n2478), .I2(n2479), .O(n2480));
  LUT3 #(.INIT(8'h96)) lut_n2481 (.I0(n2167), .I1(n2245), .I2(n2323), .O(n2481));
  LUT3 #(.INIT(8'hE8)) lut_n2482 (.I0(n2402), .I1(n2480), .I2(n2481), .O(n2482));
  LUT3 #(.INIT(8'hE8)) lut_n2483 (.I0(x576), .I1(x577), .I2(x578), .O(n2483));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2484 (.I0(x567), .I1(x568), .I2(x569), .I3(n2470), .I4(n2471), .O(n2484));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2485 (.I0(x573), .I1(x574), .I2(x575), .I3(n2483), .I4(n2484), .O(n2485));
  LUT3 #(.INIT(8'hE8)) lut_n2486 (.I0(x582), .I1(x583), .I2(x584), .O(n2486));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2487 (.I0(x573), .I1(x574), .I2(x575), .I3(n2483), .I4(n2484), .O(n2487));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2488 (.I0(x579), .I1(x580), .I2(x581), .I3(n2486), .I4(n2487), .O(n2488));
  LUT3 #(.INIT(8'h96)) lut_n2489 (.I0(n2469), .I1(n2472), .I2(n2473), .O(n2489));
  LUT3 #(.INIT(8'hE8)) lut_n2490 (.I0(n2485), .I1(n2488), .I2(n2489), .O(n2490));
  LUT3 #(.INIT(8'hE8)) lut_n2491 (.I0(x588), .I1(x589), .I2(x590), .O(n2491));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2492 (.I0(x579), .I1(x580), .I2(x581), .I3(n2486), .I4(n2487), .O(n2492));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2493 (.I0(x585), .I1(x586), .I2(x587), .I3(n2491), .I4(n2492), .O(n2493));
  LUT3 #(.INIT(8'hE8)) lut_n2494 (.I0(x594), .I1(x595), .I2(x596), .O(n2494));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2495 (.I0(x585), .I1(x586), .I2(x587), .I3(n2491), .I4(n2492), .O(n2495));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2496 (.I0(x591), .I1(x592), .I2(x593), .I3(n2494), .I4(n2495), .O(n2496));
  LUT3 #(.INIT(8'h96)) lut_n2497 (.I0(n2485), .I1(n2488), .I2(n2489), .O(n2497));
  LUT3 #(.INIT(8'hE8)) lut_n2498 (.I0(n2493), .I1(n2496), .I2(n2497), .O(n2498));
  LUT3 #(.INIT(8'h96)) lut_n2499 (.I0(n2466), .I1(n2474), .I2(n2475), .O(n2499));
  LUT3 #(.INIT(8'hE8)) lut_n2500 (.I0(n2490), .I1(n2498), .I2(n2499), .O(n2500));
  LUT3 #(.INIT(8'hE8)) lut_n2501 (.I0(x600), .I1(x601), .I2(x602), .O(n2501));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2502 (.I0(x591), .I1(x592), .I2(x593), .I3(n2494), .I4(n2495), .O(n2502));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2503 (.I0(x597), .I1(x598), .I2(x599), .I3(n2501), .I4(n2502), .O(n2503));
  LUT3 #(.INIT(8'hE8)) lut_n2504 (.I0(x606), .I1(x607), .I2(x608), .O(n2504));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2505 (.I0(x597), .I1(x598), .I2(x599), .I3(n2501), .I4(n2502), .O(n2505));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2506 (.I0(x603), .I1(x604), .I2(x605), .I3(n2504), .I4(n2505), .O(n2506));
  LUT3 #(.INIT(8'h96)) lut_n2507 (.I0(n2493), .I1(n2496), .I2(n2497), .O(n2507));
  LUT3 #(.INIT(8'hE8)) lut_n2508 (.I0(n2503), .I1(n2506), .I2(n2507), .O(n2508));
  LUT3 #(.INIT(8'hE8)) lut_n2509 (.I0(x612), .I1(x613), .I2(x614), .O(n2509));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2510 (.I0(x603), .I1(x604), .I2(x605), .I3(n2504), .I4(n2505), .O(n2510));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2511 (.I0(x609), .I1(x610), .I2(x611), .I3(n2509), .I4(n2510), .O(n2511));
  LUT3 #(.INIT(8'hE8)) lut_n2512 (.I0(x618), .I1(x619), .I2(x620), .O(n2512));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2513 (.I0(x609), .I1(x610), .I2(x611), .I3(n2509), .I4(n2510), .O(n2513));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2514 (.I0(x615), .I1(x616), .I2(x617), .I3(n2512), .I4(n2513), .O(n2514));
  LUT3 #(.INIT(8'h96)) lut_n2515 (.I0(n2503), .I1(n2506), .I2(n2507), .O(n2515));
  LUT3 #(.INIT(8'hE8)) lut_n2516 (.I0(n2511), .I1(n2514), .I2(n2515), .O(n2516));
  LUT3 #(.INIT(8'h96)) lut_n2517 (.I0(n2490), .I1(n2498), .I2(n2499), .O(n2517));
  LUT3 #(.INIT(8'hE8)) lut_n2518 (.I0(n2508), .I1(n2516), .I2(n2517), .O(n2518));
  LUT3 #(.INIT(8'h96)) lut_n2519 (.I0(n2458), .I1(n2476), .I2(n2477), .O(n2519));
  LUT3 #(.INIT(8'hE8)) lut_n2520 (.I0(n2500), .I1(n2518), .I2(n2519), .O(n2520));
  LUT3 #(.INIT(8'hE8)) lut_n2521 (.I0(x624), .I1(x625), .I2(x626), .O(n2521));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2522 (.I0(x615), .I1(x616), .I2(x617), .I3(n2512), .I4(n2513), .O(n2522));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2523 (.I0(x621), .I1(x622), .I2(x623), .I3(n2521), .I4(n2522), .O(n2523));
  LUT3 #(.INIT(8'hE8)) lut_n2524 (.I0(x630), .I1(x631), .I2(x632), .O(n2524));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2525 (.I0(x621), .I1(x622), .I2(x623), .I3(n2521), .I4(n2522), .O(n2525));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2526 (.I0(x627), .I1(x628), .I2(x629), .I3(n2524), .I4(n2525), .O(n2526));
  LUT3 #(.INIT(8'h96)) lut_n2527 (.I0(n2511), .I1(n2514), .I2(n2515), .O(n2527));
  LUT3 #(.INIT(8'hE8)) lut_n2528 (.I0(n2523), .I1(n2526), .I2(n2527), .O(n2528));
  LUT3 #(.INIT(8'hE8)) lut_n2529 (.I0(x636), .I1(x637), .I2(x638), .O(n2529));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2530 (.I0(x627), .I1(x628), .I2(x629), .I3(n2524), .I4(n2525), .O(n2530));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2531 (.I0(x633), .I1(x634), .I2(x635), .I3(n2529), .I4(n2530), .O(n2531));
  LUT3 #(.INIT(8'hE8)) lut_n2532 (.I0(x642), .I1(x643), .I2(x644), .O(n2532));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2533 (.I0(x633), .I1(x634), .I2(x635), .I3(n2529), .I4(n2530), .O(n2533));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2534 (.I0(x639), .I1(x640), .I2(x641), .I3(n2532), .I4(n2533), .O(n2534));
  LUT3 #(.INIT(8'h96)) lut_n2535 (.I0(n2523), .I1(n2526), .I2(n2527), .O(n2535));
  LUT3 #(.INIT(8'hE8)) lut_n2536 (.I0(n2531), .I1(n2534), .I2(n2535), .O(n2536));
  LUT3 #(.INIT(8'h96)) lut_n2537 (.I0(n2508), .I1(n2516), .I2(n2517), .O(n2537));
  LUT3 #(.INIT(8'hE8)) lut_n2538 (.I0(n2528), .I1(n2536), .I2(n2537), .O(n2538));
  LUT3 #(.INIT(8'hE8)) lut_n2539 (.I0(x648), .I1(x649), .I2(x650), .O(n2539));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2540 (.I0(x639), .I1(x640), .I2(x641), .I3(n2532), .I4(n2533), .O(n2540));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2541 (.I0(x645), .I1(x646), .I2(x647), .I3(n2539), .I4(n2540), .O(n2541));
  LUT3 #(.INIT(8'hE8)) lut_n2542 (.I0(x654), .I1(x655), .I2(x656), .O(n2542));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2543 (.I0(x645), .I1(x646), .I2(x647), .I3(n2539), .I4(n2540), .O(n2543));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2544 (.I0(x651), .I1(x652), .I2(x653), .I3(n2542), .I4(n2543), .O(n2544));
  LUT3 #(.INIT(8'h96)) lut_n2545 (.I0(n2531), .I1(n2534), .I2(n2535), .O(n2545));
  LUT3 #(.INIT(8'hE8)) lut_n2546 (.I0(n2541), .I1(n2544), .I2(n2545), .O(n2546));
  LUT3 #(.INIT(8'hE8)) lut_n2547 (.I0(x660), .I1(x661), .I2(x662), .O(n2547));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2548 (.I0(x651), .I1(x652), .I2(x653), .I3(n2542), .I4(n2543), .O(n2548));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2549 (.I0(x657), .I1(x658), .I2(x659), .I3(n2547), .I4(n2548), .O(n2549));
  LUT3 #(.INIT(8'hE8)) lut_n2550 (.I0(x666), .I1(x667), .I2(x668), .O(n2550));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2551 (.I0(x657), .I1(x658), .I2(x659), .I3(n2547), .I4(n2548), .O(n2551));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2552 (.I0(x663), .I1(x664), .I2(x665), .I3(n2550), .I4(n2551), .O(n2552));
  LUT3 #(.INIT(8'h96)) lut_n2553 (.I0(n2541), .I1(n2544), .I2(n2545), .O(n2553));
  LUT3 #(.INIT(8'hE8)) lut_n2554 (.I0(n2549), .I1(n2552), .I2(n2553), .O(n2554));
  LUT3 #(.INIT(8'h96)) lut_n2555 (.I0(n2528), .I1(n2536), .I2(n2537), .O(n2555));
  LUT3 #(.INIT(8'hE8)) lut_n2556 (.I0(n2546), .I1(n2554), .I2(n2555), .O(n2556));
  LUT3 #(.INIT(8'h96)) lut_n2557 (.I0(n2500), .I1(n2518), .I2(n2519), .O(n2557));
  LUT3 #(.INIT(8'hE8)) lut_n2558 (.I0(n2538), .I1(n2556), .I2(n2557), .O(n2558));
  LUT3 #(.INIT(8'h96)) lut_n2559 (.I0(n2440), .I1(n2478), .I2(n2479), .O(n2559));
  LUT3 #(.INIT(8'hE8)) lut_n2560 (.I0(n2520), .I1(n2558), .I2(n2559), .O(n2560));
  LUT3 #(.INIT(8'hE8)) lut_n2561 (.I0(x672), .I1(x673), .I2(x674), .O(n2561));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2562 (.I0(x663), .I1(x664), .I2(x665), .I3(n2550), .I4(n2551), .O(n2562));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2563 (.I0(x669), .I1(x670), .I2(x671), .I3(n2561), .I4(n2562), .O(n2563));
  LUT3 #(.INIT(8'hE8)) lut_n2564 (.I0(x678), .I1(x679), .I2(x680), .O(n2564));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2565 (.I0(x669), .I1(x670), .I2(x671), .I3(n2561), .I4(n2562), .O(n2565));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2566 (.I0(x675), .I1(x676), .I2(x677), .I3(n2564), .I4(n2565), .O(n2566));
  LUT3 #(.INIT(8'h96)) lut_n2567 (.I0(n2549), .I1(n2552), .I2(n2553), .O(n2567));
  LUT3 #(.INIT(8'hE8)) lut_n2568 (.I0(n2563), .I1(n2566), .I2(n2567), .O(n2568));
  LUT3 #(.INIT(8'hE8)) lut_n2569 (.I0(x684), .I1(x685), .I2(x686), .O(n2569));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2570 (.I0(x675), .I1(x676), .I2(x677), .I3(n2564), .I4(n2565), .O(n2570));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2571 (.I0(x681), .I1(x682), .I2(x683), .I3(n2569), .I4(n2570), .O(n2571));
  LUT3 #(.INIT(8'hE8)) lut_n2572 (.I0(x690), .I1(x691), .I2(x692), .O(n2572));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2573 (.I0(x681), .I1(x682), .I2(x683), .I3(n2569), .I4(n2570), .O(n2573));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2574 (.I0(x687), .I1(x688), .I2(x689), .I3(n2572), .I4(n2573), .O(n2574));
  LUT3 #(.INIT(8'h96)) lut_n2575 (.I0(n2563), .I1(n2566), .I2(n2567), .O(n2575));
  LUT3 #(.INIT(8'hE8)) lut_n2576 (.I0(n2571), .I1(n2574), .I2(n2575), .O(n2576));
  LUT3 #(.INIT(8'h96)) lut_n2577 (.I0(n2546), .I1(n2554), .I2(n2555), .O(n2577));
  LUT3 #(.INIT(8'hE8)) lut_n2578 (.I0(n2568), .I1(n2576), .I2(n2577), .O(n2578));
  LUT3 #(.INIT(8'hE8)) lut_n2579 (.I0(x696), .I1(x697), .I2(x698), .O(n2579));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2580 (.I0(x687), .I1(x688), .I2(x689), .I3(n2572), .I4(n2573), .O(n2580));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2581 (.I0(x693), .I1(x694), .I2(x695), .I3(n2579), .I4(n2580), .O(n2581));
  LUT3 #(.INIT(8'hE8)) lut_n2582 (.I0(x702), .I1(x703), .I2(x704), .O(n2582));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2583 (.I0(x693), .I1(x694), .I2(x695), .I3(n2579), .I4(n2580), .O(n2583));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2584 (.I0(x699), .I1(x700), .I2(x701), .I3(n2582), .I4(n2583), .O(n2584));
  LUT3 #(.INIT(8'h96)) lut_n2585 (.I0(n2571), .I1(n2574), .I2(n2575), .O(n2585));
  LUT3 #(.INIT(8'hE8)) lut_n2586 (.I0(n2581), .I1(n2584), .I2(n2585), .O(n2586));
  LUT3 #(.INIT(8'hE8)) lut_n2587 (.I0(x708), .I1(x709), .I2(x710), .O(n2587));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2588 (.I0(x699), .I1(x700), .I2(x701), .I3(n2582), .I4(n2583), .O(n2588));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2589 (.I0(x705), .I1(x706), .I2(x707), .I3(n2587), .I4(n2588), .O(n2589));
  LUT3 #(.INIT(8'hE8)) lut_n2590 (.I0(x714), .I1(x715), .I2(x716), .O(n2590));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2591 (.I0(x705), .I1(x706), .I2(x707), .I3(n2587), .I4(n2588), .O(n2591));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2592 (.I0(x711), .I1(x712), .I2(x713), .I3(n2590), .I4(n2591), .O(n2592));
  LUT3 #(.INIT(8'h96)) lut_n2593 (.I0(n2581), .I1(n2584), .I2(n2585), .O(n2593));
  LUT3 #(.INIT(8'hE8)) lut_n2594 (.I0(n2589), .I1(n2592), .I2(n2593), .O(n2594));
  LUT3 #(.INIT(8'h96)) lut_n2595 (.I0(n2568), .I1(n2576), .I2(n2577), .O(n2595));
  LUT3 #(.INIT(8'hE8)) lut_n2596 (.I0(n2586), .I1(n2594), .I2(n2595), .O(n2596));
  LUT3 #(.INIT(8'h96)) lut_n2597 (.I0(n2538), .I1(n2556), .I2(n2557), .O(n2597));
  LUT3 #(.INIT(8'hE8)) lut_n2598 (.I0(n2578), .I1(n2596), .I2(n2597), .O(n2598));
  LUT3 #(.INIT(8'hE8)) lut_n2599 (.I0(x720), .I1(x721), .I2(x722), .O(n2599));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2600 (.I0(x711), .I1(x712), .I2(x713), .I3(n2590), .I4(n2591), .O(n2600));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2601 (.I0(x717), .I1(x718), .I2(x719), .I3(n2599), .I4(n2600), .O(n2601));
  LUT3 #(.INIT(8'hE8)) lut_n2602 (.I0(x726), .I1(x727), .I2(x728), .O(n2602));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2603 (.I0(x717), .I1(x718), .I2(x719), .I3(n2599), .I4(n2600), .O(n2603));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2604 (.I0(x723), .I1(x724), .I2(x725), .I3(n2602), .I4(n2603), .O(n2604));
  LUT3 #(.INIT(8'h96)) lut_n2605 (.I0(n2589), .I1(n2592), .I2(n2593), .O(n2605));
  LUT3 #(.INIT(8'hE8)) lut_n2606 (.I0(n2601), .I1(n2604), .I2(n2605), .O(n2606));
  LUT3 #(.INIT(8'hE8)) lut_n2607 (.I0(x732), .I1(x733), .I2(x734), .O(n2607));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2608 (.I0(x723), .I1(x724), .I2(x725), .I3(n2602), .I4(n2603), .O(n2608));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2609 (.I0(x729), .I1(x730), .I2(x731), .I3(n2607), .I4(n2608), .O(n2609));
  LUT3 #(.INIT(8'hE8)) lut_n2610 (.I0(x738), .I1(x739), .I2(x740), .O(n2610));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2611 (.I0(x729), .I1(x730), .I2(x731), .I3(n2607), .I4(n2608), .O(n2611));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2612 (.I0(x735), .I1(x736), .I2(x737), .I3(n2610), .I4(n2611), .O(n2612));
  LUT3 #(.INIT(8'h96)) lut_n2613 (.I0(n2601), .I1(n2604), .I2(n2605), .O(n2613));
  LUT3 #(.INIT(8'hE8)) lut_n2614 (.I0(n2609), .I1(n2612), .I2(n2613), .O(n2614));
  LUT3 #(.INIT(8'h96)) lut_n2615 (.I0(n2586), .I1(n2594), .I2(n2595), .O(n2615));
  LUT3 #(.INIT(8'hE8)) lut_n2616 (.I0(n2606), .I1(n2614), .I2(n2615), .O(n2616));
  LUT3 #(.INIT(8'hE8)) lut_n2617 (.I0(x744), .I1(x745), .I2(x746), .O(n2617));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2618 (.I0(x735), .I1(x736), .I2(x737), .I3(n2610), .I4(n2611), .O(n2618));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2619 (.I0(x741), .I1(x742), .I2(x743), .I3(n2617), .I4(n2618), .O(n2619));
  LUT3 #(.INIT(8'hE8)) lut_n2620 (.I0(x750), .I1(x751), .I2(x752), .O(n2620));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2621 (.I0(x741), .I1(x742), .I2(x743), .I3(n2617), .I4(n2618), .O(n2621));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2622 (.I0(x747), .I1(x748), .I2(x749), .I3(n2620), .I4(n2621), .O(n2622));
  LUT3 #(.INIT(8'h96)) lut_n2623 (.I0(n2609), .I1(n2612), .I2(n2613), .O(n2623));
  LUT3 #(.INIT(8'hE8)) lut_n2624 (.I0(n2619), .I1(n2622), .I2(n2623), .O(n2624));
  LUT3 #(.INIT(8'hE8)) lut_n2625 (.I0(x756), .I1(x757), .I2(x758), .O(n2625));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2626 (.I0(x747), .I1(x748), .I2(x749), .I3(n2620), .I4(n2621), .O(n2626));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2627 (.I0(x753), .I1(x754), .I2(x755), .I3(n2625), .I4(n2626), .O(n2627));
  LUT3 #(.INIT(8'hE8)) lut_n2628 (.I0(x762), .I1(x763), .I2(x764), .O(n2628));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2629 (.I0(x753), .I1(x754), .I2(x755), .I3(n2625), .I4(n2626), .O(n2629));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2630 (.I0(x759), .I1(x760), .I2(x761), .I3(n2628), .I4(n2629), .O(n2630));
  LUT3 #(.INIT(8'h96)) lut_n2631 (.I0(n2619), .I1(n2622), .I2(n2623), .O(n2631));
  LUT3 #(.INIT(8'hE8)) lut_n2632 (.I0(n2627), .I1(n2630), .I2(n2631), .O(n2632));
  LUT3 #(.INIT(8'h96)) lut_n2633 (.I0(n2606), .I1(n2614), .I2(n2615), .O(n2633));
  LUT3 #(.INIT(8'hE8)) lut_n2634 (.I0(n2624), .I1(n2632), .I2(n2633), .O(n2634));
  LUT3 #(.INIT(8'h96)) lut_n2635 (.I0(n2578), .I1(n2596), .I2(n2597), .O(n2635));
  LUT3 #(.INIT(8'hE8)) lut_n2636 (.I0(n2616), .I1(n2634), .I2(n2635), .O(n2636));
  LUT3 #(.INIT(8'h96)) lut_n2637 (.I0(n2520), .I1(n2558), .I2(n2559), .O(n2637));
  LUT3 #(.INIT(8'hE8)) lut_n2638 (.I0(n2598), .I1(n2636), .I2(n2637), .O(n2638));
  LUT3 #(.INIT(8'h96)) lut_n2639 (.I0(n2402), .I1(n2480), .I2(n2481), .O(n2639));
  LUT3 #(.INIT(8'hE8)) lut_n2640 (.I0(n2560), .I1(n2638), .I2(n2639), .O(n2640));
  LUT3 #(.INIT(8'hE8)) lut_n2641 (.I0(n2324), .I1(n2482), .I2(n2640), .O(n2641));
  LUT3 #(.INIT(8'hE8)) lut_n2642 (.I0(x768), .I1(x769), .I2(x770), .O(n2642));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2643 (.I0(x759), .I1(x760), .I2(x761), .I3(n2628), .I4(n2629), .O(n2643));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2644 (.I0(x765), .I1(x766), .I2(x767), .I3(n2642), .I4(n2643), .O(n2644));
  LUT3 #(.INIT(8'hE8)) lut_n2645 (.I0(x774), .I1(x775), .I2(x776), .O(n2645));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2646 (.I0(x765), .I1(x766), .I2(x767), .I3(n2642), .I4(n2643), .O(n2646));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2647 (.I0(x771), .I1(x772), .I2(x773), .I3(n2645), .I4(n2646), .O(n2647));
  LUT3 #(.INIT(8'h96)) lut_n2648 (.I0(n2627), .I1(n2630), .I2(n2631), .O(n2648));
  LUT3 #(.INIT(8'hE8)) lut_n2649 (.I0(n2644), .I1(n2647), .I2(n2648), .O(n2649));
  LUT3 #(.INIT(8'hE8)) lut_n2650 (.I0(x780), .I1(x781), .I2(x782), .O(n2650));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2651 (.I0(x771), .I1(x772), .I2(x773), .I3(n2645), .I4(n2646), .O(n2651));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2652 (.I0(x777), .I1(x778), .I2(x779), .I3(n2650), .I4(n2651), .O(n2652));
  LUT3 #(.INIT(8'hE8)) lut_n2653 (.I0(x786), .I1(x787), .I2(x788), .O(n2653));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2654 (.I0(x777), .I1(x778), .I2(x779), .I3(n2650), .I4(n2651), .O(n2654));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2655 (.I0(x783), .I1(x784), .I2(x785), .I3(n2653), .I4(n2654), .O(n2655));
  LUT3 #(.INIT(8'h96)) lut_n2656 (.I0(n2644), .I1(n2647), .I2(n2648), .O(n2656));
  LUT3 #(.INIT(8'hE8)) lut_n2657 (.I0(n2652), .I1(n2655), .I2(n2656), .O(n2657));
  LUT3 #(.INIT(8'h96)) lut_n2658 (.I0(n2624), .I1(n2632), .I2(n2633), .O(n2658));
  LUT3 #(.INIT(8'hE8)) lut_n2659 (.I0(n2649), .I1(n2657), .I2(n2658), .O(n2659));
  LUT3 #(.INIT(8'hE8)) lut_n2660 (.I0(x792), .I1(x793), .I2(x794), .O(n2660));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2661 (.I0(x783), .I1(x784), .I2(x785), .I3(n2653), .I4(n2654), .O(n2661));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2662 (.I0(x789), .I1(x790), .I2(x791), .I3(n2660), .I4(n2661), .O(n2662));
  LUT3 #(.INIT(8'hE8)) lut_n2663 (.I0(x798), .I1(x799), .I2(x800), .O(n2663));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2664 (.I0(x789), .I1(x790), .I2(x791), .I3(n2660), .I4(n2661), .O(n2664));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2665 (.I0(x795), .I1(x796), .I2(x797), .I3(n2663), .I4(n2664), .O(n2665));
  LUT3 #(.INIT(8'h96)) lut_n2666 (.I0(n2652), .I1(n2655), .I2(n2656), .O(n2666));
  LUT3 #(.INIT(8'hE8)) lut_n2667 (.I0(n2662), .I1(n2665), .I2(n2666), .O(n2667));
  LUT3 #(.INIT(8'hE8)) lut_n2668 (.I0(x804), .I1(x805), .I2(x806), .O(n2668));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2669 (.I0(x795), .I1(x796), .I2(x797), .I3(n2663), .I4(n2664), .O(n2669));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2670 (.I0(x801), .I1(x802), .I2(x803), .I3(n2668), .I4(n2669), .O(n2670));
  LUT3 #(.INIT(8'hE8)) lut_n2671 (.I0(x810), .I1(x811), .I2(x812), .O(n2671));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2672 (.I0(x801), .I1(x802), .I2(x803), .I3(n2668), .I4(n2669), .O(n2672));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2673 (.I0(x807), .I1(x808), .I2(x809), .I3(n2671), .I4(n2672), .O(n2673));
  LUT3 #(.INIT(8'h96)) lut_n2674 (.I0(n2662), .I1(n2665), .I2(n2666), .O(n2674));
  LUT3 #(.INIT(8'hE8)) lut_n2675 (.I0(n2670), .I1(n2673), .I2(n2674), .O(n2675));
  LUT3 #(.INIT(8'h96)) lut_n2676 (.I0(n2649), .I1(n2657), .I2(n2658), .O(n2676));
  LUT3 #(.INIT(8'hE8)) lut_n2677 (.I0(n2667), .I1(n2675), .I2(n2676), .O(n2677));
  LUT3 #(.INIT(8'h96)) lut_n2678 (.I0(n2616), .I1(n2634), .I2(n2635), .O(n2678));
  LUT3 #(.INIT(8'hE8)) lut_n2679 (.I0(n2659), .I1(n2677), .I2(n2678), .O(n2679));
  LUT3 #(.INIT(8'hE8)) lut_n2680 (.I0(x816), .I1(x817), .I2(x818), .O(n2680));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2681 (.I0(x807), .I1(x808), .I2(x809), .I3(n2671), .I4(n2672), .O(n2681));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2682 (.I0(x813), .I1(x814), .I2(x815), .I3(n2680), .I4(n2681), .O(n2682));
  LUT3 #(.INIT(8'hE8)) lut_n2683 (.I0(x822), .I1(x823), .I2(x824), .O(n2683));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2684 (.I0(x813), .I1(x814), .I2(x815), .I3(n2680), .I4(n2681), .O(n2684));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2685 (.I0(x819), .I1(x820), .I2(x821), .I3(n2683), .I4(n2684), .O(n2685));
  LUT3 #(.INIT(8'h96)) lut_n2686 (.I0(n2670), .I1(n2673), .I2(n2674), .O(n2686));
  LUT3 #(.INIT(8'hE8)) lut_n2687 (.I0(n2682), .I1(n2685), .I2(n2686), .O(n2687));
  LUT3 #(.INIT(8'hE8)) lut_n2688 (.I0(x828), .I1(x829), .I2(x830), .O(n2688));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2689 (.I0(x819), .I1(x820), .I2(x821), .I3(n2683), .I4(n2684), .O(n2689));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2690 (.I0(x825), .I1(x826), .I2(x827), .I3(n2688), .I4(n2689), .O(n2690));
  LUT3 #(.INIT(8'hE8)) lut_n2691 (.I0(x834), .I1(x835), .I2(x836), .O(n2691));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2692 (.I0(x825), .I1(x826), .I2(x827), .I3(n2688), .I4(n2689), .O(n2692));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2693 (.I0(x831), .I1(x832), .I2(x833), .I3(n2691), .I4(n2692), .O(n2693));
  LUT3 #(.INIT(8'h96)) lut_n2694 (.I0(n2682), .I1(n2685), .I2(n2686), .O(n2694));
  LUT3 #(.INIT(8'hE8)) lut_n2695 (.I0(n2690), .I1(n2693), .I2(n2694), .O(n2695));
  LUT3 #(.INIT(8'h96)) lut_n2696 (.I0(n2667), .I1(n2675), .I2(n2676), .O(n2696));
  LUT3 #(.INIT(8'hE8)) lut_n2697 (.I0(n2687), .I1(n2695), .I2(n2696), .O(n2697));
  LUT3 #(.INIT(8'hE8)) lut_n2698 (.I0(x840), .I1(x841), .I2(x842), .O(n2698));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2699 (.I0(x831), .I1(x832), .I2(x833), .I3(n2691), .I4(n2692), .O(n2699));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2700 (.I0(x837), .I1(x838), .I2(x839), .I3(n2698), .I4(n2699), .O(n2700));
  LUT3 #(.INIT(8'hE8)) lut_n2701 (.I0(x846), .I1(x847), .I2(x848), .O(n2701));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2702 (.I0(x837), .I1(x838), .I2(x839), .I3(n2698), .I4(n2699), .O(n2702));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2703 (.I0(x843), .I1(x844), .I2(x845), .I3(n2701), .I4(n2702), .O(n2703));
  LUT3 #(.INIT(8'h96)) lut_n2704 (.I0(n2690), .I1(n2693), .I2(n2694), .O(n2704));
  LUT3 #(.INIT(8'hE8)) lut_n2705 (.I0(n2700), .I1(n2703), .I2(n2704), .O(n2705));
  LUT3 #(.INIT(8'hE8)) lut_n2706 (.I0(x852), .I1(x853), .I2(x854), .O(n2706));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2707 (.I0(x843), .I1(x844), .I2(x845), .I3(n2701), .I4(n2702), .O(n2707));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2708 (.I0(x849), .I1(x850), .I2(x851), .I3(n2706), .I4(n2707), .O(n2708));
  LUT3 #(.INIT(8'hE8)) lut_n2709 (.I0(x858), .I1(x859), .I2(x860), .O(n2709));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2710 (.I0(x849), .I1(x850), .I2(x851), .I3(n2706), .I4(n2707), .O(n2710));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2711 (.I0(x855), .I1(x856), .I2(x857), .I3(n2709), .I4(n2710), .O(n2711));
  LUT3 #(.INIT(8'h96)) lut_n2712 (.I0(n2700), .I1(n2703), .I2(n2704), .O(n2712));
  LUT3 #(.INIT(8'hE8)) lut_n2713 (.I0(n2708), .I1(n2711), .I2(n2712), .O(n2713));
  LUT3 #(.INIT(8'h96)) lut_n2714 (.I0(n2687), .I1(n2695), .I2(n2696), .O(n2714));
  LUT3 #(.INIT(8'hE8)) lut_n2715 (.I0(n2705), .I1(n2713), .I2(n2714), .O(n2715));
  LUT3 #(.INIT(8'h96)) lut_n2716 (.I0(n2659), .I1(n2677), .I2(n2678), .O(n2716));
  LUT3 #(.INIT(8'hE8)) lut_n2717 (.I0(n2697), .I1(n2715), .I2(n2716), .O(n2717));
  LUT3 #(.INIT(8'h96)) lut_n2718 (.I0(n2598), .I1(n2636), .I2(n2637), .O(n2718));
  LUT3 #(.INIT(8'hE8)) lut_n2719 (.I0(n2679), .I1(n2717), .I2(n2718), .O(n2719));
  LUT3 #(.INIT(8'hE8)) lut_n2720 (.I0(x864), .I1(x865), .I2(x866), .O(n2720));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2721 (.I0(x855), .I1(x856), .I2(x857), .I3(n2709), .I4(n2710), .O(n2721));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2722 (.I0(x861), .I1(x862), .I2(x863), .I3(n2720), .I4(n2721), .O(n2722));
  LUT3 #(.INIT(8'hE8)) lut_n2723 (.I0(x870), .I1(x871), .I2(x872), .O(n2723));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2724 (.I0(x861), .I1(x862), .I2(x863), .I3(n2720), .I4(n2721), .O(n2724));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2725 (.I0(x867), .I1(x868), .I2(x869), .I3(n2723), .I4(n2724), .O(n2725));
  LUT3 #(.INIT(8'h96)) lut_n2726 (.I0(n2708), .I1(n2711), .I2(n2712), .O(n2726));
  LUT3 #(.INIT(8'hE8)) lut_n2727 (.I0(n2722), .I1(n2725), .I2(n2726), .O(n2727));
  LUT3 #(.INIT(8'hE8)) lut_n2728 (.I0(x876), .I1(x877), .I2(x878), .O(n2728));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2729 (.I0(x867), .I1(x868), .I2(x869), .I3(n2723), .I4(n2724), .O(n2729));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2730 (.I0(x873), .I1(x874), .I2(x875), .I3(n2728), .I4(n2729), .O(n2730));
  LUT3 #(.INIT(8'hE8)) lut_n2731 (.I0(x882), .I1(x883), .I2(x884), .O(n2731));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2732 (.I0(x873), .I1(x874), .I2(x875), .I3(n2728), .I4(n2729), .O(n2732));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2733 (.I0(x879), .I1(x880), .I2(x881), .I3(n2731), .I4(n2732), .O(n2733));
  LUT3 #(.INIT(8'h96)) lut_n2734 (.I0(n2722), .I1(n2725), .I2(n2726), .O(n2734));
  LUT3 #(.INIT(8'hE8)) lut_n2735 (.I0(n2730), .I1(n2733), .I2(n2734), .O(n2735));
  LUT3 #(.INIT(8'h96)) lut_n2736 (.I0(n2705), .I1(n2713), .I2(n2714), .O(n2736));
  LUT3 #(.INIT(8'hE8)) lut_n2737 (.I0(n2727), .I1(n2735), .I2(n2736), .O(n2737));
  LUT3 #(.INIT(8'hE8)) lut_n2738 (.I0(x888), .I1(x889), .I2(x890), .O(n2738));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2739 (.I0(x879), .I1(x880), .I2(x881), .I3(n2731), .I4(n2732), .O(n2739));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2740 (.I0(x885), .I1(x886), .I2(x887), .I3(n2738), .I4(n2739), .O(n2740));
  LUT3 #(.INIT(8'hE8)) lut_n2741 (.I0(x894), .I1(x895), .I2(x896), .O(n2741));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2742 (.I0(x885), .I1(x886), .I2(x887), .I3(n2738), .I4(n2739), .O(n2742));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2743 (.I0(x891), .I1(x892), .I2(x893), .I3(n2741), .I4(n2742), .O(n2743));
  LUT3 #(.INIT(8'h96)) lut_n2744 (.I0(n2730), .I1(n2733), .I2(n2734), .O(n2744));
  LUT3 #(.INIT(8'hE8)) lut_n2745 (.I0(n2740), .I1(n2743), .I2(n2744), .O(n2745));
  LUT3 #(.INIT(8'hE8)) lut_n2746 (.I0(x900), .I1(x901), .I2(x902), .O(n2746));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2747 (.I0(x891), .I1(x892), .I2(x893), .I3(n2741), .I4(n2742), .O(n2747));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2748 (.I0(x897), .I1(x898), .I2(x899), .I3(n2746), .I4(n2747), .O(n2748));
  LUT3 #(.INIT(8'hE8)) lut_n2749 (.I0(x906), .I1(x907), .I2(x908), .O(n2749));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2750 (.I0(x897), .I1(x898), .I2(x899), .I3(n2746), .I4(n2747), .O(n2750));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2751 (.I0(x903), .I1(x904), .I2(x905), .I3(n2749), .I4(n2750), .O(n2751));
  LUT3 #(.INIT(8'h96)) lut_n2752 (.I0(n2740), .I1(n2743), .I2(n2744), .O(n2752));
  LUT3 #(.INIT(8'hE8)) lut_n2753 (.I0(n2748), .I1(n2751), .I2(n2752), .O(n2753));
  LUT3 #(.INIT(8'h96)) lut_n2754 (.I0(n2727), .I1(n2735), .I2(n2736), .O(n2754));
  LUT3 #(.INIT(8'hE8)) lut_n2755 (.I0(n2745), .I1(n2753), .I2(n2754), .O(n2755));
  LUT3 #(.INIT(8'h96)) lut_n2756 (.I0(n2697), .I1(n2715), .I2(n2716), .O(n2756));
  LUT3 #(.INIT(8'hE8)) lut_n2757 (.I0(n2737), .I1(n2755), .I2(n2756), .O(n2757));
  LUT3 #(.INIT(8'hE8)) lut_n2758 (.I0(x912), .I1(x913), .I2(x914), .O(n2758));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2759 (.I0(x903), .I1(x904), .I2(x905), .I3(n2749), .I4(n2750), .O(n2759));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2760 (.I0(x909), .I1(x910), .I2(x911), .I3(n2758), .I4(n2759), .O(n2760));
  LUT3 #(.INIT(8'hE8)) lut_n2761 (.I0(x918), .I1(x919), .I2(x920), .O(n2761));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2762 (.I0(x909), .I1(x910), .I2(x911), .I3(n2758), .I4(n2759), .O(n2762));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2763 (.I0(x915), .I1(x916), .I2(x917), .I3(n2761), .I4(n2762), .O(n2763));
  LUT3 #(.INIT(8'h96)) lut_n2764 (.I0(n2748), .I1(n2751), .I2(n2752), .O(n2764));
  LUT3 #(.INIT(8'hE8)) lut_n2765 (.I0(n2760), .I1(n2763), .I2(n2764), .O(n2765));
  LUT3 #(.INIT(8'hE8)) lut_n2766 (.I0(x924), .I1(x925), .I2(x926), .O(n2766));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2767 (.I0(x915), .I1(x916), .I2(x917), .I3(n2761), .I4(n2762), .O(n2767));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2768 (.I0(x921), .I1(x922), .I2(x923), .I3(n2766), .I4(n2767), .O(n2768));
  LUT3 #(.INIT(8'hE8)) lut_n2769 (.I0(x930), .I1(x931), .I2(x932), .O(n2769));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2770 (.I0(x921), .I1(x922), .I2(x923), .I3(n2766), .I4(n2767), .O(n2770));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2771 (.I0(x927), .I1(x928), .I2(x929), .I3(n2769), .I4(n2770), .O(n2771));
  LUT3 #(.INIT(8'h96)) lut_n2772 (.I0(n2760), .I1(n2763), .I2(n2764), .O(n2772));
  LUT3 #(.INIT(8'hE8)) lut_n2773 (.I0(n2768), .I1(n2771), .I2(n2772), .O(n2773));
  LUT3 #(.INIT(8'h96)) lut_n2774 (.I0(n2745), .I1(n2753), .I2(n2754), .O(n2774));
  LUT3 #(.INIT(8'hE8)) lut_n2775 (.I0(n2765), .I1(n2773), .I2(n2774), .O(n2775));
  LUT3 #(.INIT(8'hE8)) lut_n2776 (.I0(x936), .I1(x937), .I2(x938), .O(n2776));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2777 (.I0(x927), .I1(x928), .I2(x929), .I3(n2769), .I4(n2770), .O(n2777));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2778 (.I0(x933), .I1(x934), .I2(x935), .I3(n2776), .I4(n2777), .O(n2778));
  LUT3 #(.INIT(8'hE8)) lut_n2779 (.I0(x942), .I1(x943), .I2(x944), .O(n2779));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2780 (.I0(x933), .I1(x934), .I2(x935), .I3(n2776), .I4(n2777), .O(n2780));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2781 (.I0(x939), .I1(x940), .I2(x941), .I3(n2779), .I4(n2780), .O(n2781));
  LUT3 #(.INIT(8'h96)) lut_n2782 (.I0(n2768), .I1(n2771), .I2(n2772), .O(n2782));
  LUT3 #(.INIT(8'hE8)) lut_n2783 (.I0(n2778), .I1(n2781), .I2(n2782), .O(n2783));
  LUT3 #(.INIT(8'hE8)) lut_n2784 (.I0(x948), .I1(x949), .I2(x950), .O(n2784));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2785 (.I0(x939), .I1(x940), .I2(x941), .I3(n2779), .I4(n2780), .O(n2785));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2786 (.I0(x945), .I1(x946), .I2(x947), .I3(n2784), .I4(n2785), .O(n2786));
  LUT3 #(.INIT(8'hE8)) lut_n2787 (.I0(x954), .I1(x955), .I2(x956), .O(n2787));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2788 (.I0(x945), .I1(x946), .I2(x947), .I3(n2784), .I4(n2785), .O(n2788));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2789 (.I0(x951), .I1(x952), .I2(x953), .I3(n2787), .I4(n2788), .O(n2789));
  LUT3 #(.INIT(8'h96)) lut_n2790 (.I0(n2778), .I1(n2781), .I2(n2782), .O(n2790));
  LUT3 #(.INIT(8'hE8)) lut_n2791 (.I0(n2786), .I1(n2789), .I2(n2790), .O(n2791));
  LUT3 #(.INIT(8'h96)) lut_n2792 (.I0(n2765), .I1(n2773), .I2(n2774), .O(n2792));
  LUT3 #(.INIT(8'hE8)) lut_n2793 (.I0(n2783), .I1(n2791), .I2(n2792), .O(n2793));
  LUT3 #(.INIT(8'h96)) lut_n2794 (.I0(n2737), .I1(n2755), .I2(n2756), .O(n2794));
  LUT3 #(.INIT(8'hE8)) lut_n2795 (.I0(n2775), .I1(n2793), .I2(n2794), .O(n2795));
  LUT3 #(.INIT(8'h96)) lut_n2796 (.I0(n2679), .I1(n2717), .I2(n2718), .O(n2796));
  LUT3 #(.INIT(8'hE8)) lut_n2797 (.I0(n2757), .I1(n2795), .I2(n2796), .O(n2797));
  LUT3 #(.INIT(8'h96)) lut_n2798 (.I0(n2560), .I1(n2638), .I2(n2639), .O(n2798));
  LUT3 #(.INIT(8'hE8)) lut_n2799 (.I0(n2719), .I1(n2797), .I2(n2798), .O(n2799));
  LUT3 #(.INIT(8'hE8)) lut_n2800 (.I0(x960), .I1(x961), .I2(x962), .O(n2800));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2801 (.I0(x951), .I1(x952), .I2(x953), .I3(n2787), .I4(n2788), .O(n2801));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2802 (.I0(x957), .I1(x958), .I2(x959), .I3(n2800), .I4(n2801), .O(n2802));
  LUT3 #(.INIT(8'hE8)) lut_n2803 (.I0(x966), .I1(x967), .I2(x968), .O(n2803));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2804 (.I0(x957), .I1(x958), .I2(x959), .I3(n2800), .I4(n2801), .O(n2804));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2805 (.I0(x963), .I1(x964), .I2(x965), .I3(n2803), .I4(n2804), .O(n2805));
  LUT3 #(.INIT(8'h96)) lut_n2806 (.I0(n2786), .I1(n2789), .I2(n2790), .O(n2806));
  LUT3 #(.INIT(8'hE8)) lut_n2807 (.I0(n2802), .I1(n2805), .I2(n2806), .O(n2807));
  LUT3 #(.INIT(8'hE8)) lut_n2808 (.I0(x972), .I1(x973), .I2(x974), .O(n2808));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2809 (.I0(x963), .I1(x964), .I2(x965), .I3(n2803), .I4(n2804), .O(n2809));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2810 (.I0(x969), .I1(x970), .I2(x971), .I3(n2808), .I4(n2809), .O(n2810));
  LUT3 #(.INIT(8'hE8)) lut_n2811 (.I0(x978), .I1(x979), .I2(x980), .O(n2811));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2812 (.I0(x969), .I1(x970), .I2(x971), .I3(n2808), .I4(n2809), .O(n2812));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2813 (.I0(x975), .I1(x976), .I2(x977), .I3(n2811), .I4(n2812), .O(n2813));
  LUT3 #(.INIT(8'h96)) lut_n2814 (.I0(n2802), .I1(n2805), .I2(n2806), .O(n2814));
  LUT3 #(.INIT(8'hE8)) lut_n2815 (.I0(n2810), .I1(n2813), .I2(n2814), .O(n2815));
  LUT3 #(.INIT(8'h96)) lut_n2816 (.I0(n2783), .I1(n2791), .I2(n2792), .O(n2816));
  LUT3 #(.INIT(8'hE8)) lut_n2817 (.I0(n2807), .I1(n2815), .I2(n2816), .O(n2817));
  LUT3 #(.INIT(8'hE8)) lut_n2818 (.I0(x984), .I1(x985), .I2(x986), .O(n2818));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2819 (.I0(x975), .I1(x976), .I2(x977), .I3(n2811), .I4(n2812), .O(n2819));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2820 (.I0(x981), .I1(x982), .I2(x983), .I3(n2818), .I4(n2819), .O(n2820));
  LUT3 #(.INIT(8'hE8)) lut_n2821 (.I0(x990), .I1(x991), .I2(x992), .O(n2821));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2822 (.I0(x981), .I1(x982), .I2(x983), .I3(n2818), .I4(n2819), .O(n2822));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2823 (.I0(x987), .I1(x988), .I2(x989), .I3(n2821), .I4(n2822), .O(n2823));
  LUT3 #(.INIT(8'h96)) lut_n2824 (.I0(n2810), .I1(n2813), .I2(n2814), .O(n2824));
  LUT3 #(.INIT(8'hE8)) lut_n2825 (.I0(n2820), .I1(n2823), .I2(n2824), .O(n2825));
  LUT3 #(.INIT(8'hE8)) lut_n2826 (.I0(x996), .I1(x997), .I2(x998), .O(n2826));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2827 (.I0(x987), .I1(x988), .I2(x989), .I3(n2821), .I4(n2822), .O(n2827));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2828 (.I0(x993), .I1(x994), .I2(x995), .I3(n2826), .I4(n2827), .O(n2828));
  LUT3 #(.INIT(8'hE8)) lut_n2829 (.I0(x1002), .I1(x1003), .I2(x1004), .O(n2829));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2830 (.I0(x993), .I1(x994), .I2(x995), .I3(n2826), .I4(n2827), .O(n2830));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2831 (.I0(x999), .I1(x1000), .I2(x1001), .I3(n2829), .I4(n2830), .O(n2831));
  LUT3 #(.INIT(8'h96)) lut_n2832 (.I0(n2820), .I1(n2823), .I2(n2824), .O(n2832));
  LUT3 #(.INIT(8'hE8)) lut_n2833 (.I0(n2828), .I1(n2831), .I2(n2832), .O(n2833));
  LUT3 #(.INIT(8'h96)) lut_n2834 (.I0(n2807), .I1(n2815), .I2(n2816), .O(n2834));
  LUT3 #(.INIT(8'hE8)) lut_n2835 (.I0(n2825), .I1(n2833), .I2(n2834), .O(n2835));
  LUT3 #(.INIT(8'h96)) lut_n2836 (.I0(n2775), .I1(n2793), .I2(n2794), .O(n2836));
  LUT3 #(.INIT(8'hE8)) lut_n2837 (.I0(n2817), .I1(n2835), .I2(n2836), .O(n2837));
  LUT3 #(.INIT(8'hE8)) lut_n2838 (.I0(x1008), .I1(x1009), .I2(x1010), .O(n2838));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2839 (.I0(x999), .I1(x1000), .I2(x1001), .I3(n2829), .I4(n2830), .O(n2839));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2840 (.I0(x1005), .I1(x1006), .I2(x1007), .I3(n2838), .I4(n2839), .O(n2840));
  LUT3 #(.INIT(8'hE8)) lut_n2841 (.I0(x1014), .I1(x1015), .I2(x1016), .O(n2841));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2842 (.I0(x1005), .I1(x1006), .I2(x1007), .I3(n2838), .I4(n2839), .O(n2842));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2843 (.I0(x1011), .I1(x1012), .I2(x1013), .I3(n2841), .I4(n2842), .O(n2843));
  LUT3 #(.INIT(8'h96)) lut_n2844 (.I0(n2828), .I1(n2831), .I2(n2832), .O(n2844));
  LUT3 #(.INIT(8'hE8)) lut_n2845 (.I0(n2840), .I1(n2843), .I2(n2844), .O(n2845));
  LUT3 #(.INIT(8'hE8)) lut_n2846 (.I0(x1020), .I1(x1021), .I2(x1022), .O(n2846));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2847 (.I0(x1011), .I1(x1012), .I2(x1013), .I3(n2841), .I4(n2842), .O(n2847));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2848 (.I0(x1017), .I1(x1018), .I2(x1019), .I3(n2846), .I4(n2847), .O(n2848));
  LUT3 #(.INIT(8'hE8)) lut_n2849 (.I0(x1026), .I1(x1027), .I2(x1028), .O(n2849));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2850 (.I0(x1017), .I1(x1018), .I2(x1019), .I3(n2846), .I4(n2847), .O(n2850));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2851 (.I0(x1023), .I1(x1024), .I2(x1025), .I3(n2849), .I4(n2850), .O(n2851));
  LUT3 #(.INIT(8'h96)) lut_n2852 (.I0(n2840), .I1(n2843), .I2(n2844), .O(n2852));
  LUT3 #(.INIT(8'hE8)) lut_n2853 (.I0(n2848), .I1(n2851), .I2(n2852), .O(n2853));
  LUT3 #(.INIT(8'h96)) lut_n2854 (.I0(n2825), .I1(n2833), .I2(n2834), .O(n2854));
  LUT3 #(.INIT(8'hE8)) lut_n2855 (.I0(n2845), .I1(n2853), .I2(n2854), .O(n2855));
  LUT3 #(.INIT(8'hE8)) lut_n2856 (.I0(x1032), .I1(x1033), .I2(x1034), .O(n2856));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2857 (.I0(x1023), .I1(x1024), .I2(x1025), .I3(n2849), .I4(n2850), .O(n2857));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2858 (.I0(x1029), .I1(x1030), .I2(x1031), .I3(n2856), .I4(n2857), .O(n2858));
  LUT3 #(.INIT(8'hE8)) lut_n2859 (.I0(x1038), .I1(x1039), .I2(x1040), .O(n2859));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2860 (.I0(x1029), .I1(x1030), .I2(x1031), .I3(n2856), .I4(n2857), .O(n2860));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2861 (.I0(x1035), .I1(x1036), .I2(x1037), .I3(n2859), .I4(n2860), .O(n2861));
  LUT3 #(.INIT(8'h96)) lut_n2862 (.I0(n2848), .I1(n2851), .I2(n2852), .O(n2862));
  LUT3 #(.INIT(8'hE8)) lut_n2863 (.I0(n2858), .I1(n2861), .I2(n2862), .O(n2863));
  LUT3 #(.INIT(8'hE8)) lut_n2864 (.I0(x1044), .I1(x1045), .I2(x1046), .O(n2864));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2865 (.I0(x1035), .I1(x1036), .I2(x1037), .I3(n2859), .I4(n2860), .O(n2865));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2866 (.I0(x1041), .I1(x1042), .I2(x1043), .I3(n2864), .I4(n2865), .O(n2866));
  LUT3 #(.INIT(8'hE8)) lut_n2867 (.I0(x1050), .I1(x1051), .I2(x1052), .O(n2867));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2868 (.I0(x1041), .I1(x1042), .I2(x1043), .I3(n2864), .I4(n2865), .O(n2868));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2869 (.I0(x1047), .I1(x1048), .I2(x1049), .I3(n2867), .I4(n2868), .O(n2869));
  LUT3 #(.INIT(8'h96)) lut_n2870 (.I0(n2858), .I1(n2861), .I2(n2862), .O(n2870));
  LUT3 #(.INIT(8'hE8)) lut_n2871 (.I0(n2866), .I1(n2869), .I2(n2870), .O(n2871));
  LUT3 #(.INIT(8'h96)) lut_n2872 (.I0(n2845), .I1(n2853), .I2(n2854), .O(n2872));
  LUT3 #(.INIT(8'hE8)) lut_n2873 (.I0(n2863), .I1(n2871), .I2(n2872), .O(n2873));
  LUT3 #(.INIT(8'h96)) lut_n2874 (.I0(n2817), .I1(n2835), .I2(n2836), .O(n2874));
  LUT3 #(.INIT(8'hE8)) lut_n2875 (.I0(n2855), .I1(n2873), .I2(n2874), .O(n2875));
  LUT3 #(.INIT(8'h96)) lut_n2876 (.I0(n2757), .I1(n2795), .I2(n2796), .O(n2876));
  LUT3 #(.INIT(8'hE8)) lut_n2877 (.I0(n2837), .I1(n2875), .I2(n2876), .O(n2877));
  LUT3 #(.INIT(8'hE8)) lut_n2878 (.I0(x1056), .I1(x1057), .I2(x1058), .O(n2878));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2879 (.I0(x1047), .I1(x1048), .I2(x1049), .I3(n2867), .I4(n2868), .O(n2879));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2880 (.I0(x1053), .I1(x1054), .I2(x1055), .I3(n2878), .I4(n2879), .O(n2880));
  LUT3 #(.INIT(8'hE8)) lut_n2881 (.I0(x1062), .I1(x1063), .I2(x1064), .O(n2881));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2882 (.I0(x1053), .I1(x1054), .I2(x1055), .I3(n2878), .I4(n2879), .O(n2882));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2883 (.I0(x1059), .I1(x1060), .I2(x1061), .I3(n2881), .I4(n2882), .O(n2883));
  LUT3 #(.INIT(8'h96)) lut_n2884 (.I0(n2866), .I1(n2869), .I2(n2870), .O(n2884));
  LUT3 #(.INIT(8'hE8)) lut_n2885 (.I0(n2880), .I1(n2883), .I2(n2884), .O(n2885));
  LUT3 #(.INIT(8'hE8)) lut_n2886 (.I0(x1068), .I1(x1069), .I2(x1070), .O(n2886));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2887 (.I0(x1059), .I1(x1060), .I2(x1061), .I3(n2881), .I4(n2882), .O(n2887));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2888 (.I0(x1065), .I1(x1066), .I2(x1067), .I3(n2886), .I4(n2887), .O(n2888));
  LUT3 #(.INIT(8'hE8)) lut_n2889 (.I0(x1074), .I1(x1075), .I2(x1076), .O(n2889));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2890 (.I0(x1065), .I1(x1066), .I2(x1067), .I3(n2886), .I4(n2887), .O(n2890));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2891 (.I0(x1071), .I1(x1072), .I2(x1073), .I3(n2889), .I4(n2890), .O(n2891));
  LUT3 #(.INIT(8'h96)) lut_n2892 (.I0(n2880), .I1(n2883), .I2(n2884), .O(n2892));
  LUT3 #(.INIT(8'hE8)) lut_n2893 (.I0(n2888), .I1(n2891), .I2(n2892), .O(n2893));
  LUT3 #(.INIT(8'h96)) lut_n2894 (.I0(n2863), .I1(n2871), .I2(n2872), .O(n2894));
  LUT3 #(.INIT(8'hE8)) lut_n2895 (.I0(n2885), .I1(n2893), .I2(n2894), .O(n2895));
  LUT3 #(.INIT(8'hE8)) lut_n2896 (.I0(x1080), .I1(x1081), .I2(x1082), .O(n2896));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2897 (.I0(x1071), .I1(x1072), .I2(x1073), .I3(n2889), .I4(n2890), .O(n2897));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2898 (.I0(x1077), .I1(x1078), .I2(x1079), .I3(n2896), .I4(n2897), .O(n2898));
  LUT3 #(.INIT(8'hE8)) lut_n2899 (.I0(x1086), .I1(x1087), .I2(x1088), .O(n2899));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2900 (.I0(x1077), .I1(x1078), .I2(x1079), .I3(n2896), .I4(n2897), .O(n2900));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2901 (.I0(x1083), .I1(x1084), .I2(x1085), .I3(n2899), .I4(n2900), .O(n2901));
  LUT3 #(.INIT(8'h96)) lut_n2902 (.I0(n2888), .I1(n2891), .I2(n2892), .O(n2902));
  LUT3 #(.INIT(8'hE8)) lut_n2903 (.I0(n2898), .I1(n2901), .I2(n2902), .O(n2903));
  LUT3 #(.INIT(8'hE8)) lut_n2904 (.I0(x1092), .I1(x1093), .I2(x1094), .O(n2904));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2905 (.I0(x1083), .I1(x1084), .I2(x1085), .I3(n2899), .I4(n2900), .O(n2905));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2906 (.I0(x1089), .I1(x1090), .I2(x1091), .I3(n2904), .I4(n2905), .O(n2906));
  LUT3 #(.INIT(8'hE8)) lut_n2907 (.I0(x1098), .I1(x1099), .I2(x1100), .O(n2907));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2908 (.I0(x1089), .I1(x1090), .I2(x1091), .I3(n2904), .I4(n2905), .O(n2908));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2909 (.I0(x1095), .I1(x1096), .I2(x1097), .I3(n2907), .I4(n2908), .O(n2909));
  LUT3 #(.INIT(8'h96)) lut_n2910 (.I0(n2898), .I1(n2901), .I2(n2902), .O(n2910));
  LUT3 #(.INIT(8'hE8)) lut_n2911 (.I0(n2906), .I1(n2909), .I2(n2910), .O(n2911));
  LUT3 #(.INIT(8'h96)) lut_n2912 (.I0(n2885), .I1(n2893), .I2(n2894), .O(n2912));
  LUT3 #(.INIT(8'hE8)) lut_n2913 (.I0(n2903), .I1(n2911), .I2(n2912), .O(n2913));
  LUT3 #(.INIT(8'h96)) lut_n2914 (.I0(n2855), .I1(n2873), .I2(n2874), .O(n2914));
  LUT3 #(.INIT(8'hE8)) lut_n2915 (.I0(n2895), .I1(n2913), .I2(n2914), .O(n2915));
  LUT3 #(.INIT(8'hE8)) lut_n2916 (.I0(x1104), .I1(x1105), .I2(x1106), .O(n2916));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2917 (.I0(x1095), .I1(x1096), .I2(x1097), .I3(n2907), .I4(n2908), .O(n2917));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2918 (.I0(x1101), .I1(x1102), .I2(x1103), .I3(n2916), .I4(n2917), .O(n2918));
  LUT3 #(.INIT(8'hE8)) lut_n2919 (.I0(x1110), .I1(x1111), .I2(x1112), .O(n2919));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2920 (.I0(x1101), .I1(x1102), .I2(x1103), .I3(n2916), .I4(n2917), .O(n2920));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2921 (.I0(x1107), .I1(x1108), .I2(x1109), .I3(n2919), .I4(n2920), .O(n2921));
  LUT3 #(.INIT(8'h96)) lut_n2922 (.I0(n2906), .I1(n2909), .I2(n2910), .O(n2922));
  LUT3 #(.INIT(8'hE8)) lut_n2923 (.I0(n2918), .I1(n2921), .I2(n2922), .O(n2923));
  LUT3 #(.INIT(8'hE8)) lut_n2924 (.I0(x1116), .I1(x1117), .I2(x1118), .O(n2924));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2925 (.I0(x1107), .I1(x1108), .I2(x1109), .I3(n2919), .I4(n2920), .O(n2925));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2926 (.I0(x1113), .I1(x1114), .I2(x1115), .I3(n2924), .I4(n2925), .O(n2926));
  LUT3 #(.INIT(8'hE8)) lut_n2927 (.I0(x1122), .I1(x1123), .I2(x1124), .O(n2927));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2928 (.I0(x1113), .I1(x1114), .I2(x1115), .I3(n2924), .I4(n2925), .O(n2928));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2929 (.I0(x1119), .I1(x1120), .I2(x1121), .I3(n2927), .I4(n2928), .O(n2929));
  LUT3 #(.INIT(8'h96)) lut_n2930 (.I0(n2918), .I1(n2921), .I2(n2922), .O(n2930));
  LUT3 #(.INIT(8'hE8)) lut_n2931 (.I0(n2926), .I1(n2929), .I2(n2930), .O(n2931));
  LUT3 #(.INIT(8'h96)) lut_n2932 (.I0(n2903), .I1(n2911), .I2(n2912), .O(n2932));
  LUT3 #(.INIT(8'hE8)) lut_n2933 (.I0(n2923), .I1(n2931), .I2(n2932), .O(n2933));
  LUT3 #(.INIT(8'hE8)) lut_n2934 (.I0(x1128), .I1(x1129), .I2(x1130), .O(n2934));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2935 (.I0(x1119), .I1(x1120), .I2(x1121), .I3(n2927), .I4(n2928), .O(n2935));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2936 (.I0(x1125), .I1(x1126), .I2(x1127), .I3(n2934), .I4(n2935), .O(n2936));
  LUT3 #(.INIT(8'hE8)) lut_n2937 (.I0(x1134), .I1(x1135), .I2(x1136), .O(n2937));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2938 (.I0(x1125), .I1(x1126), .I2(x1127), .I3(n2934), .I4(n2935), .O(n2938));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2939 (.I0(x1131), .I1(x1132), .I2(x1133), .I3(n2937), .I4(n2938), .O(n2939));
  LUT3 #(.INIT(8'h96)) lut_n2940 (.I0(n2926), .I1(n2929), .I2(n2930), .O(n2940));
  LUT3 #(.INIT(8'hE8)) lut_n2941 (.I0(n2936), .I1(n2939), .I2(n2940), .O(n2941));
  LUT3 #(.INIT(8'hE8)) lut_n2942 (.I0(x1140), .I1(x1141), .I2(x1142), .O(n2942));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2943 (.I0(x1131), .I1(x1132), .I2(x1133), .I3(n2937), .I4(n2938), .O(n2943));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2944 (.I0(x1137), .I1(x1138), .I2(x1139), .I3(n2942), .I4(n2943), .O(n2944));
  LUT3 #(.INIT(8'hE8)) lut_n2945 (.I0(x1146), .I1(x1147), .I2(x1148), .O(n2945));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2946 (.I0(x1137), .I1(x1138), .I2(x1139), .I3(n2942), .I4(n2943), .O(n2946));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2947 (.I0(x1143), .I1(x1144), .I2(x1145), .I3(n2945), .I4(n2946), .O(n2947));
  LUT3 #(.INIT(8'h96)) lut_n2948 (.I0(n2936), .I1(n2939), .I2(n2940), .O(n2948));
  LUT3 #(.INIT(8'hE8)) lut_n2949 (.I0(n2944), .I1(n2947), .I2(n2948), .O(n2949));
  LUT3 #(.INIT(8'h96)) lut_n2950 (.I0(n2923), .I1(n2931), .I2(n2932), .O(n2950));
  LUT3 #(.INIT(8'hE8)) lut_n2951 (.I0(n2941), .I1(n2949), .I2(n2950), .O(n2951));
  LUT3 #(.INIT(8'h96)) lut_n2952 (.I0(n2895), .I1(n2913), .I2(n2914), .O(n2952));
  LUT3 #(.INIT(8'hE8)) lut_n2953 (.I0(n2933), .I1(n2951), .I2(n2952), .O(n2953));
  LUT3 #(.INIT(8'h96)) lut_n2954 (.I0(n2837), .I1(n2875), .I2(n2876), .O(n2954));
  LUT3 #(.INIT(8'hE8)) lut_n2955 (.I0(n2915), .I1(n2953), .I2(n2954), .O(n2955));
  LUT3 #(.INIT(8'h96)) lut_n2956 (.I0(n2719), .I1(n2797), .I2(n2798), .O(n2956));
  LUT3 #(.INIT(8'hE8)) lut_n2957 (.I0(n2877), .I1(n2955), .I2(n2956), .O(n2957));
  LUT3 #(.INIT(8'h96)) lut_n2958 (.I0(n2324), .I1(n2482), .I2(n2640), .O(n2958));
  LUT3 #(.INIT(8'hE8)) lut_n2959 (.I0(n2799), .I1(n2957), .I2(n2958), .O(n2959));
  LUT3 #(.INIT(8'hE8)) lut_n2960 (.I0(x1152), .I1(x1153), .I2(x1154), .O(n2960));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2961 (.I0(x1143), .I1(x1144), .I2(x1145), .I3(n2945), .I4(n2946), .O(n2961));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2962 (.I0(x1149), .I1(x1150), .I2(x1151), .I3(n2960), .I4(n2961), .O(n2962));
  LUT3 #(.INIT(8'hE8)) lut_n2963 (.I0(x1158), .I1(x1159), .I2(x1160), .O(n2963));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2964 (.I0(x1149), .I1(x1150), .I2(x1151), .I3(n2960), .I4(n2961), .O(n2964));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2965 (.I0(x1155), .I1(x1156), .I2(x1157), .I3(n2963), .I4(n2964), .O(n2965));
  LUT3 #(.INIT(8'h96)) lut_n2966 (.I0(n2944), .I1(n2947), .I2(n2948), .O(n2966));
  LUT3 #(.INIT(8'hE8)) lut_n2967 (.I0(n2962), .I1(n2965), .I2(n2966), .O(n2967));
  LUT3 #(.INIT(8'hE8)) lut_n2968 (.I0(x1164), .I1(x1165), .I2(x1166), .O(n2968));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2969 (.I0(x1155), .I1(x1156), .I2(x1157), .I3(n2963), .I4(n2964), .O(n2969));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2970 (.I0(x1161), .I1(x1162), .I2(x1163), .I3(n2968), .I4(n2969), .O(n2970));
  LUT3 #(.INIT(8'hE8)) lut_n2971 (.I0(x1170), .I1(x1171), .I2(x1172), .O(n2971));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2972 (.I0(x1161), .I1(x1162), .I2(x1163), .I3(n2968), .I4(n2969), .O(n2972));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2973 (.I0(x1167), .I1(x1168), .I2(x1169), .I3(n2971), .I4(n2972), .O(n2973));
  LUT3 #(.INIT(8'h96)) lut_n2974 (.I0(n2962), .I1(n2965), .I2(n2966), .O(n2974));
  LUT3 #(.INIT(8'hE8)) lut_n2975 (.I0(n2970), .I1(n2973), .I2(n2974), .O(n2975));
  LUT3 #(.INIT(8'h96)) lut_n2976 (.I0(n2941), .I1(n2949), .I2(n2950), .O(n2976));
  LUT3 #(.INIT(8'hE8)) lut_n2977 (.I0(n2967), .I1(n2975), .I2(n2976), .O(n2977));
  LUT3 #(.INIT(8'hE8)) lut_n2978 (.I0(x1176), .I1(x1177), .I2(x1178), .O(n2978));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2979 (.I0(x1167), .I1(x1168), .I2(x1169), .I3(n2971), .I4(n2972), .O(n2979));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2980 (.I0(x1173), .I1(x1174), .I2(x1175), .I3(n2978), .I4(n2979), .O(n2980));
  LUT3 #(.INIT(8'hE8)) lut_n2981 (.I0(x1182), .I1(x1183), .I2(x1184), .O(n2981));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2982 (.I0(x1173), .I1(x1174), .I2(x1175), .I3(n2978), .I4(n2979), .O(n2982));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2983 (.I0(x1179), .I1(x1180), .I2(x1181), .I3(n2981), .I4(n2982), .O(n2983));
  LUT3 #(.INIT(8'h96)) lut_n2984 (.I0(n2970), .I1(n2973), .I2(n2974), .O(n2984));
  LUT3 #(.INIT(8'hE8)) lut_n2985 (.I0(n2980), .I1(n2983), .I2(n2984), .O(n2985));
  LUT3 #(.INIT(8'hE8)) lut_n2986 (.I0(x1188), .I1(x1189), .I2(x1190), .O(n2986));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2987 (.I0(x1179), .I1(x1180), .I2(x1181), .I3(n2981), .I4(n2982), .O(n2987));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2988 (.I0(x1185), .I1(x1186), .I2(x1187), .I3(n2986), .I4(n2987), .O(n2988));
  LUT3 #(.INIT(8'hE8)) lut_n2989 (.I0(x1194), .I1(x1195), .I2(x1196), .O(n2989));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2990 (.I0(x1185), .I1(x1186), .I2(x1187), .I3(n2986), .I4(n2987), .O(n2990));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2991 (.I0(x1191), .I1(x1192), .I2(x1193), .I3(n2989), .I4(n2990), .O(n2991));
  LUT3 #(.INIT(8'h96)) lut_n2992 (.I0(n2980), .I1(n2983), .I2(n2984), .O(n2992));
  LUT3 #(.INIT(8'hE8)) lut_n2993 (.I0(n2988), .I1(n2991), .I2(n2992), .O(n2993));
  LUT3 #(.INIT(8'h96)) lut_n2994 (.I0(n2967), .I1(n2975), .I2(n2976), .O(n2994));
  LUT3 #(.INIT(8'hE8)) lut_n2995 (.I0(n2985), .I1(n2993), .I2(n2994), .O(n2995));
  LUT3 #(.INIT(8'h96)) lut_n2996 (.I0(n2933), .I1(n2951), .I2(n2952), .O(n2996));
  LUT3 #(.INIT(8'hE8)) lut_n2997 (.I0(n2977), .I1(n2995), .I2(n2996), .O(n2997));
  LUT3 #(.INIT(8'hE8)) lut_n2998 (.I0(x1200), .I1(x1201), .I2(x1202), .O(n2998));
  LUT5 #(.INIT(32'hE81717E8)) lut_n2999 (.I0(x1191), .I1(x1192), .I2(x1193), .I3(n2989), .I4(n2990), .O(n2999));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3000 (.I0(x1197), .I1(x1198), .I2(x1199), .I3(n2998), .I4(n2999), .O(n3000));
  LUT3 #(.INIT(8'hE8)) lut_n3001 (.I0(x1206), .I1(x1207), .I2(x1208), .O(n3001));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3002 (.I0(x1197), .I1(x1198), .I2(x1199), .I3(n2998), .I4(n2999), .O(n3002));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3003 (.I0(x1203), .I1(x1204), .I2(x1205), .I3(n3001), .I4(n3002), .O(n3003));
  LUT3 #(.INIT(8'h96)) lut_n3004 (.I0(n2988), .I1(n2991), .I2(n2992), .O(n3004));
  LUT3 #(.INIT(8'hE8)) lut_n3005 (.I0(n3000), .I1(n3003), .I2(n3004), .O(n3005));
  LUT3 #(.INIT(8'hE8)) lut_n3006 (.I0(x1212), .I1(x1213), .I2(x1214), .O(n3006));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3007 (.I0(x1203), .I1(x1204), .I2(x1205), .I3(n3001), .I4(n3002), .O(n3007));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3008 (.I0(x1209), .I1(x1210), .I2(x1211), .I3(n3006), .I4(n3007), .O(n3008));
  LUT3 #(.INIT(8'hE8)) lut_n3009 (.I0(x1218), .I1(x1219), .I2(x1220), .O(n3009));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3010 (.I0(x1209), .I1(x1210), .I2(x1211), .I3(n3006), .I4(n3007), .O(n3010));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3011 (.I0(x1215), .I1(x1216), .I2(x1217), .I3(n3009), .I4(n3010), .O(n3011));
  LUT3 #(.INIT(8'h96)) lut_n3012 (.I0(n3000), .I1(n3003), .I2(n3004), .O(n3012));
  LUT3 #(.INIT(8'hE8)) lut_n3013 (.I0(n3008), .I1(n3011), .I2(n3012), .O(n3013));
  LUT3 #(.INIT(8'h96)) lut_n3014 (.I0(n2985), .I1(n2993), .I2(n2994), .O(n3014));
  LUT3 #(.INIT(8'hE8)) lut_n3015 (.I0(n3005), .I1(n3013), .I2(n3014), .O(n3015));
  LUT3 #(.INIT(8'hE8)) lut_n3016 (.I0(x1224), .I1(x1225), .I2(x1226), .O(n3016));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3017 (.I0(x1215), .I1(x1216), .I2(x1217), .I3(n3009), .I4(n3010), .O(n3017));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3018 (.I0(x1221), .I1(x1222), .I2(x1223), .I3(n3016), .I4(n3017), .O(n3018));
  LUT3 #(.INIT(8'hE8)) lut_n3019 (.I0(x1230), .I1(x1231), .I2(x1232), .O(n3019));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3020 (.I0(x1221), .I1(x1222), .I2(x1223), .I3(n3016), .I4(n3017), .O(n3020));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3021 (.I0(x1227), .I1(x1228), .I2(x1229), .I3(n3019), .I4(n3020), .O(n3021));
  LUT3 #(.INIT(8'h96)) lut_n3022 (.I0(n3008), .I1(n3011), .I2(n3012), .O(n3022));
  LUT3 #(.INIT(8'hE8)) lut_n3023 (.I0(n3018), .I1(n3021), .I2(n3022), .O(n3023));
  LUT3 #(.INIT(8'hE8)) lut_n3024 (.I0(x1236), .I1(x1237), .I2(x1238), .O(n3024));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3025 (.I0(x1227), .I1(x1228), .I2(x1229), .I3(n3019), .I4(n3020), .O(n3025));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3026 (.I0(x1233), .I1(x1234), .I2(x1235), .I3(n3024), .I4(n3025), .O(n3026));
  LUT3 #(.INIT(8'hE8)) lut_n3027 (.I0(x1242), .I1(x1243), .I2(x1244), .O(n3027));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3028 (.I0(x1233), .I1(x1234), .I2(x1235), .I3(n3024), .I4(n3025), .O(n3028));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3029 (.I0(x1239), .I1(x1240), .I2(x1241), .I3(n3027), .I4(n3028), .O(n3029));
  LUT3 #(.INIT(8'h96)) lut_n3030 (.I0(n3018), .I1(n3021), .I2(n3022), .O(n3030));
  LUT3 #(.INIT(8'hE8)) lut_n3031 (.I0(n3026), .I1(n3029), .I2(n3030), .O(n3031));
  LUT3 #(.INIT(8'h96)) lut_n3032 (.I0(n3005), .I1(n3013), .I2(n3014), .O(n3032));
  LUT3 #(.INIT(8'hE8)) lut_n3033 (.I0(n3023), .I1(n3031), .I2(n3032), .O(n3033));
  LUT3 #(.INIT(8'h96)) lut_n3034 (.I0(n2977), .I1(n2995), .I2(n2996), .O(n3034));
  LUT3 #(.INIT(8'hE8)) lut_n3035 (.I0(n3015), .I1(n3033), .I2(n3034), .O(n3035));
  LUT3 #(.INIT(8'h96)) lut_n3036 (.I0(n2915), .I1(n2953), .I2(n2954), .O(n3036));
  LUT3 #(.INIT(8'hE8)) lut_n3037 (.I0(n2997), .I1(n3035), .I2(n3036), .O(n3037));
  LUT3 #(.INIT(8'hE8)) lut_n3038 (.I0(x1248), .I1(x1249), .I2(x1250), .O(n3038));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3039 (.I0(x1239), .I1(x1240), .I2(x1241), .I3(n3027), .I4(n3028), .O(n3039));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3040 (.I0(x1245), .I1(x1246), .I2(x1247), .I3(n3038), .I4(n3039), .O(n3040));
  LUT3 #(.INIT(8'hE8)) lut_n3041 (.I0(x1254), .I1(x1255), .I2(x1256), .O(n3041));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3042 (.I0(x1245), .I1(x1246), .I2(x1247), .I3(n3038), .I4(n3039), .O(n3042));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3043 (.I0(x1251), .I1(x1252), .I2(x1253), .I3(n3041), .I4(n3042), .O(n3043));
  LUT3 #(.INIT(8'h96)) lut_n3044 (.I0(n3026), .I1(n3029), .I2(n3030), .O(n3044));
  LUT3 #(.INIT(8'hE8)) lut_n3045 (.I0(n3040), .I1(n3043), .I2(n3044), .O(n3045));
  LUT3 #(.INIT(8'hE8)) lut_n3046 (.I0(x1260), .I1(x1261), .I2(x1262), .O(n3046));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3047 (.I0(x1251), .I1(x1252), .I2(x1253), .I3(n3041), .I4(n3042), .O(n3047));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3048 (.I0(x1257), .I1(x1258), .I2(x1259), .I3(n3046), .I4(n3047), .O(n3048));
  LUT3 #(.INIT(8'hE8)) lut_n3049 (.I0(x1266), .I1(x1267), .I2(x1268), .O(n3049));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3050 (.I0(x1257), .I1(x1258), .I2(x1259), .I3(n3046), .I4(n3047), .O(n3050));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3051 (.I0(x1263), .I1(x1264), .I2(x1265), .I3(n3049), .I4(n3050), .O(n3051));
  LUT3 #(.INIT(8'h96)) lut_n3052 (.I0(n3040), .I1(n3043), .I2(n3044), .O(n3052));
  LUT3 #(.INIT(8'hE8)) lut_n3053 (.I0(n3048), .I1(n3051), .I2(n3052), .O(n3053));
  LUT3 #(.INIT(8'h96)) lut_n3054 (.I0(n3023), .I1(n3031), .I2(n3032), .O(n3054));
  LUT3 #(.INIT(8'hE8)) lut_n3055 (.I0(n3045), .I1(n3053), .I2(n3054), .O(n3055));
  LUT3 #(.INIT(8'hE8)) lut_n3056 (.I0(x1272), .I1(x1273), .I2(x1274), .O(n3056));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3057 (.I0(x1263), .I1(x1264), .I2(x1265), .I3(n3049), .I4(n3050), .O(n3057));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3058 (.I0(x1269), .I1(x1270), .I2(x1271), .I3(n3056), .I4(n3057), .O(n3058));
  LUT3 #(.INIT(8'hE8)) lut_n3059 (.I0(x1278), .I1(x1279), .I2(x1280), .O(n3059));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3060 (.I0(x1269), .I1(x1270), .I2(x1271), .I3(n3056), .I4(n3057), .O(n3060));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3061 (.I0(x1275), .I1(x1276), .I2(x1277), .I3(n3059), .I4(n3060), .O(n3061));
  LUT3 #(.INIT(8'h96)) lut_n3062 (.I0(n3048), .I1(n3051), .I2(n3052), .O(n3062));
  LUT3 #(.INIT(8'hE8)) lut_n3063 (.I0(n3058), .I1(n3061), .I2(n3062), .O(n3063));
  LUT3 #(.INIT(8'hE8)) lut_n3064 (.I0(x1284), .I1(x1285), .I2(x1286), .O(n3064));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3065 (.I0(x1275), .I1(x1276), .I2(x1277), .I3(n3059), .I4(n3060), .O(n3065));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3066 (.I0(x1281), .I1(x1282), .I2(x1283), .I3(n3064), .I4(n3065), .O(n3066));
  LUT3 #(.INIT(8'hE8)) lut_n3067 (.I0(x1290), .I1(x1291), .I2(x1292), .O(n3067));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3068 (.I0(x1281), .I1(x1282), .I2(x1283), .I3(n3064), .I4(n3065), .O(n3068));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3069 (.I0(x1287), .I1(x1288), .I2(x1289), .I3(n3067), .I4(n3068), .O(n3069));
  LUT3 #(.INIT(8'h96)) lut_n3070 (.I0(n3058), .I1(n3061), .I2(n3062), .O(n3070));
  LUT3 #(.INIT(8'hE8)) lut_n3071 (.I0(n3066), .I1(n3069), .I2(n3070), .O(n3071));
  LUT3 #(.INIT(8'h96)) lut_n3072 (.I0(n3045), .I1(n3053), .I2(n3054), .O(n3072));
  LUT3 #(.INIT(8'hE8)) lut_n3073 (.I0(n3063), .I1(n3071), .I2(n3072), .O(n3073));
  LUT3 #(.INIT(8'h96)) lut_n3074 (.I0(n3015), .I1(n3033), .I2(n3034), .O(n3074));
  LUT3 #(.INIT(8'hE8)) lut_n3075 (.I0(n3055), .I1(n3073), .I2(n3074), .O(n3075));
  LUT3 #(.INIT(8'hE8)) lut_n3076 (.I0(x1296), .I1(x1297), .I2(x1298), .O(n3076));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3077 (.I0(x1287), .I1(x1288), .I2(x1289), .I3(n3067), .I4(n3068), .O(n3077));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3078 (.I0(x1293), .I1(x1294), .I2(x1295), .I3(n3076), .I4(n3077), .O(n3078));
  LUT3 #(.INIT(8'hE8)) lut_n3079 (.I0(x1302), .I1(x1303), .I2(x1304), .O(n3079));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3080 (.I0(x1293), .I1(x1294), .I2(x1295), .I3(n3076), .I4(n3077), .O(n3080));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3081 (.I0(x1299), .I1(x1300), .I2(x1301), .I3(n3079), .I4(n3080), .O(n3081));
  LUT3 #(.INIT(8'h96)) lut_n3082 (.I0(n3066), .I1(n3069), .I2(n3070), .O(n3082));
  LUT3 #(.INIT(8'hE8)) lut_n3083 (.I0(n3078), .I1(n3081), .I2(n3082), .O(n3083));
  LUT3 #(.INIT(8'hE8)) lut_n3084 (.I0(x1308), .I1(x1309), .I2(x1310), .O(n3084));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3085 (.I0(x1299), .I1(x1300), .I2(x1301), .I3(n3079), .I4(n3080), .O(n3085));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3086 (.I0(x1305), .I1(x1306), .I2(x1307), .I3(n3084), .I4(n3085), .O(n3086));
  LUT3 #(.INIT(8'hE8)) lut_n3087 (.I0(x1314), .I1(x1315), .I2(x1316), .O(n3087));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3088 (.I0(x1305), .I1(x1306), .I2(x1307), .I3(n3084), .I4(n3085), .O(n3088));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3089 (.I0(x1311), .I1(x1312), .I2(x1313), .I3(n3087), .I4(n3088), .O(n3089));
  LUT3 #(.INIT(8'h96)) lut_n3090 (.I0(n3078), .I1(n3081), .I2(n3082), .O(n3090));
  LUT3 #(.INIT(8'hE8)) lut_n3091 (.I0(n3086), .I1(n3089), .I2(n3090), .O(n3091));
  LUT3 #(.INIT(8'h96)) lut_n3092 (.I0(n3063), .I1(n3071), .I2(n3072), .O(n3092));
  LUT3 #(.INIT(8'hE8)) lut_n3093 (.I0(n3083), .I1(n3091), .I2(n3092), .O(n3093));
  LUT3 #(.INIT(8'hE8)) lut_n3094 (.I0(x1320), .I1(x1321), .I2(x1322), .O(n3094));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3095 (.I0(x1311), .I1(x1312), .I2(x1313), .I3(n3087), .I4(n3088), .O(n3095));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3096 (.I0(x1317), .I1(x1318), .I2(x1319), .I3(n3094), .I4(n3095), .O(n3096));
  LUT3 #(.INIT(8'hE8)) lut_n3097 (.I0(x1326), .I1(x1327), .I2(x1328), .O(n3097));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3098 (.I0(x1317), .I1(x1318), .I2(x1319), .I3(n3094), .I4(n3095), .O(n3098));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3099 (.I0(x1323), .I1(x1324), .I2(x1325), .I3(n3097), .I4(n3098), .O(n3099));
  LUT3 #(.INIT(8'h96)) lut_n3100 (.I0(n3086), .I1(n3089), .I2(n3090), .O(n3100));
  LUT3 #(.INIT(8'hE8)) lut_n3101 (.I0(n3096), .I1(n3099), .I2(n3100), .O(n3101));
  LUT3 #(.INIT(8'hE8)) lut_n3102 (.I0(x1332), .I1(x1333), .I2(x1334), .O(n3102));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3103 (.I0(x1323), .I1(x1324), .I2(x1325), .I3(n3097), .I4(n3098), .O(n3103));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3104 (.I0(x1329), .I1(x1330), .I2(x1331), .I3(n3102), .I4(n3103), .O(n3104));
  LUT3 #(.INIT(8'hE8)) lut_n3105 (.I0(x1338), .I1(x1339), .I2(x1340), .O(n3105));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3106 (.I0(x1329), .I1(x1330), .I2(x1331), .I3(n3102), .I4(n3103), .O(n3106));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3107 (.I0(x1335), .I1(x1336), .I2(x1337), .I3(n3105), .I4(n3106), .O(n3107));
  LUT3 #(.INIT(8'h96)) lut_n3108 (.I0(n3096), .I1(n3099), .I2(n3100), .O(n3108));
  LUT3 #(.INIT(8'hE8)) lut_n3109 (.I0(n3104), .I1(n3107), .I2(n3108), .O(n3109));
  LUT3 #(.INIT(8'h96)) lut_n3110 (.I0(n3083), .I1(n3091), .I2(n3092), .O(n3110));
  LUT3 #(.INIT(8'hE8)) lut_n3111 (.I0(n3101), .I1(n3109), .I2(n3110), .O(n3111));
  LUT3 #(.INIT(8'h96)) lut_n3112 (.I0(n3055), .I1(n3073), .I2(n3074), .O(n3112));
  LUT3 #(.INIT(8'hE8)) lut_n3113 (.I0(n3093), .I1(n3111), .I2(n3112), .O(n3113));
  LUT3 #(.INIT(8'h96)) lut_n3114 (.I0(n2997), .I1(n3035), .I2(n3036), .O(n3114));
  LUT3 #(.INIT(8'hE8)) lut_n3115 (.I0(n3075), .I1(n3113), .I2(n3114), .O(n3115));
  LUT3 #(.INIT(8'h96)) lut_n3116 (.I0(n2877), .I1(n2955), .I2(n2956), .O(n3116));
  LUT3 #(.INIT(8'hE8)) lut_n3117 (.I0(n3037), .I1(n3115), .I2(n3116), .O(n3117));
  LUT3 #(.INIT(8'hE8)) lut_n3118 (.I0(x1344), .I1(x1345), .I2(x1346), .O(n3118));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3119 (.I0(x1335), .I1(x1336), .I2(x1337), .I3(n3105), .I4(n3106), .O(n3119));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3120 (.I0(x1341), .I1(x1342), .I2(x1343), .I3(n3118), .I4(n3119), .O(n3120));
  LUT3 #(.INIT(8'hE8)) lut_n3121 (.I0(x1350), .I1(x1351), .I2(x1352), .O(n3121));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3122 (.I0(x1341), .I1(x1342), .I2(x1343), .I3(n3118), .I4(n3119), .O(n3122));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3123 (.I0(x1347), .I1(x1348), .I2(x1349), .I3(n3121), .I4(n3122), .O(n3123));
  LUT3 #(.INIT(8'h96)) lut_n3124 (.I0(n3104), .I1(n3107), .I2(n3108), .O(n3124));
  LUT3 #(.INIT(8'hE8)) lut_n3125 (.I0(n3120), .I1(n3123), .I2(n3124), .O(n3125));
  LUT3 #(.INIT(8'hE8)) lut_n3126 (.I0(x1356), .I1(x1357), .I2(x1358), .O(n3126));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3127 (.I0(x1347), .I1(x1348), .I2(x1349), .I3(n3121), .I4(n3122), .O(n3127));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3128 (.I0(x1353), .I1(x1354), .I2(x1355), .I3(n3126), .I4(n3127), .O(n3128));
  LUT3 #(.INIT(8'hE8)) lut_n3129 (.I0(x1362), .I1(x1363), .I2(x1364), .O(n3129));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3130 (.I0(x1353), .I1(x1354), .I2(x1355), .I3(n3126), .I4(n3127), .O(n3130));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3131 (.I0(x1359), .I1(x1360), .I2(x1361), .I3(n3129), .I4(n3130), .O(n3131));
  LUT3 #(.INIT(8'h96)) lut_n3132 (.I0(n3120), .I1(n3123), .I2(n3124), .O(n3132));
  LUT3 #(.INIT(8'hE8)) lut_n3133 (.I0(n3128), .I1(n3131), .I2(n3132), .O(n3133));
  LUT3 #(.INIT(8'h96)) lut_n3134 (.I0(n3101), .I1(n3109), .I2(n3110), .O(n3134));
  LUT3 #(.INIT(8'hE8)) lut_n3135 (.I0(n3125), .I1(n3133), .I2(n3134), .O(n3135));
  LUT3 #(.INIT(8'hE8)) lut_n3136 (.I0(x1368), .I1(x1369), .I2(x1370), .O(n3136));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3137 (.I0(x1359), .I1(x1360), .I2(x1361), .I3(n3129), .I4(n3130), .O(n3137));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3138 (.I0(x1365), .I1(x1366), .I2(x1367), .I3(n3136), .I4(n3137), .O(n3138));
  LUT3 #(.INIT(8'hE8)) lut_n3139 (.I0(x1374), .I1(x1375), .I2(x1376), .O(n3139));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3140 (.I0(x1365), .I1(x1366), .I2(x1367), .I3(n3136), .I4(n3137), .O(n3140));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3141 (.I0(x1371), .I1(x1372), .I2(x1373), .I3(n3139), .I4(n3140), .O(n3141));
  LUT3 #(.INIT(8'h96)) lut_n3142 (.I0(n3128), .I1(n3131), .I2(n3132), .O(n3142));
  LUT3 #(.INIT(8'hE8)) lut_n3143 (.I0(n3138), .I1(n3141), .I2(n3142), .O(n3143));
  LUT3 #(.INIT(8'hE8)) lut_n3144 (.I0(x1380), .I1(x1381), .I2(x1382), .O(n3144));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3145 (.I0(x1371), .I1(x1372), .I2(x1373), .I3(n3139), .I4(n3140), .O(n3145));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3146 (.I0(x1377), .I1(x1378), .I2(x1379), .I3(n3144), .I4(n3145), .O(n3146));
  LUT3 #(.INIT(8'hE8)) lut_n3147 (.I0(x1386), .I1(x1387), .I2(x1388), .O(n3147));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3148 (.I0(x1377), .I1(x1378), .I2(x1379), .I3(n3144), .I4(n3145), .O(n3148));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3149 (.I0(x1383), .I1(x1384), .I2(x1385), .I3(n3147), .I4(n3148), .O(n3149));
  LUT3 #(.INIT(8'h96)) lut_n3150 (.I0(n3138), .I1(n3141), .I2(n3142), .O(n3150));
  LUT3 #(.INIT(8'hE8)) lut_n3151 (.I0(n3146), .I1(n3149), .I2(n3150), .O(n3151));
  LUT3 #(.INIT(8'h96)) lut_n3152 (.I0(n3125), .I1(n3133), .I2(n3134), .O(n3152));
  LUT3 #(.INIT(8'hE8)) lut_n3153 (.I0(n3143), .I1(n3151), .I2(n3152), .O(n3153));
  LUT3 #(.INIT(8'h96)) lut_n3154 (.I0(n3093), .I1(n3111), .I2(n3112), .O(n3154));
  LUT3 #(.INIT(8'hE8)) lut_n3155 (.I0(n3135), .I1(n3153), .I2(n3154), .O(n3155));
  LUT3 #(.INIT(8'hE8)) lut_n3156 (.I0(x1392), .I1(x1393), .I2(x1394), .O(n3156));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3157 (.I0(x1383), .I1(x1384), .I2(x1385), .I3(n3147), .I4(n3148), .O(n3157));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3158 (.I0(x1389), .I1(x1390), .I2(x1391), .I3(n3156), .I4(n3157), .O(n3158));
  LUT3 #(.INIT(8'hE8)) lut_n3159 (.I0(x1398), .I1(x1399), .I2(x1400), .O(n3159));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3160 (.I0(x1389), .I1(x1390), .I2(x1391), .I3(n3156), .I4(n3157), .O(n3160));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3161 (.I0(x1395), .I1(x1396), .I2(x1397), .I3(n3159), .I4(n3160), .O(n3161));
  LUT3 #(.INIT(8'h96)) lut_n3162 (.I0(n3146), .I1(n3149), .I2(n3150), .O(n3162));
  LUT3 #(.INIT(8'hE8)) lut_n3163 (.I0(n3158), .I1(n3161), .I2(n3162), .O(n3163));
  LUT3 #(.INIT(8'hE8)) lut_n3164 (.I0(x1404), .I1(x1405), .I2(x1406), .O(n3164));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3165 (.I0(x1395), .I1(x1396), .I2(x1397), .I3(n3159), .I4(n3160), .O(n3165));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3166 (.I0(x1401), .I1(x1402), .I2(x1403), .I3(n3164), .I4(n3165), .O(n3166));
  LUT3 #(.INIT(8'hE8)) lut_n3167 (.I0(x1410), .I1(x1411), .I2(x1412), .O(n3167));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3168 (.I0(x1401), .I1(x1402), .I2(x1403), .I3(n3164), .I4(n3165), .O(n3168));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3169 (.I0(x1407), .I1(x1408), .I2(x1409), .I3(n3167), .I4(n3168), .O(n3169));
  LUT3 #(.INIT(8'h96)) lut_n3170 (.I0(n3158), .I1(n3161), .I2(n3162), .O(n3170));
  LUT3 #(.INIT(8'hE8)) lut_n3171 (.I0(n3166), .I1(n3169), .I2(n3170), .O(n3171));
  LUT3 #(.INIT(8'h96)) lut_n3172 (.I0(n3143), .I1(n3151), .I2(n3152), .O(n3172));
  LUT3 #(.INIT(8'hE8)) lut_n3173 (.I0(n3163), .I1(n3171), .I2(n3172), .O(n3173));
  LUT3 #(.INIT(8'hE8)) lut_n3174 (.I0(x1416), .I1(x1417), .I2(x1418), .O(n3174));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3175 (.I0(x1407), .I1(x1408), .I2(x1409), .I3(n3167), .I4(n3168), .O(n3175));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3176 (.I0(x1413), .I1(x1414), .I2(x1415), .I3(n3174), .I4(n3175), .O(n3176));
  LUT3 #(.INIT(8'hE8)) lut_n3177 (.I0(x1422), .I1(x1423), .I2(x1424), .O(n3177));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3178 (.I0(x1413), .I1(x1414), .I2(x1415), .I3(n3174), .I4(n3175), .O(n3178));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3179 (.I0(x1419), .I1(x1420), .I2(x1421), .I3(n3177), .I4(n3178), .O(n3179));
  LUT3 #(.INIT(8'h96)) lut_n3180 (.I0(n3166), .I1(n3169), .I2(n3170), .O(n3180));
  LUT3 #(.INIT(8'hE8)) lut_n3181 (.I0(n3176), .I1(n3179), .I2(n3180), .O(n3181));
  LUT3 #(.INIT(8'hE8)) lut_n3182 (.I0(x1428), .I1(x1429), .I2(x1430), .O(n3182));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3183 (.I0(x1419), .I1(x1420), .I2(x1421), .I3(n3177), .I4(n3178), .O(n3183));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3184 (.I0(x1425), .I1(x1426), .I2(x1427), .I3(n3182), .I4(n3183), .O(n3184));
  LUT3 #(.INIT(8'hE8)) lut_n3185 (.I0(x1434), .I1(x1435), .I2(x1436), .O(n3185));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3186 (.I0(x1425), .I1(x1426), .I2(x1427), .I3(n3182), .I4(n3183), .O(n3186));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3187 (.I0(x1431), .I1(x1432), .I2(x1433), .I3(n3185), .I4(n3186), .O(n3187));
  LUT3 #(.INIT(8'h96)) lut_n3188 (.I0(n3176), .I1(n3179), .I2(n3180), .O(n3188));
  LUT3 #(.INIT(8'hE8)) lut_n3189 (.I0(n3184), .I1(n3187), .I2(n3188), .O(n3189));
  LUT3 #(.INIT(8'h96)) lut_n3190 (.I0(n3163), .I1(n3171), .I2(n3172), .O(n3190));
  LUT3 #(.INIT(8'hE8)) lut_n3191 (.I0(n3181), .I1(n3189), .I2(n3190), .O(n3191));
  LUT3 #(.INIT(8'h96)) lut_n3192 (.I0(n3135), .I1(n3153), .I2(n3154), .O(n3192));
  LUT3 #(.INIT(8'hE8)) lut_n3193 (.I0(n3173), .I1(n3191), .I2(n3192), .O(n3193));
  LUT3 #(.INIT(8'h96)) lut_n3194 (.I0(n3075), .I1(n3113), .I2(n3114), .O(n3194));
  LUT3 #(.INIT(8'hE8)) lut_n3195 (.I0(n3155), .I1(n3193), .I2(n3194), .O(n3195));
  LUT3 #(.INIT(8'hE8)) lut_n3196 (.I0(x1440), .I1(x1441), .I2(x1442), .O(n3196));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3197 (.I0(x1431), .I1(x1432), .I2(x1433), .I3(n3185), .I4(n3186), .O(n3197));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3198 (.I0(x1437), .I1(x1438), .I2(x1439), .I3(n3196), .I4(n3197), .O(n3198));
  LUT3 #(.INIT(8'hE8)) lut_n3199 (.I0(x1446), .I1(x1447), .I2(x1448), .O(n3199));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3200 (.I0(x1437), .I1(x1438), .I2(x1439), .I3(n3196), .I4(n3197), .O(n3200));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3201 (.I0(x1443), .I1(x1444), .I2(x1445), .I3(n3199), .I4(n3200), .O(n3201));
  LUT3 #(.INIT(8'h96)) lut_n3202 (.I0(n3184), .I1(n3187), .I2(n3188), .O(n3202));
  LUT3 #(.INIT(8'hE8)) lut_n3203 (.I0(n3198), .I1(n3201), .I2(n3202), .O(n3203));
  LUT3 #(.INIT(8'hE8)) lut_n3204 (.I0(x1452), .I1(x1453), .I2(x1454), .O(n3204));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3205 (.I0(x1443), .I1(x1444), .I2(x1445), .I3(n3199), .I4(n3200), .O(n3205));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3206 (.I0(x1449), .I1(x1450), .I2(x1451), .I3(n3204), .I4(n3205), .O(n3206));
  LUT3 #(.INIT(8'hE8)) lut_n3207 (.I0(x1458), .I1(x1459), .I2(x1460), .O(n3207));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3208 (.I0(x1449), .I1(x1450), .I2(x1451), .I3(n3204), .I4(n3205), .O(n3208));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3209 (.I0(x1455), .I1(x1456), .I2(x1457), .I3(n3207), .I4(n3208), .O(n3209));
  LUT3 #(.INIT(8'h96)) lut_n3210 (.I0(n3198), .I1(n3201), .I2(n3202), .O(n3210));
  LUT3 #(.INIT(8'hE8)) lut_n3211 (.I0(n3206), .I1(n3209), .I2(n3210), .O(n3211));
  LUT3 #(.INIT(8'h96)) lut_n3212 (.I0(n3181), .I1(n3189), .I2(n3190), .O(n3212));
  LUT3 #(.INIT(8'hE8)) lut_n3213 (.I0(n3203), .I1(n3211), .I2(n3212), .O(n3213));
  LUT3 #(.INIT(8'hE8)) lut_n3214 (.I0(x1464), .I1(x1465), .I2(x1466), .O(n3214));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3215 (.I0(x1455), .I1(x1456), .I2(x1457), .I3(n3207), .I4(n3208), .O(n3215));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3216 (.I0(x1461), .I1(x1462), .I2(x1463), .I3(n3214), .I4(n3215), .O(n3216));
  LUT3 #(.INIT(8'hE8)) lut_n3217 (.I0(x1470), .I1(x1471), .I2(x1472), .O(n3217));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3218 (.I0(x1461), .I1(x1462), .I2(x1463), .I3(n3214), .I4(n3215), .O(n3218));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3219 (.I0(x1467), .I1(x1468), .I2(x1469), .I3(n3217), .I4(n3218), .O(n3219));
  LUT3 #(.INIT(8'h96)) lut_n3220 (.I0(n3206), .I1(n3209), .I2(n3210), .O(n3220));
  LUT3 #(.INIT(8'hE8)) lut_n3221 (.I0(n3216), .I1(n3219), .I2(n3220), .O(n3221));
  LUT3 #(.INIT(8'hE8)) lut_n3222 (.I0(x1476), .I1(x1477), .I2(x1478), .O(n3222));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3223 (.I0(x1467), .I1(x1468), .I2(x1469), .I3(n3217), .I4(n3218), .O(n3223));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3224 (.I0(x1473), .I1(x1474), .I2(x1475), .I3(n3222), .I4(n3223), .O(n3224));
  LUT3 #(.INIT(8'hE8)) lut_n3225 (.I0(x1482), .I1(x1483), .I2(x1484), .O(n3225));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3226 (.I0(x1473), .I1(x1474), .I2(x1475), .I3(n3222), .I4(n3223), .O(n3226));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3227 (.I0(x1479), .I1(x1480), .I2(x1481), .I3(n3225), .I4(n3226), .O(n3227));
  LUT3 #(.INIT(8'h96)) lut_n3228 (.I0(n3216), .I1(n3219), .I2(n3220), .O(n3228));
  LUT3 #(.INIT(8'hE8)) lut_n3229 (.I0(n3224), .I1(n3227), .I2(n3228), .O(n3229));
  LUT3 #(.INIT(8'h96)) lut_n3230 (.I0(n3203), .I1(n3211), .I2(n3212), .O(n3230));
  LUT3 #(.INIT(8'hE8)) lut_n3231 (.I0(n3221), .I1(n3229), .I2(n3230), .O(n3231));
  LUT3 #(.INIT(8'h96)) lut_n3232 (.I0(n3173), .I1(n3191), .I2(n3192), .O(n3232));
  LUT3 #(.INIT(8'hE8)) lut_n3233 (.I0(n3213), .I1(n3231), .I2(n3232), .O(n3233));
  LUT3 #(.INIT(8'hE8)) lut_n3234 (.I0(x1488), .I1(x1489), .I2(x1490), .O(n3234));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3235 (.I0(x1479), .I1(x1480), .I2(x1481), .I3(n3225), .I4(n3226), .O(n3235));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3236 (.I0(x1485), .I1(x1486), .I2(x1487), .I3(n3234), .I4(n3235), .O(n3236));
  LUT3 #(.INIT(8'hE8)) lut_n3237 (.I0(x1494), .I1(x1495), .I2(x1496), .O(n3237));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3238 (.I0(x1485), .I1(x1486), .I2(x1487), .I3(n3234), .I4(n3235), .O(n3238));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3239 (.I0(x1491), .I1(x1492), .I2(x1493), .I3(n3237), .I4(n3238), .O(n3239));
  LUT3 #(.INIT(8'h96)) lut_n3240 (.I0(n3224), .I1(n3227), .I2(n3228), .O(n3240));
  LUT3 #(.INIT(8'hE8)) lut_n3241 (.I0(n3236), .I1(n3239), .I2(n3240), .O(n3241));
  LUT3 #(.INIT(8'hE8)) lut_n3242 (.I0(x1500), .I1(x1501), .I2(x1502), .O(n3242));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3243 (.I0(x1491), .I1(x1492), .I2(x1493), .I3(n3237), .I4(n3238), .O(n3243));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3244 (.I0(x1497), .I1(x1498), .I2(x1499), .I3(n3242), .I4(n3243), .O(n3244));
  LUT3 #(.INIT(8'hE8)) lut_n3245 (.I0(x1506), .I1(x1507), .I2(x1508), .O(n3245));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3246 (.I0(x1497), .I1(x1498), .I2(x1499), .I3(n3242), .I4(n3243), .O(n3246));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3247 (.I0(x1503), .I1(x1504), .I2(x1505), .I3(n3245), .I4(n3246), .O(n3247));
  LUT3 #(.INIT(8'h96)) lut_n3248 (.I0(n3236), .I1(n3239), .I2(n3240), .O(n3248));
  LUT3 #(.INIT(8'hE8)) lut_n3249 (.I0(n3244), .I1(n3247), .I2(n3248), .O(n3249));
  LUT3 #(.INIT(8'h96)) lut_n3250 (.I0(n3221), .I1(n3229), .I2(n3230), .O(n3250));
  LUT3 #(.INIT(8'hE8)) lut_n3251 (.I0(n3241), .I1(n3249), .I2(n3250), .O(n3251));
  LUT3 #(.INIT(8'hE8)) lut_n3252 (.I0(x1512), .I1(x1513), .I2(x1514), .O(n3252));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3253 (.I0(x1503), .I1(x1504), .I2(x1505), .I3(n3245), .I4(n3246), .O(n3253));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3254 (.I0(x1509), .I1(x1510), .I2(x1511), .I3(n3252), .I4(n3253), .O(n3254));
  LUT3 #(.INIT(8'hE8)) lut_n3255 (.I0(x1518), .I1(x1519), .I2(x1520), .O(n3255));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3256 (.I0(x1509), .I1(x1510), .I2(x1511), .I3(n3252), .I4(n3253), .O(n3256));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3257 (.I0(x1515), .I1(x1516), .I2(x1517), .I3(n3255), .I4(n3256), .O(n3257));
  LUT3 #(.INIT(8'h96)) lut_n3258 (.I0(n3244), .I1(n3247), .I2(n3248), .O(n3258));
  LUT3 #(.INIT(8'hE8)) lut_n3259 (.I0(n3254), .I1(n3257), .I2(n3258), .O(n3259));
  LUT3 #(.INIT(8'hE8)) lut_n3260 (.I0(x1524), .I1(x1525), .I2(x1526), .O(n3260));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3261 (.I0(x1515), .I1(x1516), .I2(x1517), .I3(n3255), .I4(n3256), .O(n3261));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3262 (.I0(x1521), .I1(x1522), .I2(x1523), .I3(n3260), .I4(n3261), .O(n3262));
  LUT3 #(.INIT(8'hE8)) lut_n3263 (.I0(x1530), .I1(x1531), .I2(x1532), .O(n3263));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3264 (.I0(x1521), .I1(x1522), .I2(x1523), .I3(n3260), .I4(n3261), .O(n3264));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3265 (.I0(x1527), .I1(x1528), .I2(x1529), .I3(n3263), .I4(n3264), .O(n3265));
  LUT3 #(.INIT(8'h96)) lut_n3266 (.I0(n3254), .I1(n3257), .I2(n3258), .O(n3266));
  LUT3 #(.INIT(8'hE8)) lut_n3267 (.I0(n3262), .I1(n3265), .I2(n3266), .O(n3267));
  LUT3 #(.INIT(8'h96)) lut_n3268 (.I0(n3241), .I1(n3249), .I2(n3250), .O(n3268));
  LUT3 #(.INIT(8'hE8)) lut_n3269 (.I0(n3259), .I1(n3267), .I2(n3268), .O(n3269));
  LUT3 #(.INIT(8'h96)) lut_n3270 (.I0(n3213), .I1(n3231), .I2(n3232), .O(n3270));
  LUT3 #(.INIT(8'hE8)) lut_n3271 (.I0(n3251), .I1(n3269), .I2(n3270), .O(n3271));
  LUT3 #(.INIT(8'h96)) lut_n3272 (.I0(n3155), .I1(n3193), .I2(n3194), .O(n3272));
  LUT3 #(.INIT(8'hE8)) lut_n3273 (.I0(n3233), .I1(n3271), .I2(n3272), .O(n3273));
  LUT3 #(.INIT(8'h96)) lut_n3274 (.I0(n3037), .I1(n3115), .I2(n3116), .O(n3274));
  LUT3 #(.INIT(8'hE8)) lut_n3275 (.I0(n3195), .I1(n3273), .I2(n3274), .O(n3275));
  LUT3 #(.INIT(8'h96)) lut_n3276 (.I0(n2799), .I1(n2957), .I2(n2958), .O(n3276));
  LUT3 #(.INIT(8'hE8)) lut_n3277 (.I0(n3117), .I1(n3275), .I2(n3276), .O(n3277));
  LUT3 #(.INIT(8'hE8)) lut_n3278 (.I0(n2641), .I1(n2959), .I2(n3277), .O(n3278));
  LUT3 #(.INIT(8'hE8)) lut_n3279 (.I0(x1536), .I1(x1537), .I2(x1538), .O(n3279));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3280 (.I0(x1527), .I1(x1528), .I2(x1529), .I3(n3263), .I4(n3264), .O(n3280));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3281 (.I0(x1533), .I1(x1534), .I2(x1535), .I3(n3279), .I4(n3280), .O(n3281));
  LUT3 #(.INIT(8'hE8)) lut_n3282 (.I0(x1542), .I1(x1543), .I2(x1544), .O(n3282));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3283 (.I0(x1533), .I1(x1534), .I2(x1535), .I3(n3279), .I4(n3280), .O(n3283));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3284 (.I0(x1539), .I1(x1540), .I2(x1541), .I3(n3282), .I4(n3283), .O(n3284));
  LUT3 #(.INIT(8'h96)) lut_n3285 (.I0(n3262), .I1(n3265), .I2(n3266), .O(n3285));
  LUT3 #(.INIT(8'hE8)) lut_n3286 (.I0(n3281), .I1(n3284), .I2(n3285), .O(n3286));
  LUT3 #(.INIT(8'hE8)) lut_n3287 (.I0(x1548), .I1(x1549), .I2(x1550), .O(n3287));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3288 (.I0(x1539), .I1(x1540), .I2(x1541), .I3(n3282), .I4(n3283), .O(n3288));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3289 (.I0(x1545), .I1(x1546), .I2(x1547), .I3(n3287), .I4(n3288), .O(n3289));
  LUT3 #(.INIT(8'hE8)) lut_n3290 (.I0(x1554), .I1(x1555), .I2(x1556), .O(n3290));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3291 (.I0(x1545), .I1(x1546), .I2(x1547), .I3(n3287), .I4(n3288), .O(n3291));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3292 (.I0(x1551), .I1(x1552), .I2(x1553), .I3(n3290), .I4(n3291), .O(n3292));
  LUT3 #(.INIT(8'h96)) lut_n3293 (.I0(n3281), .I1(n3284), .I2(n3285), .O(n3293));
  LUT3 #(.INIT(8'hE8)) lut_n3294 (.I0(n3289), .I1(n3292), .I2(n3293), .O(n3294));
  LUT3 #(.INIT(8'h96)) lut_n3295 (.I0(n3259), .I1(n3267), .I2(n3268), .O(n3295));
  LUT3 #(.INIT(8'hE8)) lut_n3296 (.I0(n3286), .I1(n3294), .I2(n3295), .O(n3296));
  LUT3 #(.INIT(8'hE8)) lut_n3297 (.I0(x1560), .I1(x1561), .I2(x1562), .O(n3297));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3298 (.I0(x1551), .I1(x1552), .I2(x1553), .I3(n3290), .I4(n3291), .O(n3298));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3299 (.I0(x1557), .I1(x1558), .I2(x1559), .I3(n3297), .I4(n3298), .O(n3299));
  LUT3 #(.INIT(8'hE8)) lut_n3300 (.I0(x1566), .I1(x1567), .I2(x1568), .O(n3300));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3301 (.I0(x1557), .I1(x1558), .I2(x1559), .I3(n3297), .I4(n3298), .O(n3301));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3302 (.I0(x1563), .I1(x1564), .I2(x1565), .I3(n3300), .I4(n3301), .O(n3302));
  LUT3 #(.INIT(8'h96)) lut_n3303 (.I0(n3289), .I1(n3292), .I2(n3293), .O(n3303));
  LUT3 #(.INIT(8'hE8)) lut_n3304 (.I0(n3299), .I1(n3302), .I2(n3303), .O(n3304));
  LUT3 #(.INIT(8'hE8)) lut_n3305 (.I0(x1572), .I1(x1573), .I2(x1574), .O(n3305));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3306 (.I0(x1563), .I1(x1564), .I2(x1565), .I3(n3300), .I4(n3301), .O(n3306));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3307 (.I0(x1569), .I1(x1570), .I2(x1571), .I3(n3305), .I4(n3306), .O(n3307));
  LUT3 #(.INIT(8'hE8)) lut_n3308 (.I0(x1578), .I1(x1579), .I2(x1580), .O(n3308));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3309 (.I0(x1569), .I1(x1570), .I2(x1571), .I3(n3305), .I4(n3306), .O(n3309));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3310 (.I0(x1575), .I1(x1576), .I2(x1577), .I3(n3308), .I4(n3309), .O(n3310));
  LUT3 #(.INIT(8'h96)) lut_n3311 (.I0(n3299), .I1(n3302), .I2(n3303), .O(n3311));
  LUT3 #(.INIT(8'hE8)) lut_n3312 (.I0(n3307), .I1(n3310), .I2(n3311), .O(n3312));
  LUT3 #(.INIT(8'h96)) lut_n3313 (.I0(n3286), .I1(n3294), .I2(n3295), .O(n3313));
  LUT3 #(.INIT(8'hE8)) lut_n3314 (.I0(n3304), .I1(n3312), .I2(n3313), .O(n3314));
  LUT3 #(.INIT(8'h96)) lut_n3315 (.I0(n3251), .I1(n3269), .I2(n3270), .O(n3315));
  LUT3 #(.INIT(8'hE8)) lut_n3316 (.I0(n3296), .I1(n3314), .I2(n3315), .O(n3316));
  LUT3 #(.INIT(8'hE8)) lut_n3317 (.I0(x1584), .I1(x1585), .I2(x1586), .O(n3317));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3318 (.I0(x1575), .I1(x1576), .I2(x1577), .I3(n3308), .I4(n3309), .O(n3318));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3319 (.I0(x1581), .I1(x1582), .I2(x1583), .I3(n3317), .I4(n3318), .O(n3319));
  LUT3 #(.INIT(8'hE8)) lut_n3320 (.I0(x1590), .I1(x1591), .I2(x1592), .O(n3320));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3321 (.I0(x1581), .I1(x1582), .I2(x1583), .I3(n3317), .I4(n3318), .O(n3321));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3322 (.I0(x1587), .I1(x1588), .I2(x1589), .I3(n3320), .I4(n3321), .O(n3322));
  LUT3 #(.INIT(8'h96)) lut_n3323 (.I0(n3307), .I1(n3310), .I2(n3311), .O(n3323));
  LUT3 #(.INIT(8'hE8)) lut_n3324 (.I0(n3319), .I1(n3322), .I2(n3323), .O(n3324));
  LUT3 #(.INIT(8'hE8)) lut_n3325 (.I0(x1596), .I1(x1597), .I2(x1598), .O(n3325));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3326 (.I0(x1587), .I1(x1588), .I2(x1589), .I3(n3320), .I4(n3321), .O(n3326));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3327 (.I0(x1593), .I1(x1594), .I2(x1595), .I3(n3325), .I4(n3326), .O(n3327));
  LUT3 #(.INIT(8'hE8)) lut_n3328 (.I0(x1602), .I1(x1603), .I2(x1604), .O(n3328));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3329 (.I0(x1593), .I1(x1594), .I2(x1595), .I3(n3325), .I4(n3326), .O(n3329));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3330 (.I0(x1599), .I1(x1600), .I2(x1601), .I3(n3328), .I4(n3329), .O(n3330));
  LUT3 #(.INIT(8'h96)) lut_n3331 (.I0(n3319), .I1(n3322), .I2(n3323), .O(n3331));
  LUT3 #(.INIT(8'hE8)) lut_n3332 (.I0(n3327), .I1(n3330), .I2(n3331), .O(n3332));
  LUT3 #(.INIT(8'h96)) lut_n3333 (.I0(n3304), .I1(n3312), .I2(n3313), .O(n3333));
  LUT3 #(.INIT(8'hE8)) lut_n3334 (.I0(n3324), .I1(n3332), .I2(n3333), .O(n3334));
  LUT3 #(.INIT(8'hE8)) lut_n3335 (.I0(x1608), .I1(x1609), .I2(x1610), .O(n3335));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3336 (.I0(x1599), .I1(x1600), .I2(x1601), .I3(n3328), .I4(n3329), .O(n3336));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3337 (.I0(x1605), .I1(x1606), .I2(x1607), .I3(n3335), .I4(n3336), .O(n3337));
  LUT3 #(.INIT(8'hE8)) lut_n3338 (.I0(x1614), .I1(x1615), .I2(x1616), .O(n3338));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3339 (.I0(x1605), .I1(x1606), .I2(x1607), .I3(n3335), .I4(n3336), .O(n3339));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3340 (.I0(x1611), .I1(x1612), .I2(x1613), .I3(n3338), .I4(n3339), .O(n3340));
  LUT3 #(.INIT(8'h96)) lut_n3341 (.I0(n3327), .I1(n3330), .I2(n3331), .O(n3341));
  LUT3 #(.INIT(8'hE8)) lut_n3342 (.I0(n3337), .I1(n3340), .I2(n3341), .O(n3342));
  LUT3 #(.INIT(8'hE8)) lut_n3343 (.I0(x1620), .I1(x1621), .I2(x1622), .O(n3343));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3344 (.I0(x1611), .I1(x1612), .I2(x1613), .I3(n3338), .I4(n3339), .O(n3344));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3345 (.I0(x1617), .I1(x1618), .I2(x1619), .I3(n3343), .I4(n3344), .O(n3345));
  LUT3 #(.INIT(8'hE8)) lut_n3346 (.I0(x1626), .I1(x1627), .I2(x1628), .O(n3346));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3347 (.I0(x1617), .I1(x1618), .I2(x1619), .I3(n3343), .I4(n3344), .O(n3347));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3348 (.I0(x1623), .I1(x1624), .I2(x1625), .I3(n3346), .I4(n3347), .O(n3348));
  LUT3 #(.INIT(8'h96)) lut_n3349 (.I0(n3337), .I1(n3340), .I2(n3341), .O(n3349));
  LUT3 #(.INIT(8'hE8)) lut_n3350 (.I0(n3345), .I1(n3348), .I2(n3349), .O(n3350));
  LUT3 #(.INIT(8'h96)) lut_n3351 (.I0(n3324), .I1(n3332), .I2(n3333), .O(n3351));
  LUT3 #(.INIT(8'hE8)) lut_n3352 (.I0(n3342), .I1(n3350), .I2(n3351), .O(n3352));
  LUT3 #(.INIT(8'h96)) lut_n3353 (.I0(n3296), .I1(n3314), .I2(n3315), .O(n3353));
  LUT3 #(.INIT(8'hE8)) lut_n3354 (.I0(n3334), .I1(n3352), .I2(n3353), .O(n3354));
  LUT3 #(.INIT(8'h96)) lut_n3355 (.I0(n3233), .I1(n3271), .I2(n3272), .O(n3355));
  LUT3 #(.INIT(8'hE8)) lut_n3356 (.I0(n3316), .I1(n3354), .I2(n3355), .O(n3356));
  LUT3 #(.INIT(8'hE8)) lut_n3357 (.I0(x1632), .I1(x1633), .I2(x1634), .O(n3357));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3358 (.I0(x1623), .I1(x1624), .I2(x1625), .I3(n3346), .I4(n3347), .O(n3358));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3359 (.I0(x1629), .I1(x1630), .I2(x1631), .I3(n3357), .I4(n3358), .O(n3359));
  LUT3 #(.INIT(8'hE8)) lut_n3360 (.I0(x1638), .I1(x1639), .I2(x1640), .O(n3360));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3361 (.I0(x1629), .I1(x1630), .I2(x1631), .I3(n3357), .I4(n3358), .O(n3361));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3362 (.I0(x1635), .I1(x1636), .I2(x1637), .I3(n3360), .I4(n3361), .O(n3362));
  LUT3 #(.INIT(8'h96)) lut_n3363 (.I0(n3345), .I1(n3348), .I2(n3349), .O(n3363));
  LUT3 #(.INIT(8'hE8)) lut_n3364 (.I0(n3359), .I1(n3362), .I2(n3363), .O(n3364));
  LUT3 #(.INIT(8'hE8)) lut_n3365 (.I0(x1644), .I1(x1645), .I2(x1646), .O(n3365));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3366 (.I0(x1635), .I1(x1636), .I2(x1637), .I3(n3360), .I4(n3361), .O(n3366));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3367 (.I0(x1641), .I1(x1642), .I2(x1643), .I3(n3365), .I4(n3366), .O(n3367));
  LUT3 #(.INIT(8'hE8)) lut_n3368 (.I0(x1650), .I1(x1651), .I2(x1652), .O(n3368));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3369 (.I0(x1641), .I1(x1642), .I2(x1643), .I3(n3365), .I4(n3366), .O(n3369));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3370 (.I0(x1647), .I1(x1648), .I2(x1649), .I3(n3368), .I4(n3369), .O(n3370));
  LUT3 #(.INIT(8'h96)) lut_n3371 (.I0(n3359), .I1(n3362), .I2(n3363), .O(n3371));
  LUT3 #(.INIT(8'hE8)) lut_n3372 (.I0(n3367), .I1(n3370), .I2(n3371), .O(n3372));
  LUT3 #(.INIT(8'h96)) lut_n3373 (.I0(n3342), .I1(n3350), .I2(n3351), .O(n3373));
  LUT3 #(.INIT(8'hE8)) lut_n3374 (.I0(n3364), .I1(n3372), .I2(n3373), .O(n3374));
  LUT3 #(.INIT(8'hE8)) lut_n3375 (.I0(x1656), .I1(x1657), .I2(x1658), .O(n3375));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3376 (.I0(x1647), .I1(x1648), .I2(x1649), .I3(n3368), .I4(n3369), .O(n3376));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3377 (.I0(x1653), .I1(x1654), .I2(x1655), .I3(n3375), .I4(n3376), .O(n3377));
  LUT3 #(.INIT(8'hE8)) lut_n3378 (.I0(x1662), .I1(x1663), .I2(x1664), .O(n3378));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3379 (.I0(x1653), .I1(x1654), .I2(x1655), .I3(n3375), .I4(n3376), .O(n3379));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3380 (.I0(x1659), .I1(x1660), .I2(x1661), .I3(n3378), .I4(n3379), .O(n3380));
  LUT3 #(.INIT(8'h96)) lut_n3381 (.I0(n3367), .I1(n3370), .I2(n3371), .O(n3381));
  LUT3 #(.INIT(8'hE8)) lut_n3382 (.I0(n3377), .I1(n3380), .I2(n3381), .O(n3382));
  LUT3 #(.INIT(8'hE8)) lut_n3383 (.I0(x1668), .I1(x1669), .I2(x1670), .O(n3383));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3384 (.I0(x1659), .I1(x1660), .I2(x1661), .I3(n3378), .I4(n3379), .O(n3384));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3385 (.I0(x1665), .I1(x1666), .I2(x1667), .I3(n3383), .I4(n3384), .O(n3385));
  LUT3 #(.INIT(8'hE8)) lut_n3386 (.I0(x1674), .I1(x1675), .I2(x1676), .O(n3386));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3387 (.I0(x1665), .I1(x1666), .I2(x1667), .I3(n3383), .I4(n3384), .O(n3387));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3388 (.I0(x1671), .I1(x1672), .I2(x1673), .I3(n3386), .I4(n3387), .O(n3388));
  LUT3 #(.INIT(8'h96)) lut_n3389 (.I0(n3377), .I1(n3380), .I2(n3381), .O(n3389));
  LUT3 #(.INIT(8'hE8)) lut_n3390 (.I0(n3385), .I1(n3388), .I2(n3389), .O(n3390));
  LUT3 #(.INIT(8'h96)) lut_n3391 (.I0(n3364), .I1(n3372), .I2(n3373), .O(n3391));
  LUT3 #(.INIT(8'hE8)) lut_n3392 (.I0(n3382), .I1(n3390), .I2(n3391), .O(n3392));
  LUT3 #(.INIT(8'h96)) lut_n3393 (.I0(n3334), .I1(n3352), .I2(n3353), .O(n3393));
  LUT3 #(.INIT(8'hE8)) lut_n3394 (.I0(n3374), .I1(n3392), .I2(n3393), .O(n3394));
  LUT3 #(.INIT(8'hE8)) lut_n3395 (.I0(x1680), .I1(x1681), .I2(x1682), .O(n3395));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3396 (.I0(x1671), .I1(x1672), .I2(x1673), .I3(n3386), .I4(n3387), .O(n3396));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3397 (.I0(x1677), .I1(x1678), .I2(x1679), .I3(n3395), .I4(n3396), .O(n3397));
  LUT3 #(.INIT(8'hE8)) lut_n3398 (.I0(x1686), .I1(x1687), .I2(x1688), .O(n3398));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3399 (.I0(x1677), .I1(x1678), .I2(x1679), .I3(n3395), .I4(n3396), .O(n3399));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3400 (.I0(x1683), .I1(x1684), .I2(x1685), .I3(n3398), .I4(n3399), .O(n3400));
  LUT3 #(.INIT(8'h96)) lut_n3401 (.I0(n3385), .I1(n3388), .I2(n3389), .O(n3401));
  LUT3 #(.INIT(8'hE8)) lut_n3402 (.I0(n3397), .I1(n3400), .I2(n3401), .O(n3402));
  LUT3 #(.INIT(8'hE8)) lut_n3403 (.I0(x1692), .I1(x1693), .I2(x1694), .O(n3403));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3404 (.I0(x1683), .I1(x1684), .I2(x1685), .I3(n3398), .I4(n3399), .O(n3404));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3405 (.I0(x1689), .I1(x1690), .I2(x1691), .I3(n3403), .I4(n3404), .O(n3405));
  LUT3 #(.INIT(8'hE8)) lut_n3406 (.I0(x1698), .I1(x1699), .I2(x1700), .O(n3406));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3407 (.I0(x1689), .I1(x1690), .I2(x1691), .I3(n3403), .I4(n3404), .O(n3407));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3408 (.I0(x1695), .I1(x1696), .I2(x1697), .I3(n3406), .I4(n3407), .O(n3408));
  LUT3 #(.INIT(8'h96)) lut_n3409 (.I0(n3397), .I1(n3400), .I2(n3401), .O(n3409));
  LUT3 #(.INIT(8'hE8)) lut_n3410 (.I0(n3405), .I1(n3408), .I2(n3409), .O(n3410));
  LUT3 #(.INIT(8'h96)) lut_n3411 (.I0(n3382), .I1(n3390), .I2(n3391), .O(n3411));
  LUT3 #(.INIT(8'hE8)) lut_n3412 (.I0(n3402), .I1(n3410), .I2(n3411), .O(n3412));
  LUT3 #(.INIT(8'hE8)) lut_n3413 (.I0(x1704), .I1(x1705), .I2(x1706), .O(n3413));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3414 (.I0(x1695), .I1(x1696), .I2(x1697), .I3(n3406), .I4(n3407), .O(n3414));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3415 (.I0(x1701), .I1(x1702), .I2(x1703), .I3(n3413), .I4(n3414), .O(n3415));
  LUT3 #(.INIT(8'hE8)) lut_n3416 (.I0(x1710), .I1(x1711), .I2(x1712), .O(n3416));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3417 (.I0(x1701), .I1(x1702), .I2(x1703), .I3(n3413), .I4(n3414), .O(n3417));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3418 (.I0(x1707), .I1(x1708), .I2(x1709), .I3(n3416), .I4(n3417), .O(n3418));
  LUT3 #(.INIT(8'h96)) lut_n3419 (.I0(n3405), .I1(n3408), .I2(n3409), .O(n3419));
  LUT3 #(.INIT(8'hE8)) lut_n3420 (.I0(n3415), .I1(n3418), .I2(n3419), .O(n3420));
  LUT3 #(.INIT(8'hE8)) lut_n3421 (.I0(x1716), .I1(x1717), .I2(x1718), .O(n3421));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3422 (.I0(x1707), .I1(x1708), .I2(x1709), .I3(n3416), .I4(n3417), .O(n3422));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3423 (.I0(x1713), .I1(x1714), .I2(x1715), .I3(n3421), .I4(n3422), .O(n3423));
  LUT3 #(.INIT(8'hE8)) lut_n3424 (.I0(x1722), .I1(x1723), .I2(x1724), .O(n3424));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3425 (.I0(x1713), .I1(x1714), .I2(x1715), .I3(n3421), .I4(n3422), .O(n3425));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3426 (.I0(x1719), .I1(x1720), .I2(x1721), .I3(n3424), .I4(n3425), .O(n3426));
  LUT3 #(.INIT(8'h96)) lut_n3427 (.I0(n3415), .I1(n3418), .I2(n3419), .O(n3427));
  LUT3 #(.INIT(8'hE8)) lut_n3428 (.I0(n3423), .I1(n3426), .I2(n3427), .O(n3428));
  LUT3 #(.INIT(8'h96)) lut_n3429 (.I0(n3402), .I1(n3410), .I2(n3411), .O(n3429));
  LUT3 #(.INIT(8'hE8)) lut_n3430 (.I0(n3420), .I1(n3428), .I2(n3429), .O(n3430));
  LUT3 #(.INIT(8'h96)) lut_n3431 (.I0(n3374), .I1(n3392), .I2(n3393), .O(n3431));
  LUT3 #(.INIT(8'hE8)) lut_n3432 (.I0(n3412), .I1(n3430), .I2(n3431), .O(n3432));
  LUT3 #(.INIT(8'h96)) lut_n3433 (.I0(n3316), .I1(n3354), .I2(n3355), .O(n3433));
  LUT3 #(.INIT(8'hE8)) lut_n3434 (.I0(n3394), .I1(n3432), .I2(n3433), .O(n3434));
  LUT3 #(.INIT(8'h96)) lut_n3435 (.I0(n3195), .I1(n3273), .I2(n3274), .O(n3435));
  LUT3 #(.INIT(8'hE8)) lut_n3436 (.I0(n3356), .I1(n3434), .I2(n3435), .O(n3436));
  LUT3 #(.INIT(8'hE8)) lut_n3437 (.I0(x1728), .I1(x1729), .I2(x1730), .O(n3437));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3438 (.I0(x1719), .I1(x1720), .I2(x1721), .I3(n3424), .I4(n3425), .O(n3438));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3439 (.I0(x1725), .I1(x1726), .I2(x1727), .I3(n3437), .I4(n3438), .O(n3439));
  LUT3 #(.INIT(8'hE8)) lut_n3440 (.I0(x1734), .I1(x1735), .I2(x1736), .O(n3440));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3441 (.I0(x1725), .I1(x1726), .I2(x1727), .I3(n3437), .I4(n3438), .O(n3441));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3442 (.I0(x1731), .I1(x1732), .I2(x1733), .I3(n3440), .I4(n3441), .O(n3442));
  LUT3 #(.INIT(8'h96)) lut_n3443 (.I0(n3423), .I1(n3426), .I2(n3427), .O(n3443));
  LUT3 #(.INIT(8'hE8)) lut_n3444 (.I0(n3439), .I1(n3442), .I2(n3443), .O(n3444));
  LUT3 #(.INIT(8'hE8)) lut_n3445 (.I0(x1740), .I1(x1741), .I2(x1742), .O(n3445));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3446 (.I0(x1731), .I1(x1732), .I2(x1733), .I3(n3440), .I4(n3441), .O(n3446));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3447 (.I0(x1737), .I1(x1738), .I2(x1739), .I3(n3445), .I4(n3446), .O(n3447));
  LUT3 #(.INIT(8'hE8)) lut_n3448 (.I0(x1746), .I1(x1747), .I2(x1748), .O(n3448));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3449 (.I0(x1737), .I1(x1738), .I2(x1739), .I3(n3445), .I4(n3446), .O(n3449));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3450 (.I0(x1743), .I1(x1744), .I2(x1745), .I3(n3448), .I4(n3449), .O(n3450));
  LUT3 #(.INIT(8'h96)) lut_n3451 (.I0(n3439), .I1(n3442), .I2(n3443), .O(n3451));
  LUT3 #(.INIT(8'hE8)) lut_n3452 (.I0(n3447), .I1(n3450), .I2(n3451), .O(n3452));
  LUT3 #(.INIT(8'h96)) lut_n3453 (.I0(n3420), .I1(n3428), .I2(n3429), .O(n3453));
  LUT3 #(.INIT(8'hE8)) lut_n3454 (.I0(n3444), .I1(n3452), .I2(n3453), .O(n3454));
  LUT3 #(.INIT(8'hE8)) lut_n3455 (.I0(x1752), .I1(x1753), .I2(x1754), .O(n3455));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3456 (.I0(x1743), .I1(x1744), .I2(x1745), .I3(n3448), .I4(n3449), .O(n3456));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3457 (.I0(x1749), .I1(x1750), .I2(x1751), .I3(n3455), .I4(n3456), .O(n3457));
  LUT3 #(.INIT(8'hE8)) lut_n3458 (.I0(x1758), .I1(x1759), .I2(x1760), .O(n3458));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3459 (.I0(x1749), .I1(x1750), .I2(x1751), .I3(n3455), .I4(n3456), .O(n3459));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3460 (.I0(x1755), .I1(x1756), .I2(x1757), .I3(n3458), .I4(n3459), .O(n3460));
  LUT3 #(.INIT(8'h96)) lut_n3461 (.I0(n3447), .I1(n3450), .I2(n3451), .O(n3461));
  LUT3 #(.INIT(8'hE8)) lut_n3462 (.I0(n3457), .I1(n3460), .I2(n3461), .O(n3462));
  LUT3 #(.INIT(8'hE8)) lut_n3463 (.I0(x1764), .I1(x1765), .I2(x1766), .O(n3463));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3464 (.I0(x1755), .I1(x1756), .I2(x1757), .I3(n3458), .I4(n3459), .O(n3464));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3465 (.I0(x1761), .I1(x1762), .I2(x1763), .I3(n3463), .I4(n3464), .O(n3465));
  LUT3 #(.INIT(8'hE8)) lut_n3466 (.I0(x1770), .I1(x1771), .I2(x1772), .O(n3466));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3467 (.I0(x1761), .I1(x1762), .I2(x1763), .I3(n3463), .I4(n3464), .O(n3467));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3468 (.I0(x1767), .I1(x1768), .I2(x1769), .I3(n3466), .I4(n3467), .O(n3468));
  LUT3 #(.INIT(8'h96)) lut_n3469 (.I0(n3457), .I1(n3460), .I2(n3461), .O(n3469));
  LUT3 #(.INIT(8'hE8)) lut_n3470 (.I0(n3465), .I1(n3468), .I2(n3469), .O(n3470));
  LUT3 #(.INIT(8'h96)) lut_n3471 (.I0(n3444), .I1(n3452), .I2(n3453), .O(n3471));
  LUT3 #(.INIT(8'hE8)) lut_n3472 (.I0(n3462), .I1(n3470), .I2(n3471), .O(n3472));
  LUT3 #(.INIT(8'h96)) lut_n3473 (.I0(n3412), .I1(n3430), .I2(n3431), .O(n3473));
  LUT3 #(.INIT(8'hE8)) lut_n3474 (.I0(n3454), .I1(n3472), .I2(n3473), .O(n3474));
  LUT3 #(.INIT(8'hE8)) lut_n3475 (.I0(x1776), .I1(x1777), .I2(x1778), .O(n3475));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3476 (.I0(x1767), .I1(x1768), .I2(x1769), .I3(n3466), .I4(n3467), .O(n3476));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3477 (.I0(x1773), .I1(x1774), .I2(x1775), .I3(n3475), .I4(n3476), .O(n3477));
  LUT3 #(.INIT(8'hE8)) lut_n3478 (.I0(x1782), .I1(x1783), .I2(x1784), .O(n3478));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3479 (.I0(x1773), .I1(x1774), .I2(x1775), .I3(n3475), .I4(n3476), .O(n3479));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3480 (.I0(x1779), .I1(x1780), .I2(x1781), .I3(n3478), .I4(n3479), .O(n3480));
  LUT3 #(.INIT(8'h96)) lut_n3481 (.I0(n3465), .I1(n3468), .I2(n3469), .O(n3481));
  LUT3 #(.INIT(8'hE8)) lut_n3482 (.I0(n3477), .I1(n3480), .I2(n3481), .O(n3482));
  LUT3 #(.INIT(8'hE8)) lut_n3483 (.I0(x1788), .I1(x1789), .I2(x1790), .O(n3483));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3484 (.I0(x1779), .I1(x1780), .I2(x1781), .I3(n3478), .I4(n3479), .O(n3484));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3485 (.I0(x1785), .I1(x1786), .I2(x1787), .I3(n3483), .I4(n3484), .O(n3485));
  LUT3 #(.INIT(8'hE8)) lut_n3486 (.I0(x1794), .I1(x1795), .I2(x1796), .O(n3486));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3487 (.I0(x1785), .I1(x1786), .I2(x1787), .I3(n3483), .I4(n3484), .O(n3487));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3488 (.I0(x1791), .I1(x1792), .I2(x1793), .I3(n3486), .I4(n3487), .O(n3488));
  LUT3 #(.INIT(8'h96)) lut_n3489 (.I0(n3477), .I1(n3480), .I2(n3481), .O(n3489));
  LUT3 #(.INIT(8'hE8)) lut_n3490 (.I0(n3485), .I1(n3488), .I2(n3489), .O(n3490));
  LUT3 #(.INIT(8'h96)) lut_n3491 (.I0(n3462), .I1(n3470), .I2(n3471), .O(n3491));
  LUT3 #(.INIT(8'hE8)) lut_n3492 (.I0(n3482), .I1(n3490), .I2(n3491), .O(n3492));
  LUT3 #(.INIT(8'hE8)) lut_n3493 (.I0(x1800), .I1(x1801), .I2(x1802), .O(n3493));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3494 (.I0(x1791), .I1(x1792), .I2(x1793), .I3(n3486), .I4(n3487), .O(n3494));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3495 (.I0(x1797), .I1(x1798), .I2(x1799), .I3(n3493), .I4(n3494), .O(n3495));
  LUT3 #(.INIT(8'hE8)) lut_n3496 (.I0(x1806), .I1(x1807), .I2(x1808), .O(n3496));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3497 (.I0(x1797), .I1(x1798), .I2(x1799), .I3(n3493), .I4(n3494), .O(n3497));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3498 (.I0(x1803), .I1(x1804), .I2(x1805), .I3(n3496), .I4(n3497), .O(n3498));
  LUT3 #(.INIT(8'h96)) lut_n3499 (.I0(n3485), .I1(n3488), .I2(n3489), .O(n3499));
  LUT3 #(.INIT(8'hE8)) lut_n3500 (.I0(n3495), .I1(n3498), .I2(n3499), .O(n3500));
  LUT3 #(.INIT(8'hE8)) lut_n3501 (.I0(x1812), .I1(x1813), .I2(x1814), .O(n3501));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3502 (.I0(x1803), .I1(x1804), .I2(x1805), .I3(n3496), .I4(n3497), .O(n3502));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3503 (.I0(x1809), .I1(x1810), .I2(x1811), .I3(n3501), .I4(n3502), .O(n3503));
  LUT3 #(.INIT(8'hE8)) lut_n3504 (.I0(x1818), .I1(x1819), .I2(x1820), .O(n3504));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3505 (.I0(x1809), .I1(x1810), .I2(x1811), .I3(n3501), .I4(n3502), .O(n3505));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3506 (.I0(x1815), .I1(x1816), .I2(x1817), .I3(n3504), .I4(n3505), .O(n3506));
  LUT3 #(.INIT(8'h96)) lut_n3507 (.I0(n3495), .I1(n3498), .I2(n3499), .O(n3507));
  LUT3 #(.INIT(8'hE8)) lut_n3508 (.I0(n3503), .I1(n3506), .I2(n3507), .O(n3508));
  LUT3 #(.INIT(8'h96)) lut_n3509 (.I0(n3482), .I1(n3490), .I2(n3491), .O(n3509));
  LUT3 #(.INIT(8'hE8)) lut_n3510 (.I0(n3500), .I1(n3508), .I2(n3509), .O(n3510));
  LUT3 #(.INIT(8'h96)) lut_n3511 (.I0(n3454), .I1(n3472), .I2(n3473), .O(n3511));
  LUT3 #(.INIT(8'hE8)) lut_n3512 (.I0(n3492), .I1(n3510), .I2(n3511), .O(n3512));
  LUT3 #(.INIT(8'h96)) lut_n3513 (.I0(n3394), .I1(n3432), .I2(n3433), .O(n3513));
  LUT3 #(.INIT(8'hE8)) lut_n3514 (.I0(n3474), .I1(n3512), .I2(n3513), .O(n3514));
  LUT3 #(.INIT(8'hE8)) lut_n3515 (.I0(x1824), .I1(x1825), .I2(x1826), .O(n3515));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3516 (.I0(x1815), .I1(x1816), .I2(x1817), .I3(n3504), .I4(n3505), .O(n3516));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3517 (.I0(x1821), .I1(x1822), .I2(x1823), .I3(n3515), .I4(n3516), .O(n3517));
  LUT3 #(.INIT(8'hE8)) lut_n3518 (.I0(x1830), .I1(x1831), .I2(x1832), .O(n3518));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3519 (.I0(x1821), .I1(x1822), .I2(x1823), .I3(n3515), .I4(n3516), .O(n3519));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3520 (.I0(x1827), .I1(x1828), .I2(x1829), .I3(n3518), .I4(n3519), .O(n3520));
  LUT3 #(.INIT(8'h96)) lut_n3521 (.I0(n3503), .I1(n3506), .I2(n3507), .O(n3521));
  LUT3 #(.INIT(8'hE8)) lut_n3522 (.I0(n3517), .I1(n3520), .I2(n3521), .O(n3522));
  LUT3 #(.INIT(8'hE8)) lut_n3523 (.I0(x1836), .I1(x1837), .I2(x1838), .O(n3523));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3524 (.I0(x1827), .I1(x1828), .I2(x1829), .I3(n3518), .I4(n3519), .O(n3524));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3525 (.I0(x1833), .I1(x1834), .I2(x1835), .I3(n3523), .I4(n3524), .O(n3525));
  LUT3 #(.INIT(8'hE8)) lut_n3526 (.I0(x1842), .I1(x1843), .I2(x1844), .O(n3526));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3527 (.I0(x1833), .I1(x1834), .I2(x1835), .I3(n3523), .I4(n3524), .O(n3527));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3528 (.I0(x1839), .I1(x1840), .I2(x1841), .I3(n3526), .I4(n3527), .O(n3528));
  LUT3 #(.INIT(8'h96)) lut_n3529 (.I0(n3517), .I1(n3520), .I2(n3521), .O(n3529));
  LUT3 #(.INIT(8'hE8)) lut_n3530 (.I0(n3525), .I1(n3528), .I2(n3529), .O(n3530));
  LUT3 #(.INIT(8'h96)) lut_n3531 (.I0(n3500), .I1(n3508), .I2(n3509), .O(n3531));
  LUT3 #(.INIT(8'hE8)) lut_n3532 (.I0(n3522), .I1(n3530), .I2(n3531), .O(n3532));
  LUT3 #(.INIT(8'hE8)) lut_n3533 (.I0(x1848), .I1(x1849), .I2(x1850), .O(n3533));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3534 (.I0(x1839), .I1(x1840), .I2(x1841), .I3(n3526), .I4(n3527), .O(n3534));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3535 (.I0(x1845), .I1(x1846), .I2(x1847), .I3(n3533), .I4(n3534), .O(n3535));
  LUT3 #(.INIT(8'hE8)) lut_n3536 (.I0(x1854), .I1(x1855), .I2(x1856), .O(n3536));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3537 (.I0(x1845), .I1(x1846), .I2(x1847), .I3(n3533), .I4(n3534), .O(n3537));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3538 (.I0(x1851), .I1(x1852), .I2(x1853), .I3(n3536), .I4(n3537), .O(n3538));
  LUT3 #(.INIT(8'h96)) lut_n3539 (.I0(n3525), .I1(n3528), .I2(n3529), .O(n3539));
  LUT3 #(.INIT(8'hE8)) lut_n3540 (.I0(n3535), .I1(n3538), .I2(n3539), .O(n3540));
  LUT3 #(.INIT(8'hE8)) lut_n3541 (.I0(x1860), .I1(x1861), .I2(x1862), .O(n3541));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3542 (.I0(x1851), .I1(x1852), .I2(x1853), .I3(n3536), .I4(n3537), .O(n3542));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3543 (.I0(x1857), .I1(x1858), .I2(x1859), .I3(n3541), .I4(n3542), .O(n3543));
  LUT3 #(.INIT(8'hE8)) lut_n3544 (.I0(x1866), .I1(x1867), .I2(x1868), .O(n3544));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3545 (.I0(x1857), .I1(x1858), .I2(x1859), .I3(n3541), .I4(n3542), .O(n3545));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3546 (.I0(x1863), .I1(x1864), .I2(x1865), .I3(n3544), .I4(n3545), .O(n3546));
  LUT3 #(.INIT(8'h96)) lut_n3547 (.I0(n3535), .I1(n3538), .I2(n3539), .O(n3547));
  LUT3 #(.INIT(8'hE8)) lut_n3548 (.I0(n3543), .I1(n3546), .I2(n3547), .O(n3548));
  LUT3 #(.INIT(8'h96)) lut_n3549 (.I0(n3522), .I1(n3530), .I2(n3531), .O(n3549));
  LUT3 #(.INIT(8'hE8)) lut_n3550 (.I0(n3540), .I1(n3548), .I2(n3549), .O(n3550));
  LUT3 #(.INIT(8'h96)) lut_n3551 (.I0(n3492), .I1(n3510), .I2(n3511), .O(n3551));
  LUT3 #(.INIT(8'hE8)) lut_n3552 (.I0(n3532), .I1(n3550), .I2(n3551), .O(n3552));
  LUT3 #(.INIT(8'hE8)) lut_n3553 (.I0(x1872), .I1(x1873), .I2(x1874), .O(n3553));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3554 (.I0(x1863), .I1(x1864), .I2(x1865), .I3(n3544), .I4(n3545), .O(n3554));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3555 (.I0(x1869), .I1(x1870), .I2(x1871), .I3(n3553), .I4(n3554), .O(n3555));
  LUT3 #(.INIT(8'hE8)) lut_n3556 (.I0(x1878), .I1(x1879), .I2(x1880), .O(n3556));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3557 (.I0(x1869), .I1(x1870), .I2(x1871), .I3(n3553), .I4(n3554), .O(n3557));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3558 (.I0(x1875), .I1(x1876), .I2(x1877), .I3(n3556), .I4(n3557), .O(n3558));
  LUT3 #(.INIT(8'h96)) lut_n3559 (.I0(n3543), .I1(n3546), .I2(n3547), .O(n3559));
  LUT3 #(.INIT(8'hE8)) lut_n3560 (.I0(n3555), .I1(n3558), .I2(n3559), .O(n3560));
  LUT3 #(.INIT(8'hE8)) lut_n3561 (.I0(x1884), .I1(x1885), .I2(x1886), .O(n3561));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3562 (.I0(x1875), .I1(x1876), .I2(x1877), .I3(n3556), .I4(n3557), .O(n3562));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3563 (.I0(x1881), .I1(x1882), .I2(x1883), .I3(n3561), .I4(n3562), .O(n3563));
  LUT3 #(.INIT(8'hE8)) lut_n3564 (.I0(x1890), .I1(x1891), .I2(x1892), .O(n3564));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3565 (.I0(x1881), .I1(x1882), .I2(x1883), .I3(n3561), .I4(n3562), .O(n3565));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3566 (.I0(x1887), .I1(x1888), .I2(x1889), .I3(n3564), .I4(n3565), .O(n3566));
  LUT3 #(.INIT(8'h96)) lut_n3567 (.I0(n3555), .I1(n3558), .I2(n3559), .O(n3567));
  LUT3 #(.INIT(8'hE8)) lut_n3568 (.I0(n3563), .I1(n3566), .I2(n3567), .O(n3568));
  LUT3 #(.INIT(8'h96)) lut_n3569 (.I0(n3540), .I1(n3548), .I2(n3549), .O(n3569));
  LUT3 #(.INIT(8'hE8)) lut_n3570 (.I0(n3560), .I1(n3568), .I2(n3569), .O(n3570));
  LUT3 #(.INIT(8'hE8)) lut_n3571 (.I0(x1896), .I1(x1897), .I2(x1898), .O(n3571));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3572 (.I0(x1887), .I1(x1888), .I2(x1889), .I3(n3564), .I4(n3565), .O(n3572));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3573 (.I0(x1893), .I1(x1894), .I2(x1895), .I3(n3571), .I4(n3572), .O(n3573));
  LUT3 #(.INIT(8'hE8)) lut_n3574 (.I0(x1902), .I1(x1903), .I2(x1904), .O(n3574));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3575 (.I0(x1893), .I1(x1894), .I2(x1895), .I3(n3571), .I4(n3572), .O(n3575));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3576 (.I0(x1899), .I1(x1900), .I2(x1901), .I3(n3574), .I4(n3575), .O(n3576));
  LUT3 #(.INIT(8'h96)) lut_n3577 (.I0(n3563), .I1(n3566), .I2(n3567), .O(n3577));
  LUT3 #(.INIT(8'hE8)) lut_n3578 (.I0(n3573), .I1(n3576), .I2(n3577), .O(n3578));
  LUT3 #(.INIT(8'hE8)) lut_n3579 (.I0(x1908), .I1(x1909), .I2(x1910), .O(n3579));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3580 (.I0(x1899), .I1(x1900), .I2(x1901), .I3(n3574), .I4(n3575), .O(n3580));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3581 (.I0(x1905), .I1(x1906), .I2(x1907), .I3(n3579), .I4(n3580), .O(n3581));
  LUT3 #(.INIT(8'hE8)) lut_n3582 (.I0(x1914), .I1(x1915), .I2(x1916), .O(n3582));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3583 (.I0(x1905), .I1(x1906), .I2(x1907), .I3(n3579), .I4(n3580), .O(n3583));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3584 (.I0(x1911), .I1(x1912), .I2(x1913), .I3(n3582), .I4(n3583), .O(n3584));
  LUT3 #(.INIT(8'h96)) lut_n3585 (.I0(n3573), .I1(n3576), .I2(n3577), .O(n3585));
  LUT3 #(.INIT(8'hE8)) lut_n3586 (.I0(n3581), .I1(n3584), .I2(n3585), .O(n3586));
  LUT3 #(.INIT(8'h96)) lut_n3587 (.I0(n3560), .I1(n3568), .I2(n3569), .O(n3587));
  LUT3 #(.INIT(8'hE8)) lut_n3588 (.I0(n3578), .I1(n3586), .I2(n3587), .O(n3588));
  LUT3 #(.INIT(8'h96)) lut_n3589 (.I0(n3532), .I1(n3550), .I2(n3551), .O(n3589));
  LUT3 #(.INIT(8'hE8)) lut_n3590 (.I0(n3570), .I1(n3588), .I2(n3589), .O(n3590));
  LUT3 #(.INIT(8'h96)) lut_n3591 (.I0(n3474), .I1(n3512), .I2(n3513), .O(n3591));
  LUT3 #(.INIT(8'hE8)) lut_n3592 (.I0(n3552), .I1(n3590), .I2(n3591), .O(n3592));
  LUT3 #(.INIT(8'h96)) lut_n3593 (.I0(n3356), .I1(n3434), .I2(n3435), .O(n3593));
  LUT3 #(.INIT(8'hE8)) lut_n3594 (.I0(n3514), .I1(n3592), .I2(n3593), .O(n3594));
  LUT3 #(.INIT(8'h96)) lut_n3595 (.I0(n3117), .I1(n3275), .I2(n3276), .O(n3595));
  LUT3 #(.INIT(8'hE8)) lut_n3596 (.I0(n3436), .I1(n3594), .I2(n3595), .O(n3596));
  LUT3 #(.INIT(8'hE8)) lut_n3597 (.I0(x1920), .I1(x1921), .I2(x1922), .O(n3597));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3598 (.I0(x1911), .I1(x1912), .I2(x1913), .I3(n3582), .I4(n3583), .O(n3598));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3599 (.I0(x1917), .I1(x1918), .I2(x1919), .I3(n3597), .I4(n3598), .O(n3599));
  LUT3 #(.INIT(8'hE8)) lut_n3600 (.I0(x1926), .I1(x1927), .I2(x1928), .O(n3600));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3601 (.I0(x1917), .I1(x1918), .I2(x1919), .I3(n3597), .I4(n3598), .O(n3601));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3602 (.I0(x1923), .I1(x1924), .I2(x1925), .I3(n3600), .I4(n3601), .O(n3602));
  LUT3 #(.INIT(8'h96)) lut_n3603 (.I0(n3581), .I1(n3584), .I2(n3585), .O(n3603));
  LUT3 #(.INIT(8'hE8)) lut_n3604 (.I0(n3599), .I1(n3602), .I2(n3603), .O(n3604));
  LUT3 #(.INIT(8'hE8)) lut_n3605 (.I0(x1932), .I1(x1933), .I2(x1934), .O(n3605));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3606 (.I0(x1923), .I1(x1924), .I2(x1925), .I3(n3600), .I4(n3601), .O(n3606));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3607 (.I0(x1929), .I1(x1930), .I2(x1931), .I3(n3605), .I4(n3606), .O(n3607));
  LUT3 #(.INIT(8'hE8)) lut_n3608 (.I0(x1938), .I1(x1939), .I2(x1940), .O(n3608));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3609 (.I0(x1929), .I1(x1930), .I2(x1931), .I3(n3605), .I4(n3606), .O(n3609));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3610 (.I0(x1935), .I1(x1936), .I2(x1937), .I3(n3608), .I4(n3609), .O(n3610));
  LUT3 #(.INIT(8'h96)) lut_n3611 (.I0(n3599), .I1(n3602), .I2(n3603), .O(n3611));
  LUT3 #(.INIT(8'hE8)) lut_n3612 (.I0(n3607), .I1(n3610), .I2(n3611), .O(n3612));
  LUT3 #(.INIT(8'h96)) lut_n3613 (.I0(n3578), .I1(n3586), .I2(n3587), .O(n3613));
  LUT3 #(.INIT(8'hE8)) lut_n3614 (.I0(n3604), .I1(n3612), .I2(n3613), .O(n3614));
  LUT3 #(.INIT(8'hE8)) lut_n3615 (.I0(x1944), .I1(x1945), .I2(x1946), .O(n3615));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3616 (.I0(x1935), .I1(x1936), .I2(x1937), .I3(n3608), .I4(n3609), .O(n3616));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3617 (.I0(x1941), .I1(x1942), .I2(x1943), .I3(n3615), .I4(n3616), .O(n3617));
  LUT3 #(.INIT(8'hE8)) lut_n3618 (.I0(x1950), .I1(x1951), .I2(x1952), .O(n3618));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3619 (.I0(x1941), .I1(x1942), .I2(x1943), .I3(n3615), .I4(n3616), .O(n3619));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3620 (.I0(x1947), .I1(x1948), .I2(x1949), .I3(n3618), .I4(n3619), .O(n3620));
  LUT3 #(.INIT(8'h96)) lut_n3621 (.I0(n3607), .I1(n3610), .I2(n3611), .O(n3621));
  LUT3 #(.INIT(8'hE8)) lut_n3622 (.I0(n3617), .I1(n3620), .I2(n3621), .O(n3622));
  LUT3 #(.INIT(8'hE8)) lut_n3623 (.I0(x1956), .I1(x1957), .I2(x1958), .O(n3623));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3624 (.I0(x1947), .I1(x1948), .I2(x1949), .I3(n3618), .I4(n3619), .O(n3624));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3625 (.I0(x1953), .I1(x1954), .I2(x1955), .I3(n3623), .I4(n3624), .O(n3625));
  LUT3 #(.INIT(8'hE8)) lut_n3626 (.I0(x1962), .I1(x1963), .I2(x1964), .O(n3626));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3627 (.I0(x1953), .I1(x1954), .I2(x1955), .I3(n3623), .I4(n3624), .O(n3627));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3628 (.I0(x1959), .I1(x1960), .I2(x1961), .I3(n3626), .I4(n3627), .O(n3628));
  LUT3 #(.INIT(8'h96)) lut_n3629 (.I0(n3617), .I1(n3620), .I2(n3621), .O(n3629));
  LUT3 #(.INIT(8'hE8)) lut_n3630 (.I0(n3625), .I1(n3628), .I2(n3629), .O(n3630));
  LUT3 #(.INIT(8'h96)) lut_n3631 (.I0(n3604), .I1(n3612), .I2(n3613), .O(n3631));
  LUT3 #(.INIT(8'hE8)) lut_n3632 (.I0(n3622), .I1(n3630), .I2(n3631), .O(n3632));
  LUT3 #(.INIT(8'h96)) lut_n3633 (.I0(n3570), .I1(n3588), .I2(n3589), .O(n3633));
  LUT3 #(.INIT(8'hE8)) lut_n3634 (.I0(n3614), .I1(n3632), .I2(n3633), .O(n3634));
  LUT3 #(.INIT(8'hE8)) lut_n3635 (.I0(x1968), .I1(x1969), .I2(x1970), .O(n3635));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3636 (.I0(x1959), .I1(x1960), .I2(x1961), .I3(n3626), .I4(n3627), .O(n3636));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3637 (.I0(x1965), .I1(x1966), .I2(x1967), .I3(n3635), .I4(n3636), .O(n3637));
  LUT3 #(.INIT(8'hE8)) lut_n3638 (.I0(x1974), .I1(x1975), .I2(x1976), .O(n3638));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3639 (.I0(x1965), .I1(x1966), .I2(x1967), .I3(n3635), .I4(n3636), .O(n3639));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3640 (.I0(x1971), .I1(x1972), .I2(x1973), .I3(n3638), .I4(n3639), .O(n3640));
  LUT3 #(.INIT(8'h96)) lut_n3641 (.I0(n3625), .I1(n3628), .I2(n3629), .O(n3641));
  LUT3 #(.INIT(8'hE8)) lut_n3642 (.I0(n3637), .I1(n3640), .I2(n3641), .O(n3642));
  LUT3 #(.INIT(8'hE8)) lut_n3643 (.I0(x1980), .I1(x1981), .I2(x1982), .O(n3643));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3644 (.I0(x1971), .I1(x1972), .I2(x1973), .I3(n3638), .I4(n3639), .O(n3644));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3645 (.I0(x1977), .I1(x1978), .I2(x1979), .I3(n3643), .I4(n3644), .O(n3645));
  LUT3 #(.INIT(8'hE8)) lut_n3646 (.I0(x1986), .I1(x1987), .I2(x1988), .O(n3646));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3647 (.I0(x1977), .I1(x1978), .I2(x1979), .I3(n3643), .I4(n3644), .O(n3647));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3648 (.I0(x1983), .I1(x1984), .I2(x1985), .I3(n3646), .I4(n3647), .O(n3648));
  LUT3 #(.INIT(8'h96)) lut_n3649 (.I0(n3637), .I1(n3640), .I2(n3641), .O(n3649));
  LUT3 #(.INIT(8'hE8)) lut_n3650 (.I0(n3645), .I1(n3648), .I2(n3649), .O(n3650));
  LUT3 #(.INIT(8'h96)) lut_n3651 (.I0(n3622), .I1(n3630), .I2(n3631), .O(n3651));
  LUT3 #(.INIT(8'hE8)) lut_n3652 (.I0(n3642), .I1(n3650), .I2(n3651), .O(n3652));
  LUT3 #(.INIT(8'hE8)) lut_n3653 (.I0(x1992), .I1(x1993), .I2(x1994), .O(n3653));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3654 (.I0(x1983), .I1(x1984), .I2(x1985), .I3(n3646), .I4(n3647), .O(n3654));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3655 (.I0(x1989), .I1(x1990), .I2(x1991), .I3(n3653), .I4(n3654), .O(n3655));
  LUT3 #(.INIT(8'hE8)) lut_n3656 (.I0(x1998), .I1(x1999), .I2(x2000), .O(n3656));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3657 (.I0(x1989), .I1(x1990), .I2(x1991), .I3(n3653), .I4(n3654), .O(n3657));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3658 (.I0(x1995), .I1(x1996), .I2(x1997), .I3(n3656), .I4(n3657), .O(n3658));
  LUT3 #(.INIT(8'h96)) lut_n3659 (.I0(n3645), .I1(n3648), .I2(n3649), .O(n3659));
  LUT3 #(.INIT(8'hE8)) lut_n3660 (.I0(n3655), .I1(n3658), .I2(n3659), .O(n3660));
  LUT3 #(.INIT(8'hE8)) lut_n3661 (.I0(x2004), .I1(x2005), .I2(x2006), .O(n3661));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3662 (.I0(x1995), .I1(x1996), .I2(x1997), .I3(n3656), .I4(n3657), .O(n3662));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3663 (.I0(x2001), .I1(x2002), .I2(x2003), .I3(n3661), .I4(n3662), .O(n3663));
  LUT3 #(.INIT(8'hE8)) lut_n3664 (.I0(x2010), .I1(x2011), .I2(x2012), .O(n3664));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3665 (.I0(x2001), .I1(x2002), .I2(x2003), .I3(n3661), .I4(n3662), .O(n3665));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3666 (.I0(x2007), .I1(x2008), .I2(x2009), .I3(n3664), .I4(n3665), .O(n3666));
  LUT3 #(.INIT(8'h96)) lut_n3667 (.I0(n3655), .I1(n3658), .I2(n3659), .O(n3667));
  LUT3 #(.INIT(8'hE8)) lut_n3668 (.I0(n3663), .I1(n3666), .I2(n3667), .O(n3668));
  LUT3 #(.INIT(8'h96)) lut_n3669 (.I0(n3642), .I1(n3650), .I2(n3651), .O(n3669));
  LUT3 #(.INIT(8'hE8)) lut_n3670 (.I0(n3660), .I1(n3668), .I2(n3669), .O(n3670));
  LUT3 #(.INIT(8'h96)) lut_n3671 (.I0(n3614), .I1(n3632), .I2(n3633), .O(n3671));
  LUT3 #(.INIT(8'hE8)) lut_n3672 (.I0(n3652), .I1(n3670), .I2(n3671), .O(n3672));
  LUT3 #(.INIT(8'h96)) lut_n3673 (.I0(n3552), .I1(n3590), .I2(n3591), .O(n3673));
  LUT3 #(.INIT(8'hE8)) lut_n3674 (.I0(n3634), .I1(n3672), .I2(n3673), .O(n3674));
  LUT3 #(.INIT(8'hE8)) lut_n3675 (.I0(x2016), .I1(x2017), .I2(x2018), .O(n3675));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3676 (.I0(x2007), .I1(x2008), .I2(x2009), .I3(n3664), .I4(n3665), .O(n3676));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3677 (.I0(x2013), .I1(x2014), .I2(x2015), .I3(n3675), .I4(n3676), .O(n3677));
  LUT3 #(.INIT(8'hE8)) lut_n3678 (.I0(x2022), .I1(x2023), .I2(x2024), .O(n3678));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3679 (.I0(x2013), .I1(x2014), .I2(x2015), .I3(n3675), .I4(n3676), .O(n3679));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n3680 (.I0(x2019), .I1(x2020), .I2(x2021), .I3(n3678), .I4(n3679), .O(n3680));
  LUT3 #(.INIT(8'h96)) lut_n3681 (.I0(n3663), .I1(n3666), .I2(n3667), .O(n3681));
  LUT3 #(.INIT(8'hE8)) lut_n3682 (.I0(n3677), .I1(n3680), .I2(n3681), .O(n3682));
  LUT3 #(.INIT(8'h96)) lut_n3683 (.I0(x0), .I1(x1), .I2(x2), .O(n3683));
  LUT3 #(.INIT(8'h96)) lut_n3684 (.I0(x6), .I1(x7), .I2(x8), .O(n3684));
  LUT5 #(.INIT(32'hFF969600)) lut_n3685 (.I0(x3), .I1(x4), .I2(x5), .I3(n3683), .I4(n3684), .O(n3685));
  LUT3 #(.INIT(8'h96)) lut_n3686 (.I0(x12), .I1(x13), .I2(x14), .O(n3686));
  LUT5 #(.INIT(32'h96696996)) lut_n3687 (.I0(x3), .I1(x4), .I2(x5), .I3(n3683), .I4(n3684), .O(n3687));
  LUT5 #(.INIT(32'hFF969600)) lut_n3688 (.I0(x9), .I1(x10), .I2(x11), .I3(n3686), .I4(n3687), .O(n3688));
  LUT5 #(.INIT(32'hE81717E8)) lut_n3689 (.I0(x2019), .I1(x2020), .I2(x2021), .I3(n3678), .I4(n3679), .O(n3689));
  LUT3 #(.INIT(8'hE8)) lut_n3690 (.I0(n3685), .I1(n3688), .I2(n3689), .O(n3690));
  LUT3 #(.INIT(8'h96)) lut_n3691 (.I0(x18), .I1(x19), .I2(x20), .O(n3691));
  LUT5 #(.INIT(32'h96696996)) lut_n3692 (.I0(x9), .I1(x10), .I2(x11), .I3(n3686), .I4(n3687), .O(n3692));
  LUT5 #(.INIT(32'hFF969600)) lut_n3693 (.I0(x15), .I1(x16), .I2(x17), .I3(n3691), .I4(n3692), .O(n3693));
  LUT3 #(.INIT(8'h96)) lut_n3694 (.I0(x24), .I1(x25), .I2(x26), .O(n3694));
  LUT5 #(.INIT(32'h96696996)) lut_n3695 (.I0(x15), .I1(x16), .I2(x17), .I3(n3691), .I4(n3692), .O(n3695));
  LUT5 #(.INIT(32'hFF969600)) lut_n3696 (.I0(x21), .I1(x22), .I2(x23), .I3(n3694), .I4(n3695), .O(n3696));
  LUT3 #(.INIT(8'h96)) lut_n3697 (.I0(n3685), .I1(n3688), .I2(n3689), .O(n3697));
  LUT3 #(.INIT(8'hE8)) lut_n3698 (.I0(n3693), .I1(n3696), .I2(n3697), .O(n3698));
  LUT3 #(.INIT(8'h96)) lut_n3699 (.I0(n3677), .I1(n3680), .I2(n3681), .O(n3699));
  LUT3 #(.INIT(8'hE8)) lut_n3700 (.I0(n3690), .I1(n3698), .I2(n3699), .O(n3700));
  LUT3 #(.INIT(8'h96)) lut_n3701 (.I0(n3660), .I1(n3668), .I2(n3669), .O(n3701));
  LUT3 #(.INIT(8'hE8)) lut_n3702 (.I0(n3682), .I1(n3700), .I2(n3701), .O(n3702));
  LUT3 #(.INIT(8'h96)) lut_n3703 (.I0(x27), .I1(x28), .I2(x29), .O(n3703));
  LUT5 #(.INIT(32'h96696996)) lut_n3704 (.I0(x21), .I1(x22), .I2(x23), .I3(n3694), .I4(n3695), .O(n3704));
  LUT5 #(.INIT(32'hFF969600)) lut_n3705 (.I0(x30), .I1(x31), .I2(x32), .I3(n3703), .I4(n3704), .O(n3705));
  LUT3 #(.INIT(8'h96)) lut_n3706 (.I0(x36), .I1(x37), .I2(x38), .O(n3706));
  LUT5 #(.INIT(32'h96696996)) lut_n3707 (.I0(x30), .I1(x31), .I2(x32), .I3(n3703), .I4(n3704), .O(n3707));
  LUT5 #(.INIT(32'hFF969600)) lut_n3708 (.I0(x33), .I1(x34), .I2(x35), .I3(n3706), .I4(n3707), .O(n3708));
  LUT3 #(.INIT(8'h96)) lut_n3709 (.I0(n3693), .I1(n3696), .I2(n3697), .O(n3709));
  LUT3 #(.INIT(8'hE8)) lut_n3710 (.I0(n3705), .I1(n3708), .I2(n3709), .O(n3710));
  LUT3 #(.INIT(8'h96)) lut_n3711 (.I0(x42), .I1(x43), .I2(x44), .O(n3711));
  LUT5 #(.INIT(32'h96696996)) lut_n3712 (.I0(x33), .I1(x34), .I2(x35), .I3(n3706), .I4(n3707), .O(n3712));
  LUT5 #(.INIT(32'hFF969600)) lut_n3713 (.I0(x39), .I1(x40), .I2(x41), .I3(n3711), .I4(n3712), .O(n3713));
  LUT3 #(.INIT(8'h96)) lut_n3714 (.I0(x48), .I1(x49), .I2(x50), .O(n3714));
  LUT5 #(.INIT(32'h96696996)) lut_n3715 (.I0(x39), .I1(x40), .I2(x41), .I3(n3711), .I4(n3712), .O(n3715));
  LUT5 #(.INIT(32'hFF969600)) lut_n3716 (.I0(x45), .I1(x46), .I2(x47), .I3(n3714), .I4(n3715), .O(n3716));
  LUT3 #(.INIT(8'h96)) lut_n3717 (.I0(n3705), .I1(n3708), .I2(n3709), .O(n3717));
  LUT3 #(.INIT(8'hE8)) lut_n3718 (.I0(n3713), .I1(n3716), .I2(n3717), .O(n3718));
  LUT3 #(.INIT(8'h96)) lut_n3719 (.I0(n3690), .I1(n3698), .I2(n3699), .O(n3719));
  LUT3 #(.INIT(8'hE8)) lut_n3720 (.I0(n3710), .I1(n3718), .I2(n3719), .O(n3720));
  LUT3 #(.INIT(8'h96)) lut_n3721 (.I0(x54), .I1(x55), .I2(x56), .O(n3721));
  LUT5 #(.INIT(32'h96696996)) lut_n3722 (.I0(x45), .I1(x46), .I2(x47), .I3(n3714), .I4(n3715), .O(n3722));
  LUT5 #(.INIT(32'hFF969600)) lut_n3723 (.I0(x51), .I1(x52), .I2(x53), .I3(n3721), .I4(n3722), .O(n3723));
  LUT3 #(.INIT(8'h96)) lut_n3724 (.I0(x60), .I1(x61), .I2(x62), .O(n3724));
  LUT5 #(.INIT(32'h96696996)) lut_n3725 (.I0(x51), .I1(x52), .I2(x53), .I3(n3721), .I4(n3722), .O(n3725));
  LUT5 #(.INIT(32'hFF969600)) lut_n3726 (.I0(x57), .I1(x58), .I2(x59), .I3(n3724), .I4(n3725), .O(n3726));
  LUT3 #(.INIT(8'h96)) lut_n3727 (.I0(n3713), .I1(n3716), .I2(n3717), .O(n3727));
  LUT3 #(.INIT(8'hE8)) lut_n3728 (.I0(n3723), .I1(n3726), .I2(n3727), .O(n3728));
  LUT3 #(.INIT(8'h96)) lut_n3729 (.I0(x66), .I1(x67), .I2(x68), .O(n3729));
  LUT5 #(.INIT(32'h96696996)) lut_n3730 (.I0(x57), .I1(x58), .I2(x59), .I3(n3724), .I4(n3725), .O(n3730));
  LUT5 #(.INIT(32'hFF969600)) lut_n3731 (.I0(x63), .I1(x64), .I2(x65), .I3(n3729), .I4(n3730), .O(n3731));
  LUT3 #(.INIT(8'h96)) lut_n3732 (.I0(x72), .I1(x73), .I2(x74), .O(n3732));
  LUT5 #(.INIT(32'h96696996)) lut_n3733 (.I0(x63), .I1(x64), .I2(x65), .I3(n3729), .I4(n3730), .O(n3733));
  LUT5 #(.INIT(32'hFF969600)) lut_n3734 (.I0(x69), .I1(x70), .I2(x71), .I3(n3732), .I4(n3733), .O(n3734));
  LUT3 #(.INIT(8'h96)) lut_n3735 (.I0(n3723), .I1(n3726), .I2(n3727), .O(n3735));
  LUT3 #(.INIT(8'hE8)) lut_n3736 (.I0(n3731), .I1(n3734), .I2(n3735), .O(n3736));
  LUT3 #(.INIT(8'h96)) lut_n3737 (.I0(n3710), .I1(n3718), .I2(n3719), .O(n3737));
  LUT3 #(.INIT(8'hE8)) lut_n3738 (.I0(n3728), .I1(n3736), .I2(n3737), .O(n3738));
  LUT3 #(.INIT(8'h96)) lut_n3739 (.I0(n3682), .I1(n3700), .I2(n3701), .O(n3739));
  LUT3 #(.INIT(8'hE8)) lut_n3740 (.I0(n3720), .I1(n3738), .I2(n3739), .O(n3740));
  LUT3 #(.INIT(8'h96)) lut_n3741 (.I0(n3652), .I1(n3670), .I2(n3671), .O(n3741));
  LUT3 #(.INIT(8'hE8)) lut_n3742 (.I0(n3702), .I1(n3740), .I2(n3741), .O(n3742));
  LUT3 #(.INIT(8'h96)) lut_n3743 (.I0(x78), .I1(x79), .I2(x80), .O(n3743));
  LUT5 #(.INIT(32'h96696996)) lut_n3744 (.I0(x69), .I1(x70), .I2(x71), .I3(n3732), .I4(n3733), .O(n3744));
  LUT5 #(.INIT(32'hFF969600)) lut_n3745 (.I0(x75), .I1(x76), .I2(x77), .I3(n3743), .I4(n3744), .O(n3745));
  LUT3 #(.INIT(8'h96)) lut_n3746 (.I0(x84), .I1(x85), .I2(x86), .O(n3746));
  LUT5 #(.INIT(32'h96696996)) lut_n3747 (.I0(x75), .I1(x76), .I2(x77), .I3(n3743), .I4(n3744), .O(n3747));
  LUT5 #(.INIT(32'hFF969600)) lut_n3748 (.I0(x81), .I1(x82), .I2(x83), .I3(n3746), .I4(n3747), .O(n3748));
  LUT3 #(.INIT(8'h96)) lut_n3749 (.I0(n3731), .I1(n3734), .I2(n3735), .O(n3749));
  LUT3 #(.INIT(8'hE8)) lut_n3750 (.I0(n3745), .I1(n3748), .I2(n3749), .O(n3750));
  LUT3 #(.INIT(8'h96)) lut_n3751 (.I0(x90), .I1(x91), .I2(x92), .O(n3751));
  LUT5 #(.INIT(32'h96696996)) lut_n3752 (.I0(x81), .I1(x82), .I2(x83), .I3(n3746), .I4(n3747), .O(n3752));
  LUT5 #(.INIT(32'hFF969600)) lut_n3753 (.I0(x87), .I1(x88), .I2(x89), .I3(n3751), .I4(n3752), .O(n3753));
  LUT3 #(.INIT(8'h96)) lut_n3754 (.I0(x96), .I1(x97), .I2(x98), .O(n3754));
  LUT5 #(.INIT(32'h96696996)) lut_n3755 (.I0(x87), .I1(x88), .I2(x89), .I3(n3751), .I4(n3752), .O(n3755));
  LUT5 #(.INIT(32'hFF969600)) lut_n3756 (.I0(x93), .I1(x94), .I2(x95), .I3(n3754), .I4(n3755), .O(n3756));
  LUT3 #(.INIT(8'h96)) lut_n3757 (.I0(n3745), .I1(n3748), .I2(n3749), .O(n3757));
  LUT3 #(.INIT(8'hE8)) lut_n3758 (.I0(n3753), .I1(n3756), .I2(n3757), .O(n3758));
  LUT3 #(.INIT(8'h96)) lut_n3759 (.I0(n3728), .I1(n3736), .I2(n3737), .O(n3759));
  LUT3 #(.INIT(8'hE8)) lut_n3760 (.I0(n3750), .I1(n3758), .I2(n3759), .O(n3760));
  LUT3 #(.INIT(8'h96)) lut_n3761 (.I0(x102), .I1(x103), .I2(x104), .O(n3761));
  LUT5 #(.INIT(32'h96696996)) lut_n3762 (.I0(x93), .I1(x94), .I2(x95), .I3(n3754), .I4(n3755), .O(n3762));
  LUT5 #(.INIT(32'hFF969600)) lut_n3763 (.I0(x99), .I1(x100), .I2(x101), .I3(n3761), .I4(n3762), .O(n3763));
  LUT3 #(.INIT(8'h96)) lut_n3764 (.I0(x108), .I1(x109), .I2(x110), .O(n3764));
  LUT5 #(.INIT(32'h96696996)) lut_n3765 (.I0(x99), .I1(x100), .I2(x101), .I3(n3761), .I4(n3762), .O(n3765));
  LUT5 #(.INIT(32'hFF969600)) lut_n3766 (.I0(x105), .I1(x106), .I2(x107), .I3(n3764), .I4(n3765), .O(n3766));
  LUT3 #(.INIT(8'h96)) lut_n3767 (.I0(n3753), .I1(n3756), .I2(n3757), .O(n3767));
  LUT3 #(.INIT(8'hE8)) lut_n3768 (.I0(n3763), .I1(n3766), .I2(n3767), .O(n3768));
  LUT3 #(.INIT(8'h96)) lut_n3769 (.I0(x114), .I1(x115), .I2(x116), .O(n3769));
  LUT5 #(.INIT(32'h96696996)) lut_n3770 (.I0(x105), .I1(x106), .I2(x107), .I3(n3764), .I4(n3765), .O(n3770));
  LUT5 #(.INIT(32'hFF969600)) lut_n3771 (.I0(x111), .I1(x112), .I2(x113), .I3(n3769), .I4(n3770), .O(n3771));
  LUT3 #(.INIT(8'h96)) lut_n3772 (.I0(x120), .I1(x121), .I2(x122), .O(n3772));
  LUT5 #(.INIT(32'h96696996)) lut_n3773 (.I0(x111), .I1(x112), .I2(x113), .I3(n3769), .I4(n3770), .O(n3773));
  LUT5 #(.INIT(32'hFF969600)) lut_n3774 (.I0(x117), .I1(x118), .I2(x119), .I3(n3772), .I4(n3773), .O(n3774));
  LUT3 #(.INIT(8'h96)) lut_n3775 (.I0(n3763), .I1(n3766), .I2(n3767), .O(n3775));
  LUT3 #(.INIT(8'hE8)) lut_n3776 (.I0(n3771), .I1(n3774), .I2(n3775), .O(n3776));
  LUT3 #(.INIT(8'h96)) lut_n3777 (.I0(n3750), .I1(n3758), .I2(n3759), .O(n3777));
  LUT3 #(.INIT(8'hE8)) lut_n3778 (.I0(n3768), .I1(n3776), .I2(n3777), .O(n3778));
  LUT3 #(.INIT(8'h96)) lut_n3779 (.I0(n3720), .I1(n3738), .I2(n3739), .O(n3779));
  LUT3 #(.INIT(8'hE8)) lut_n3780 (.I0(n3760), .I1(n3778), .I2(n3779), .O(n3780));
  LUT3 #(.INIT(8'h96)) lut_n3781 (.I0(x126), .I1(x127), .I2(x128), .O(n3781));
  LUT5 #(.INIT(32'h96696996)) lut_n3782 (.I0(x117), .I1(x118), .I2(x119), .I3(n3772), .I4(n3773), .O(n3782));
  LUT5 #(.INIT(32'hFF969600)) lut_n3783 (.I0(x123), .I1(x124), .I2(x125), .I3(n3781), .I4(n3782), .O(n3783));
  LUT3 #(.INIT(8'h96)) lut_n3784 (.I0(x132), .I1(x133), .I2(x134), .O(n3784));
  LUT5 #(.INIT(32'h96696996)) lut_n3785 (.I0(x123), .I1(x124), .I2(x125), .I3(n3781), .I4(n3782), .O(n3785));
  LUT5 #(.INIT(32'hFF969600)) lut_n3786 (.I0(x129), .I1(x130), .I2(x131), .I3(n3784), .I4(n3785), .O(n3786));
  LUT3 #(.INIT(8'h96)) lut_n3787 (.I0(n3771), .I1(n3774), .I2(n3775), .O(n3787));
  LUT3 #(.INIT(8'hE8)) lut_n3788 (.I0(n3783), .I1(n3786), .I2(n3787), .O(n3788));
  LUT3 #(.INIT(8'h96)) lut_n3789 (.I0(x138), .I1(x139), .I2(x140), .O(n3789));
  LUT5 #(.INIT(32'h96696996)) lut_n3790 (.I0(x129), .I1(x130), .I2(x131), .I3(n3784), .I4(n3785), .O(n3790));
  LUT5 #(.INIT(32'hFF969600)) lut_n3791 (.I0(x135), .I1(x136), .I2(x137), .I3(n3789), .I4(n3790), .O(n3791));
  LUT3 #(.INIT(8'h96)) lut_n3792 (.I0(x144), .I1(x145), .I2(x146), .O(n3792));
  LUT5 #(.INIT(32'h96696996)) lut_n3793 (.I0(x135), .I1(x136), .I2(x137), .I3(n3789), .I4(n3790), .O(n3793));
  LUT5 #(.INIT(32'hFF969600)) lut_n3794 (.I0(x141), .I1(x142), .I2(x143), .I3(n3792), .I4(n3793), .O(n3794));
  LUT3 #(.INIT(8'h96)) lut_n3795 (.I0(n3783), .I1(n3786), .I2(n3787), .O(n3795));
  LUT3 #(.INIT(8'hE8)) lut_n3796 (.I0(n3791), .I1(n3794), .I2(n3795), .O(n3796));
  LUT3 #(.INIT(8'h96)) lut_n3797 (.I0(n3768), .I1(n3776), .I2(n3777), .O(n3797));
  LUT3 #(.INIT(8'hE8)) lut_n3798 (.I0(n3788), .I1(n3796), .I2(n3797), .O(n3798));
  LUT3 #(.INIT(8'h96)) lut_n3799 (.I0(x150), .I1(x151), .I2(x152), .O(n3799));
  LUT5 #(.INIT(32'h96696996)) lut_n3800 (.I0(x141), .I1(x142), .I2(x143), .I3(n3792), .I4(n3793), .O(n3800));
  LUT5 #(.INIT(32'hFF969600)) lut_n3801 (.I0(x147), .I1(x148), .I2(x149), .I3(n3799), .I4(n3800), .O(n3801));
  LUT3 #(.INIT(8'h96)) lut_n3802 (.I0(x156), .I1(x157), .I2(x158), .O(n3802));
  LUT5 #(.INIT(32'h96696996)) lut_n3803 (.I0(x147), .I1(x148), .I2(x149), .I3(n3799), .I4(n3800), .O(n3803));
  LUT5 #(.INIT(32'hFF969600)) lut_n3804 (.I0(x153), .I1(x154), .I2(x155), .I3(n3802), .I4(n3803), .O(n3804));
  LUT3 #(.INIT(8'h96)) lut_n3805 (.I0(n3791), .I1(n3794), .I2(n3795), .O(n3805));
  LUT3 #(.INIT(8'hE8)) lut_n3806 (.I0(n3801), .I1(n3804), .I2(n3805), .O(n3806));
  LUT3 #(.INIT(8'h96)) lut_n3807 (.I0(x162), .I1(x163), .I2(x164), .O(n3807));
  LUT5 #(.INIT(32'h96696996)) lut_n3808 (.I0(x153), .I1(x154), .I2(x155), .I3(n3802), .I4(n3803), .O(n3808));
  LUT5 #(.INIT(32'hFF969600)) lut_n3809 (.I0(x159), .I1(x160), .I2(x161), .I3(n3807), .I4(n3808), .O(n3809));
  LUT3 #(.INIT(8'h96)) lut_n3810 (.I0(x168), .I1(x169), .I2(x170), .O(n3810));
  LUT5 #(.INIT(32'h96696996)) lut_n3811 (.I0(x159), .I1(x160), .I2(x161), .I3(n3807), .I4(n3808), .O(n3811));
  LUT5 #(.INIT(32'hFF969600)) lut_n3812 (.I0(x165), .I1(x166), .I2(x167), .I3(n3810), .I4(n3811), .O(n3812));
  LUT3 #(.INIT(8'h96)) lut_n3813 (.I0(n3801), .I1(n3804), .I2(n3805), .O(n3813));
  LUT3 #(.INIT(8'hE8)) lut_n3814 (.I0(n3809), .I1(n3812), .I2(n3813), .O(n3814));
  LUT3 #(.INIT(8'h96)) lut_n3815 (.I0(n3788), .I1(n3796), .I2(n3797), .O(n3815));
  LUT3 #(.INIT(8'hE8)) lut_n3816 (.I0(n3806), .I1(n3814), .I2(n3815), .O(n3816));
  LUT3 #(.INIT(8'h96)) lut_n3817 (.I0(n3760), .I1(n3778), .I2(n3779), .O(n3817));
  LUT3 #(.INIT(8'hE8)) lut_n3818 (.I0(n3798), .I1(n3816), .I2(n3817), .O(n3818));
  LUT3 #(.INIT(8'h96)) lut_n3819 (.I0(n3702), .I1(n3740), .I2(n3741), .O(n3819));
  LUT3 #(.INIT(8'hE8)) lut_n3820 (.I0(n3780), .I1(n3818), .I2(n3819), .O(n3820));
  LUT3 #(.INIT(8'h96)) lut_n3821 (.I0(n3634), .I1(n3672), .I2(n3673), .O(n3821));
  LUT3 #(.INIT(8'hE8)) lut_n3822 (.I0(n3742), .I1(n3820), .I2(n3821), .O(n3822));
  LUT3 #(.INIT(8'h96)) lut_n3823 (.I0(n3514), .I1(n3592), .I2(n3593), .O(n3823));
  LUT3 #(.INIT(8'hE8)) lut_n3824 (.I0(n3674), .I1(n3822), .I2(n3823), .O(n3824));
  LUT3 #(.INIT(8'h96)) lut_n3825 (.I0(x174), .I1(x175), .I2(x176), .O(n3825));
  LUT5 #(.INIT(32'h96696996)) lut_n3826 (.I0(x165), .I1(x166), .I2(x167), .I3(n3810), .I4(n3811), .O(n3826));
  LUT5 #(.INIT(32'hFF969600)) lut_n3827 (.I0(x171), .I1(x172), .I2(x173), .I3(n3825), .I4(n3826), .O(n3827));
  LUT3 #(.INIT(8'h96)) lut_n3828 (.I0(x180), .I1(x181), .I2(x182), .O(n3828));
  LUT5 #(.INIT(32'h96696996)) lut_n3829 (.I0(x171), .I1(x172), .I2(x173), .I3(n3825), .I4(n3826), .O(n3829));
  LUT5 #(.INIT(32'hFF969600)) lut_n3830 (.I0(x177), .I1(x178), .I2(x179), .I3(n3828), .I4(n3829), .O(n3830));
  LUT3 #(.INIT(8'h96)) lut_n3831 (.I0(n3809), .I1(n3812), .I2(n3813), .O(n3831));
  LUT3 #(.INIT(8'hE8)) lut_n3832 (.I0(n3827), .I1(n3830), .I2(n3831), .O(n3832));
  LUT3 #(.INIT(8'h96)) lut_n3833 (.I0(x186), .I1(x187), .I2(x188), .O(n3833));
  LUT5 #(.INIT(32'h96696996)) lut_n3834 (.I0(x177), .I1(x178), .I2(x179), .I3(n3828), .I4(n3829), .O(n3834));
  LUT5 #(.INIT(32'hFF969600)) lut_n3835 (.I0(x183), .I1(x184), .I2(x185), .I3(n3833), .I4(n3834), .O(n3835));
  LUT3 #(.INIT(8'h96)) lut_n3836 (.I0(x192), .I1(x193), .I2(x194), .O(n3836));
  LUT5 #(.INIT(32'h96696996)) lut_n3837 (.I0(x183), .I1(x184), .I2(x185), .I3(n3833), .I4(n3834), .O(n3837));
  LUT5 #(.INIT(32'hFF969600)) lut_n3838 (.I0(x189), .I1(x190), .I2(x191), .I3(n3836), .I4(n3837), .O(n3838));
  LUT3 #(.INIT(8'h96)) lut_n3839 (.I0(n3827), .I1(n3830), .I2(n3831), .O(n3839));
  LUT3 #(.INIT(8'hE8)) lut_n3840 (.I0(n3835), .I1(n3838), .I2(n3839), .O(n3840));
  LUT3 #(.INIT(8'h96)) lut_n3841 (.I0(n3806), .I1(n3814), .I2(n3815), .O(n3841));
  LUT3 #(.INIT(8'hE8)) lut_n3842 (.I0(n3832), .I1(n3840), .I2(n3841), .O(n3842));
  LUT3 #(.INIT(8'h96)) lut_n3843 (.I0(x198), .I1(x199), .I2(x200), .O(n3843));
  LUT5 #(.INIT(32'h96696996)) lut_n3844 (.I0(x189), .I1(x190), .I2(x191), .I3(n3836), .I4(n3837), .O(n3844));
  LUT5 #(.INIT(32'hFF969600)) lut_n3845 (.I0(x195), .I1(x196), .I2(x197), .I3(n3843), .I4(n3844), .O(n3845));
  LUT3 #(.INIT(8'h96)) lut_n3846 (.I0(x204), .I1(x205), .I2(x206), .O(n3846));
  LUT5 #(.INIT(32'h96696996)) lut_n3847 (.I0(x195), .I1(x196), .I2(x197), .I3(n3843), .I4(n3844), .O(n3847));
  LUT5 #(.INIT(32'hFF969600)) lut_n3848 (.I0(x201), .I1(x202), .I2(x203), .I3(n3846), .I4(n3847), .O(n3848));
  LUT3 #(.INIT(8'h96)) lut_n3849 (.I0(n3835), .I1(n3838), .I2(n3839), .O(n3849));
  LUT3 #(.INIT(8'hE8)) lut_n3850 (.I0(n3845), .I1(n3848), .I2(n3849), .O(n3850));
  LUT3 #(.INIT(8'h96)) lut_n3851 (.I0(x210), .I1(x211), .I2(x212), .O(n3851));
  LUT5 #(.INIT(32'h96696996)) lut_n3852 (.I0(x201), .I1(x202), .I2(x203), .I3(n3846), .I4(n3847), .O(n3852));
  LUT5 #(.INIT(32'hFF969600)) lut_n3853 (.I0(x207), .I1(x208), .I2(x209), .I3(n3851), .I4(n3852), .O(n3853));
  LUT3 #(.INIT(8'h96)) lut_n3854 (.I0(x216), .I1(x217), .I2(x218), .O(n3854));
  LUT5 #(.INIT(32'h96696996)) lut_n3855 (.I0(x207), .I1(x208), .I2(x209), .I3(n3851), .I4(n3852), .O(n3855));
  LUT5 #(.INIT(32'hFF969600)) lut_n3856 (.I0(x213), .I1(x214), .I2(x215), .I3(n3854), .I4(n3855), .O(n3856));
  LUT3 #(.INIT(8'h96)) lut_n3857 (.I0(n3845), .I1(n3848), .I2(n3849), .O(n3857));
  LUT3 #(.INIT(8'hE8)) lut_n3858 (.I0(n3853), .I1(n3856), .I2(n3857), .O(n3858));
  LUT3 #(.INIT(8'h96)) lut_n3859 (.I0(n3832), .I1(n3840), .I2(n3841), .O(n3859));
  LUT3 #(.INIT(8'hE8)) lut_n3860 (.I0(n3850), .I1(n3858), .I2(n3859), .O(n3860));
  LUT3 #(.INIT(8'h96)) lut_n3861 (.I0(n3798), .I1(n3816), .I2(n3817), .O(n3861));
  LUT3 #(.INIT(8'hE8)) lut_n3862 (.I0(n3842), .I1(n3860), .I2(n3861), .O(n3862));
  LUT3 #(.INIT(8'h96)) lut_n3863 (.I0(x222), .I1(x223), .I2(x224), .O(n3863));
  LUT5 #(.INIT(32'h96696996)) lut_n3864 (.I0(x213), .I1(x214), .I2(x215), .I3(n3854), .I4(n3855), .O(n3864));
  LUT5 #(.INIT(32'hFF969600)) lut_n3865 (.I0(x219), .I1(x220), .I2(x221), .I3(n3863), .I4(n3864), .O(n3865));
  LUT3 #(.INIT(8'h96)) lut_n3866 (.I0(x228), .I1(x229), .I2(x230), .O(n3866));
  LUT5 #(.INIT(32'h96696996)) lut_n3867 (.I0(x219), .I1(x220), .I2(x221), .I3(n3863), .I4(n3864), .O(n3867));
  LUT5 #(.INIT(32'hFF969600)) lut_n3868 (.I0(x225), .I1(x226), .I2(x227), .I3(n3866), .I4(n3867), .O(n3868));
  LUT3 #(.INIT(8'h96)) lut_n3869 (.I0(n3853), .I1(n3856), .I2(n3857), .O(n3869));
  LUT3 #(.INIT(8'hE8)) lut_n3870 (.I0(n3865), .I1(n3868), .I2(n3869), .O(n3870));
  LUT3 #(.INIT(8'h96)) lut_n3871 (.I0(x234), .I1(x235), .I2(x236), .O(n3871));
  LUT5 #(.INIT(32'h96696996)) lut_n3872 (.I0(x225), .I1(x226), .I2(x227), .I3(n3866), .I4(n3867), .O(n3872));
  LUT5 #(.INIT(32'hFF969600)) lut_n3873 (.I0(x231), .I1(x232), .I2(x233), .I3(n3871), .I4(n3872), .O(n3873));
  LUT3 #(.INIT(8'h96)) lut_n3874 (.I0(x240), .I1(x241), .I2(x242), .O(n3874));
  LUT5 #(.INIT(32'h96696996)) lut_n3875 (.I0(x231), .I1(x232), .I2(x233), .I3(n3871), .I4(n3872), .O(n3875));
  LUT5 #(.INIT(32'hFF969600)) lut_n3876 (.I0(x237), .I1(x238), .I2(x239), .I3(n3874), .I4(n3875), .O(n3876));
  LUT3 #(.INIT(8'h96)) lut_n3877 (.I0(n3865), .I1(n3868), .I2(n3869), .O(n3877));
  LUT3 #(.INIT(8'hE8)) lut_n3878 (.I0(n3873), .I1(n3876), .I2(n3877), .O(n3878));
  LUT3 #(.INIT(8'h96)) lut_n3879 (.I0(n3850), .I1(n3858), .I2(n3859), .O(n3879));
  LUT3 #(.INIT(8'hE8)) lut_n3880 (.I0(n3870), .I1(n3878), .I2(n3879), .O(n3880));
  LUT3 #(.INIT(8'h96)) lut_n3881 (.I0(x246), .I1(x247), .I2(x248), .O(n3881));
  LUT5 #(.INIT(32'h96696996)) lut_n3882 (.I0(x237), .I1(x238), .I2(x239), .I3(n3874), .I4(n3875), .O(n3882));
  LUT5 #(.INIT(32'hFF969600)) lut_n3883 (.I0(x243), .I1(x244), .I2(x245), .I3(n3881), .I4(n3882), .O(n3883));
  LUT3 #(.INIT(8'h96)) lut_n3884 (.I0(x252), .I1(x253), .I2(x254), .O(n3884));
  LUT5 #(.INIT(32'h96696996)) lut_n3885 (.I0(x243), .I1(x244), .I2(x245), .I3(n3881), .I4(n3882), .O(n3885));
  LUT5 #(.INIT(32'hFF969600)) lut_n3886 (.I0(x249), .I1(x250), .I2(x251), .I3(n3884), .I4(n3885), .O(n3886));
  LUT3 #(.INIT(8'h96)) lut_n3887 (.I0(n3873), .I1(n3876), .I2(n3877), .O(n3887));
  LUT3 #(.INIT(8'hE8)) lut_n3888 (.I0(n3883), .I1(n3886), .I2(n3887), .O(n3888));
  LUT3 #(.INIT(8'h96)) lut_n3889 (.I0(x258), .I1(x259), .I2(x260), .O(n3889));
  LUT5 #(.INIT(32'h96696996)) lut_n3890 (.I0(x249), .I1(x250), .I2(x251), .I3(n3884), .I4(n3885), .O(n3890));
  LUT5 #(.INIT(32'hFF969600)) lut_n3891 (.I0(x255), .I1(x256), .I2(x257), .I3(n3889), .I4(n3890), .O(n3891));
  LUT3 #(.INIT(8'h96)) lut_n3892 (.I0(x264), .I1(x265), .I2(x266), .O(n3892));
  LUT5 #(.INIT(32'h96696996)) lut_n3893 (.I0(x255), .I1(x256), .I2(x257), .I3(n3889), .I4(n3890), .O(n3893));
  LUT5 #(.INIT(32'hFF969600)) lut_n3894 (.I0(x261), .I1(x262), .I2(x263), .I3(n3892), .I4(n3893), .O(n3894));
  LUT3 #(.INIT(8'h96)) lut_n3895 (.I0(n3883), .I1(n3886), .I2(n3887), .O(n3895));
  LUT3 #(.INIT(8'hE8)) lut_n3896 (.I0(n3891), .I1(n3894), .I2(n3895), .O(n3896));
  LUT3 #(.INIT(8'h96)) lut_n3897 (.I0(n3870), .I1(n3878), .I2(n3879), .O(n3897));
  LUT3 #(.INIT(8'hE8)) lut_n3898 (.I0(n3888), .I1(n3896), .I2(n3897), .O(n3898));
  LUT3 #(.INIT(8'h96)) lut_n3899 (.I0(n3842), .I1(n3860), .I2(n3861), .O(n3899));
  LUT3 #(.INIT(8'hE8)) lut_n3900 (.I0(n3880), .I1(n3898), .I2(n3899), .O(n3900));
  LUT3 #(.INIT(8'h96)) lut_n3901 (.I0(n3780), .I1(n3818), .I2(n3819), .O(n3901));
  LUT3 #(.INIT(8'hE8)) lut_n3902 (.I0(n3862), .I1(n3900), .I2(n3901), .O(n3902));
  LUT3 #(.INIT(8'h96)) lut_n3903 (.I0(x270), .I1(x271), .I2(x272), .O(n3903));
  LUT5 #(.INIT(32'h96696996)) lut_n3904 (.I0(x261), .I1(x262), .I2(x263), .I3(n3892), .I4(n3893), .O(n3904));
  LUT5 #(.INIT(32'hFF969600)) lut_n3905 (.I0(x267), .I1(x268), .I2(x269), .I3(n3903), .I4(n3904), .O(n3905));
  LUT3 #(.INIT(8'h96)) lut_n3906 (.I0(x276), .I1(x277), .I2(x278), .O(n3906));
  LUT5 #(.INIT(32'h96696996)) lut_n3907 (.I0(x267), .I1(x268), .I2(x269), .I3(n3903), .I4(n3904), .O(n3907));
  LUT5 #(.INIT(32'hFF969600)) lut_n3908 (.I0(x273), .I1(x274), .I2(x275), .I3(n3906), .I4(n3907), .O(n3908));
  LUT3 #(.INIT(8'h96)) lut_n3909 (.I0(n3891), .I1(n3894), .I2(n3895), .O(n3909));
  LUT3 #(.INIT(8'hE8)) lut_n3910 (.I0(n3905), .I1(n3908), .I2(n3909), .O(n3910));
  LUT3 #(.INIT(8'h96)) lut_n3911 (.I0(x282), .I1(x283), .I2(x284), .O(n3911));
  LUT5 #(.INIT(32'h96696996)) lut_n3912 (.I0(x273), .I1(x274), .I2(x275), .I3(n3906), .I4(n3907), .O(n3912));
  LUT5 #(.INIT(32'hFF969600)) lut_n3913 (.I0(x279), .I1(x280), .I2(x281), .I3(n3911), .I4(n3912), .O(n3913));
  LUT3 #(.INIT(8'h96)) lut_n3914 (.I0(x288), .I1(x289), .I2(x290), .O(n3914));
  LUT5 #(.INIT(32'h96696996)) lut_n3915 (.I0(x279), .I1(x280), .I2(x281), .I3(n3911), .I4(n3912), .O(n3915));
  LUT5 #(.INIT(32'hFF969600)) lut_n3916 (.I0(x285), .I1(x286), .I2(x287), .I3(n3914), .I4(n3915), .O(n3916));
  LUT3 #(.INIT(8'h96)) lut_n3917 (.I0(n3905), .I1(n3908), .I2(n3909), .O(n3917));
  LUT3 #(.INIT(8'hE8)) lut_n3918 (.I0(n3913), .I1(n3916), .I2(n3917), .O(n3918));
  LUT3 #(.INIT(8'h96)) lut_n3919 (.I0(n3888), .I1(n3896), .I2(n3897), .O(n3919));
  LUT3 #(.INIT(8'hE8)) lut_n3920 (.I0(n3910), .I1(n3918), .I2(n3919), .O(n3920));
  LUT3 #(.INIT(8'h96)) lut_n3921 (.I0(x294), .I1(x295), .I2(x296), .O(n3921));
  LUT5 #(.INIT(32'h96696996)) lut_n3922 (.I0(x285), .I1(x286), .I2(x287), .I3(n3914), .I4(n3915), .O(n3922));
  LUT5 #(.INIT(32'hFF969600)) lut_n3923 (.I0(x291), .I1(x292), .I2(x293), .I3(n3921), .I4(n3922), .O(n3923));
  LUT3 #(.INIT(8'h96)) lut_n3924 (.I0(x297), .I1(x298), .I2(x299), .O(n3924));
  LUT5 #(.INIT(32'h96696996)) lut_n3925 (.I0(x291), .I1(x292), .I2(x293), .I3(n3921), .I4(n3922), .O(n3925));
  LUT5 #(.INIT(32'hFF969600)) lut_n3926 (.I0(x300), .I1(x301), .I2(x302), .I3(n3924), .I4(n3925), .O(n3926));
  LUT3 #(.INIT(8'h96)) lut_n3927 (.I0(n3913), .I1(n3916), .I2(n3917), .O(n3927));
  LUT3 #(.INIT(8'hE8)) lut_n3928 (.I0(n3923), .I1(n3926), .I2(n3927), .O(n3928));
  LUT3 #(.INIT(8'h96)) lut_n3929 (.I0(x306), .I1(x307), .I2(x308), .O(n3929));
  LUT5 #(.INIT(32'h96696996)) lut_n3930 (.I0(x300), .I1(x301), .I2(x302), .I3(n3924), .I4(n3925), .O(n3930));
  LUT5 #(.INIT(32'hFF969600)) lut_n3931 (.I0(x303), .I1(x304), .I2(x305), .I3(n3929), .I4(n3930), .O(n3931));
  LUT3 #(.INIT(8'h96)) lut_n3932 (.I0(x312), .I1(x313), .I2(x314), .O(n3932));
  LUT5 #(.INIT(32'h96696996)) lut_n3933 (.I0(x303), .I1(x304), .I2(x305), .I3(n3929), .I4(n3930), .O(n3933));
  LUT5 #(.INIT(32'hFF969600)) lut_n3934 (.I0(x309), .I1(x310), .I2(x311), .I3(n3932), .I4(n3933), .O(n3934));
  LUT3 #(.INIT(8'h96)) lut_n3935 (.I0(n3923), .I1(n3926), .I2(n3927), .O(n3935));
  LUT3 #(.INIT(8'hE8)) lut_n3936 (.I0(n3931), .I1(n3934), .I2(n3935), .O(n3936));
  LUT3 #(.INIT(8'h96)) lut_n3937 (.I0(n3910), .I1(n3918), .I2(n3919), .O(n3937));
  LUT3 #(.INIT(8'hE8)) lut_n3938 (.I0(n3928), .I1(n3936), .I2(n3937), .O(n3938));
  LUT3 #(.INIT(8'h96)) lut_n3939 (.I0(n3880), .I1(n3898), .I2(n3899), .O(n3939));
  LUT3 #(.INIT(8'hE8)) lut_n3940 (.I0(n3920), .I1(n3938), .I2(n3939), .O(n3940));
  LUT3 #(.INIT(8'h96)) lut_n3941 (.I0(x318), .I1(x319), .I2(x320), .O(n3941));
  LUT5 #(.INIT(32'h96696996)) lut_n3942 (.I0(x309), .I1(x310), .I2(x311), .I3(n3932), .I4(n3933), .O(n3942));
  LUT5 #(.INIT(32'hFF969600)) lut_n3943 (.I0(x315), .I1(x316), .I2(x317), .I3(n3941), .I4(n3942), .O(n3943));
  LUT3 #(.INIT(8'h96)) lut_n3944 (.I0(x324), .I1(x325), .I2(x326), .O(n3944));
  LUT5 #(.INIT(32'h96696996)) lut_n3945 (.I0(x315), .I1(x316), .I2(x317), .I3(n3941), .I4(n3942), .O(n3945));
  LUT5 #(.INIT(32'hFF969600)) lut_n3946 (.I0(x321), .I1(x322), .I2(x323), .I3(n3944), .I4(n3945), .O(n3946));
  LUT3 #(.INIT(8'h96)) lut_n3947 (.I0(n3931), .I1(n3934), .I2(n3935), .O(n3947));
  LUT3 #(.INIT(8'hE8)) lut_n3948 (.I0(n3943), .I1(n3946), .I2(n3947), .O(n3948));
  LUT3 #(.INIT(8'h96)) lut_n3949 (.I0(x330), .I1(x331), .I2(x332), .O(n3949));
  LUT5 #(.INIT(32'h96696996)) lut_n3950 (.I0(x321), .I1(x322), .I2(x323), .I3(n3944), .I4(n3945), .O(n3950));
  LUT5 #(.INIT(32'hFF969600)) lut_n3951 (.I0(x327), .I1(x328), .I2(x329), .I3(n3949), .I4(n3950), .O(n3951));
  LUT3 #(.INIT(8'h96)) lut_n3952 (.I0(x336), .I1(x337), .I2(x338), .O(n3952));
  LUT5 #(.INIT(32'h96696996)) lut_n3953 (.I0(x327), .I1(x328), .I2(x329), .I3(n3949), .I4(n3950), .O(n3953));
  LUT5 #(.INIT(32'hFF969600)) lut_n3954 (.I0(x333), .I1(x334), .I2(x335), .I3(n3952), .I4(n3953), .O(n3954));
  LUT3 #(.INIT(8'h96)) lut_n3955 (.I0(n3943), .I1(n3946), .I2(n3947), .O(n3955));
  LUT3 #(.INIT(8'hE8)) lut_n3956 (.I0(n3951), .I1(n3954), .I2(n3955), .O(n3956));
  LUT3 #(.INIT(8'h96)) lut_n3957 (.I0(n3928), .I1(n3936), .I2(n3937), .O(n3957));
  LUT3 #(.INIT(8'hE8)) lut_n3958 (.I0(n3948), .I1(n3956), .I2(n3957), .O(n3958));
  LUT3 #(.INIT(8'h96)) lut_n3959 (.I0(x342), .I1(x343), .I2(x344), .O(n3959));
  LUT5 #(.INIT(32'h96696996)) lut_n3960 (.I0(x333), .I1(x334), .I2(x335), .I3(n3952), .I4(n3953), .O(n3960));
  LUT5 #(.INIT(32'hFF969600)) lut_n3961 (.I0(x339), .I1(x340), .I2(x341), .I3(n3959), .I4(n3960), .O(n3961));
  LUT3 #(.INIT(8'h96)) lut_n3962 (.I0(x348), .I1(x349), .I2(x350), .O(n3962));
  LUT5 #(.INIT(32'h96696996)) lut_n3963 (.I0(x339), .I1(x340), .I2(x341), .I3(n3959), .I4(n3960), .O(n3963));
  LUT5 #(.INIT(32'hFF969600)) lut_n3964 (.I0(x345), .I1(x346), .I2(x347), .I3(n3962), .I4(n3963), .O(n3964));
  LUT3 #(.INIT(8'h96)) lut_n3965 (.I0(n3951), .I1(n3954), .I2(n3955), .O(n3965));
  LUT3 #(.INIT(8'hE8)) lut_n3966 (.I0(n3961), .I1(n3964), .I2(n3965), .O(n3966));
  LUT3 #(.INIT(8'h96)) lut_n3967 (.I0(x354), .I1(x355), .I2(x356), .O(n3967));
  LUT5 #(.INIT(32'h96696996)) lut_n3968 (.I0(x345), .I1(x346), .I2(x347), .I3(n3962), .I4(n3963), .O(n3968));
  LUT5 #(.INIT(32'hFF969600)) lut_n3969 (.I0(x351), .I1(x352), .I2(x353), .I3(n3967), .I4(n3968), .O(n3969));
  LUT3 #(.INIT(8'h96)) lut_n3970 (.I0(x360), .I1(x361), .I2(x362), .O(n3970));
  LUT5 #(.INIT(32'h96696996)) lut_n3971 (.I0(x351), .I1(x352), .I2(x353), .I3(n3967), .I4(n3968), .O(n3971));
  LUT5 #(.INIT(32'hFF969600)) lut_n3972 (.I0(x357), .I1(x358), .I2(x359), .I3(n3970), .I4(n3971), .O(n3972));
  LUT3 #(.INIT(8'h96)) lut_n3973 (.I0(n3961), .I1(n3964), .I2(n3965), .O(n3973));
  LUT3 #(.INIT(8'hE8)) lut_n3974 (.I0(n3969), .I1(n3972), .I2(n3973), .O(n3974));
  LUT3 #(.INIT(8'h96)) lut_n3975 (.I0(n3948), .I1(n3956), .I2(n3957), .O(n3975));
  LUT3 #(.INIT(8'hE8)) lut_n3976 (.I0(n3966), .I1(n3974), .I2(n3975), .O(n3976));
  LUT3 #(.INIT(8'h96)) lut_n3977 (.I0(n3920), .I1(n3938), .I2(n3939), .O(n3977));
  LUT3 #(.INIT(8'hE8)) lut_n3978 (.I0(n3958), .I1(n3976), .I2(n3977), .O(n3978));
  LUT3 #(.INIT(8'h96)) lut_n3979 (.I0(n3862), .I1(n3900), .I2(n3901), .O(n3979));
  LUT3 #(.INIT(8'hE8)) lut_n3980 (.I0(n3940), .I1(n3978), .I2(n3979), .O(n3980));
  LUT3 #(.INIT(8'h96)) lut_n3981 (.I0(n3742), .I1(n3820), .I2(n3821), .O(n3981));
  LUT3 #(.INIT(8'hE8)) lut_n3982 (.I0(n3902), .I1(n3980), .I2(n3981), .O(n3982));
  LUT3 #(.INIT(8'h96)) lut_n3983 (.I0(x366), .I1(x367), .I2(x368), .O(n3983));
  LUT5 #(.INIT(32'h96696996)) lut_n3984 (.I0(x357), .I1(x358), .I2(x359), .I3(n3970), .I4(n3971), .O(n3984));
  LUT5 #(.INIT(32'hFF969600)) lut_n3985 (.I0(x363), .I1(x364), .I2(x365), .I3(n3983), .I4(n3984), .O(n3985));
  LUT3 #(.INIT(8'h96)) lut_n3986 (.I0(x372), .I1(x373), .I2(x374), .O(n3986));
  LUT5 #(.INIT(32'h96696996)) lut_n3987 (.I0(x363), .I1(x364), .I2(x365), .I3(n3983), .I4(n3984), .O(n3987));
  LUT5 #(.INIT(32'hFF969600)) lut_n3988 (.I0(x369), .I1(x370), .I2(x371), .I3(n3986), .I4(n3987), .O(n3988));
  LUT3 #(.INIT(8'h96)) lut_n3989 (.I0(n3969), .I1(n3972), .I2(n3973), .O(n3989));
  LUT3 #(.INIT(8'hE8)) lut_n3990 (.I0(n3985), .I1(n3988), .I2(n3989), .O(n3990));
  LUT3 #(.INIT(8'h96)) lut_n3991 (.I0(x378), .I1(x379), .I2(x380), .O(n3991));
  LUT5 #(.INIT(32'h96696996)) lut_n3992 (.I0(x369), .I1(x370), .I2(x371), .I3(n3986), .I4(n3987), .O(n3992));
  LUT5 #(.INIT(32'hFF969600)) lut_n3993 (.I0(x375), .I1(x376), .I2(x377), .I3(n3991), .I4(n3992), .O(n3993));
  LUT3 #(.INIT(8'h96)) lut_n3994 (.I0(x384), .I1(x385), .I2(x386), .O(n3994));
  LUT5 #(.INIT(32'h96696996)) lut_n3995 (.I0(x375), .I1(x376), .I2(x377), .I3(n3991), .I4(n3992), .O(n3995));
  LUT5 #(.INIT(32'hFF969600)) lut_n3996 (.I0(x381), .I1(x382), .I2(x383), .I3(n3994), .I4(n3995), .O(n3996));
  LUT3 #(.INIT(8'h96)) lut_n3997 (.I0(n3985), .I1(n3988), .I2(n3989), .O(n3997));
  LUT3 #(.INIT(8'hE8)) lut_n3998 (.I0(n3993), .I1(n3996), .I2(n3997), .O(n3998));
  LUT3 #(.INIT(8'h96)) lut_n3999 (.I0(n3966), .I1(n3974), .I2(n3975), .O(n3999));
  LUT3 #(.INIT(8'hE8)) lut_n4000 (.I0(n3990), .I1(n3998), .I2(n3999), .O(n4000));
  LUT3 #(.INIT(8'h96)) lut_n4001 (.I0(x390), .I1(x391), .I2(x392), .O(n4001));
  LUT5 #(.INIT(32'h96696996)) lut_n4002 (.I0(x381), .I1(x382), .I2(x383), .I3(n3994), .I4(n3995), .O(n4002));
  LUT5 #(.INIT(32'hFF969600)) lut_n4003 (.I0(x387), .I1(x388), .I2(x389), .I3(n4001), .I4(n4002), .O(n4003));
  LUT3 #(.INIT(8'h96)) lut_n4004 (.I0(x396), .I1(x397), .I2(x398), .O(n4004));
  LUT5 #(.INIT(32'h96696996)) lut_n4005 (.I0(x387), .I1(x388), .I2(x389), .I3(n4001), .I4(n4002), .O(n4005));
  LUT5 #(.INIT(32'hFF969600)) lut_n4006 (.I0(x393), .I1(x394), .I2(x395), .I3(n4004), .I4(n4005), .O(n4006));
  LUT3 #(.INIT(8'h96)) lut_n4007 (.I0(n3993), .I1(n3996), .I2(n3997), .O(n4007));
  LUT3 #(.INIT(8'hE8)) lut_n4008 (.I0(n4003), .I1(n4006), .I2(n4007), .O(n4008));
  LUT3 #(.INIT(8'h96)) lut_n4009 (.I0(x402), .I1(x403), .I2(x404), .O(n4009));
  LUT5 #(.INIT(32'h96696996)) lut_n4010 (.I0(x393), .I1(x394), .I2(x395), .I3(n4004), .I4(n4005), .O(n4010));
  LUT5 #(.INIT(32'hFF969600)) lut_n4011 (.I0(x399), .I1(x400), .I2(x401), .I3(n4009), .I4(n4010), .O(n4011));
  LUT3 #(.INIT(8'h96)) lut_n4012 (.I0(x408), .I1(x409), .I2(x410), .O(n4012));
  LUT5 #(.INIT(32'h96696996)) lut_n4013 (.I0(x399), .I1(x400), .I2(x401), .I3(n4009), .I4(n4010), .O(n4013));
  LUT5 #(.INIT(32'hFF969600)) lut_n4014 (.I0(x405), .I1(x406), .I2(x407), .I3(n4012), .I4(n4013), .O(n4014));
  LUT3 #(.INIT(8'h96)) lut_n4015 (.I0(n4003), .I1(n4006), .I2(n4007), .O(n4015));
  LUT3 #(.INIT(8'hE8)) lut_n4016 (.I0(n4011), .I1(n4014), .I2(n4015), .O(n4016));
  LUT3 #(.INIT(8'h96)) lut_n4017 (.I0(n3990), .I1(n3998), .I2(n3999), .O(n4017));
  LUT3 #(.INIT(8'hE8)) lut_n4018 (.I0(n4008), .I1(n4016), .I2(n4017), .O(n4018));
  LUT3 #(.INIT(8'h96)) lut_n4019 (.I0(n3958), .I1(n3976), .I2(n3977), .O(n4019));
  LUT3 #(.INIT(8'hE8)) lut_n4020 (.I0(n4000), .I1(n4018), .I2(n4019), .O(n4020));
  LUT3 #(.INIT(8'h96)) lut_n4021 (.I0(x414), .I1(x415), .I2(x416), .O(n4021));
  LUT5 #(.INIT(32'h96696996)) lut_n4022 (.I0(x405), .I1(x406), .I2(x407), .I3(n4012), .I4(n4013), .O(n4022));
  LUT5 #(.INIT(32'hFF969600)) lut_n4023 (.I0(x411), .I1(x412), .I2(x413), .I3(n4021), .I4(n4022), .O(n4023));
  LUT3 #(.INIT(8'h96)) lut_n4024 (.I0(x420), .I1(x421), .I2(x422), .O(n4024));
  LUT5 #(.INIT(32'h96696996)) lut_n4025 (.I0(x411), .I1(x412), .I2(x413), .I3(n4021), .I4(n4022), .O(n4025));
  LUT5 #(.INIT(32'hFF969600)) lut_n4026 (.I0(x417), .I1(x418), .I2(x419), .I3(n4024), .I4(n4025), .O(n4026));
  LUT3 #(.INIT(8'h96)) lut_n4027 (.I0(n4011), .I1(n4014), .I2(n4015), .O(n4027));
  LUT3 #(.INIT(8'hE8)) lut_n4028 (.I0(n4023), .I1(n4026), .I2(n4027), .O(n4028));
  LUT3 #(.INIT(8'h96)) lut_n4029 (.I0(x426), .I1(x427), .I2(x428), .O(n4029));
  LUT5 #(.INIT(32'h96696996)) lut_n4030 (.I0(x417), .I1(x418), .I2(x419), .I3(n4024), .I4(n4025), .O(n4030));
  LUT5 #(.INIT(32'hFF969600)) lut_n4031 (.I0(x423), .I1(x424), .I2(x425), .I3(n4029), .I4(n4030), .O(n4031));
  LUT3 #(.INIT(8'h96)) lut_n4032 (.I0(x432), .I1(x433), .I2(x434), .O(n4032));
  LUT5 #(.INIT(32'h96696996)) lut_n4033 (.I0(x423), .I1(x424), .I2(x425), .I3(n4029), .I4(n4030), .O(n4033));
  LUT5 #(.INIT(32'hFF969600)) lut_n4034 (.I0(x429), .I1(x430), .I2(x431), .I3(n4032), .I4(n4033), .O(n4034));
  LUT3 #(.INIT(8'h96)) lut_n4035 (.I0(n4023), .I1(n4026), .I2(n4027), .O(n4035));
  LUT3 #(.INIT(8'hE8)) lut_n4036 (.I0(n4031), .I1(n4034), .I2(n4035), .O(n4036));
  LUT3 #(.INIT(8'h96)) lut_n4037 (.I0(n4008), .I1(n4016), .I2(n4017), .O(n4037));
  LUT3 #(.INIT(8'hE8)) lut_n4038 (.I0(n4028), .I1(n4036), .I2(n4037), .O(n4038));
  LUT3 #(.INIT(8'h96)) lut_n4039 (.I0(x438), .I1(x439), .I2(x440), .O(n4039));
  LUT5 #(.INIT(32'h96696996)) lut_n4040 (.I0(x429), .I1(x430), .I2(x431), .I3(n4032), .I4(n4033), .O(n4040));
  LUT5 #(.INIT(32'hFF969600)) lut_n4041 (.I0(x435), .I1(x436), .I2(x437), .I3(n4039), .I4(n4040), .O(n4041));
  LUT3 #(.INIT(8'h96)) lut_n4042 (.I0(x444), .I1(x445), .I2(x446), .O(n4042));
  LUT5 #(.INIT(32'h96696996)) lut_n4043 (.I0(x435), .I1(x436), .I2(x437), .I3(n4039), .I4(n4040), .O(n4043));
  LUT5 #(.INIT(32'hFF969600)) lut_n4044 (.I0(x441), .I1(x442), .I2(x443), .I3(n4042), .I4(n4043), .O(n4044));
  LUT3 #(.INIT(8'h96)) lut_n4045 (.I0(n4031), .I1(n4034), .I2(n4035), .O(n4045));
  LUT3 #(.INIT(8'hE8)) lut_n4046 (.I0(n4041), .I1(n4044), .I2(n4045), .O(n4046));
  LUT3 #(.INIT(8'h96)) lut_n4047 (.I0(x450), .I1(x451), .I2(x452), .O(n4047));
  LUT5 #(.INIT(32'h96696996)) lut_n4048 (.I0(x441), .I1(x442), .I2(x443), .I3(n4042), .I4(n4043), .O(n4048));
  LUT5 #(.INIT(32'hFF969600)) lut_n4049 (.I0(x447), .I1(x448), .I2(x449), .I3(n4047), .I4(n4048), .O(n4049));
  LUT3 #(.INIT(8'h96)) lut_n4050 (.I0(x456), .I1(x457), .I2(x458), .O(n4050));
  LUT5 #(.INIT(32'h96696996)) lut_n4051 (.I0(x447), .I1(x448), .I2(x449), .I3(n4047), .I4(n4048), .O(n4051));
  LUT5 #(.INIT(32'hFF969600)) lut_n4052 (.I0(x453), .I1(x454), .I2(x455), .I3(n4050), .I4(n4051), .O(n4052));
  LUT3 #(.INIT(8'h96)) lut_n4053 (.I0(n4041), .I1(n4044), .I2(n4045), .O(n4053));
  LUT3 #(.INIT(8'hE8)) lut_n4054 (.I0(n4049), .I1(n4052), .I2(n4053), .O(n4054));
  LUT3 #(.INIT(8'h96)) lut_n4055 (.I0(n4028), .I1(n4036), .I2(n4037), .O(n4055));
  LUT3 #(.INIT(8'hE8)) lut_n4056 (.I0(n4046), .I1(n4054), .I2(n4055), .O(n4056));
  LUT3 #(.INIT(8'h96)) lut_n4057 (.I0(n4000), .I1(n4018), .I2(n4019), .O(n4057));
  LUT3 #(.INIT(8'hE8)) lut_n4058 (.I0(n4038), .I1(n4056), .I2(n4057), .O(n4058));
  LUT3 #(.INIT(8'h96)) lut_n4059 (.I0(n3940), .I1(n3978), .I2(n3979), .O(n4059));
  LUT3 #(.INIT(8'hE8)) lut_n4060 (.I0(n4020), .I1(n4058), .I2(n4059), .O(n4060));
  LUT3 #(.INIT(8'h96)) lut_n4061 (.I0(x462), .I1(x463), .I2(x464), .O(n4061));
  LUT5 #(.INIT(32'h96696996)) lut_n4062 (.I0(x453), .I1(x454), .I2(x455), .I3(n4050), .I4(n4051), .O(n4062));
  LUT5 #(.INIT(32'hFF969600)) lut_n4063 (.I0(x459), .I1(x460), .I2(x461), .I3(n4061), .I4(n4062), .O(n4063));
  LUT3 #(.INIT(8'h96)) lut_n4064 (.I0(x468), .I1(x469), .I2(x470), .O(n4064));
  LUT5 #(.INIT(32'h96696996)) lut_n4065 (.I0(x459), .I1(x460), .I2(x461), .I3(n4061), .I4(n4062), .O(n4065));
  LUT5 #(.INIT(32'hFF969600)) lut_n4066 (.I0(x465), .I1(x466), .I2(x467), .I3(n4064), .I4(n4065), .O(n4066));
  LUT3 #(.INIT(8'h96)) lut_n4067 (.I0(n4049), .I1(n4052), .I2(n4053), .O(n4067));
  LUT3 #(.INIT(8'hE8)) lut_n4068 (.I0(n4063), .I1(n4066), .I2(n4067), .O(n4068));
  LUT3 #(.INIT(8'h96)) lut_n4069 (.I0(x474), .I1(x475), .I2(x476), .O(n4069));
  LUT5 #(.INIT(32'h96696996)) lut_n4070 (.I0(x465), .I1(x466), .I2(x467), .I3(n4064), .I4(n4065), .O(n4070));
  LUT5 #(.INIT(32'hFF969600)) lut_n4071 (.I0(x471), .I1(x472), .I2(x473), .I3(n4069), .I4(n4070), .O(n4071));
  LUT3 #(.INIT(8'h96)) lut_n4072 (.I0(x480), .I1(x481), .I2(x482), .O(n4072));
  LUT5 #(.INIT(32'h96696996)) lut_n4073 (.I0(x471), .I1(x472), .I2(x473), .I3(n4069), .I4(n4070), .O(n4073));
  LUT5 #(.INIT(32'hFF969600)) lut_n4074 (.I0(x477), .I1(x478), .I2(x479), .I3(n4072), .I4(n4073), .O(n4074));
  LUT3 #(.INIT(8'h96)) lut_n4075 (.I0(n4063), .I1(n4066), .I2(n4067), .O(n4075));
  LUT3 #(.INIT(8'hE8)) lut_n4076 (.I0(n4071), .I1(n4074), .I2(n4075), .O(n4076));
  LUT3 #(.INIT(8'h96)) lut_n4077 (.I0(n4046), .I1(n4054), .I2(n4055), .O(n4077));
  LUT3 #(.INIT(8'hE8)) lut_n4078 (.I0(n4068), .I1(n4076), .I2(n4077), .O(n4078));
  LUT3 #(.INIT(8'h96)) lut_n4079 (.I0(x486), .I1(x487), .I2(x488), .O(n4079));
  LUT5 #(.INIT(32'h96696996)) lut_n4080 (.I0(x477), .I1(x478), .I2(x479), .I3(n4072), .I4(n4073), .O(n4080));
  LUT5 #(.INIT(32'hFF969600)) lut_n4081 (.I0(x483), .I1(x484), .I2(x485), .I3(n4079), .I4(n4080), .O(n4081));
  LUT3 #(.INIT(8'h96)) lut_n4082 (.I0(x492), .I1(x493), .I2(x494), .O(n4082));
  LUT5 #(.INIT(32'h96696996)) lut_n4083 (.I0(x483), .I1(x484), .I2(x485), .I3(n4079), .I4(n4080), .O(n4083));
  LUT5 #(.INIT(32'hFF969600)) lut_n4084 (.I0(x489), .I1(x490), .I2(x491), .I3(n4082), .I4(n4083), .O(n4084));
  LUT3 #(.INIT(8'h96)) lut_n4085 (.I0(n4071), .I1(n4074), .I2(n4075), .O(n4085));
  LUT3 #(.INIT(8'hE8)) lut_n4086 (.I0(n4081), .I1(n4084), .I2(n4085), .O(n4086));
  LUT3 #(.INIT(8'h96)) lut_n4087 (.I0(x498), .I1(x499), .I2(x500), .O(n4087));
  LUT5 #(.INIT(32'h96696996)) lut_n4088 (.I0(x489), .I1(x490), .I2(x491), .I3(n4082), .I4(n4083), .O(n4088));
  LUT5 #(.INIT(32'hFF969600)) lut_n4089 (.I0(x495), .I1(x496), .I2(x497), .I3(n4087), .I4(n4088), .O(n4089));
  LUT3 #(.INIT(8'h96)) lut_n4090 (.I0(x504), .I1(x505), .I2(x506), .O(n4090));
  LUT5 #(.INIT(32'h96696996)) lut_n4091 (.I0(x495), .I1(x496), .I2(x497), .I3(n4087), .I4(n4088), .O(n4091));
  LUT5 #(.INIT(32'hFF969600)) lut_n4092 (.I0(x501), .I1(x502), .I2(x503), .I3(n4090), .I4(n4091), .O(n4092));
  LUT3 #(.INIT(8'h96)) lut_n4093 (.I0(n4081), .I1(n4084), .I2(n4085), .O(n4093));
  LUT3 #(.INIT(8'hE8)) lut_n4094 (.I0(n4089), .I1(n4092), .I2(n4093), .O(n4094));
  LUT3 #(.INIT(8'h96)) lut_n4095 (.I0(n4068), .I1(n4076), .I2(n4077), .O(n4095));
  LUT3 #(.INIT(8'hE8)) lut_n4096 (.I0(n4086), .I1(n4094), .I2(n4095), .O(n4096));
  LUT3 #(.INIT(8'h96)) lut_n4097 (.I0(n4038), .I1(n4056), .I2(n4057), .O(n4097));
  LUT3 #(.INIT(8'hE8)) lut_n4098 (.I0(n4078), .I1(n4096), .I2(n4097), .O(n4098));
  LUT3 #(.INIT(8'h96)) lut_n4099 (.I0(x510), .I1(x511), .I2(x512), .O(n4099));
  LUT5 #(.INIT(32'h96696996)) lut_n4100 (.I0(x501), .I1(x502), .I2(x503), .I3(n4090), .I4(n4091), .O(n4100));
  LUT5 #(.INIT(32'hFF969600)) lut_n4101 (.I0(x507), .I1(x508), .I2(x509), .I3(n4099), .I4(n4100), .O(n4101));
  LUT3 #(.INIT(8'h96)) lut_n4102 (.I0(x516), .I1(x517), .I2(x518), .O(n4102));
  LUT5 #(.INIT(32'h96696996)) lut_n4103 (.I0(x507), .I1(x508), .I2(x509), .I3(n4099), .I4(n4100), .O(n4103));
  LUT5 #(.INIT(32'hFF969600)) lut_n4104 (.I0(x513), .I1(x514), .I2(x515), .I3(n4102), .I4(n4103), .O(n4104));
  LUT3 #(.INIT(8'h96)) lut_n4105 (.I0(n4089), .I1(n4092), .I2(n4093), .O(n4105));
  LUT3 #(.INIT(8'hE8)) lut_n4106 (.I0(n4101), .I1(n4104), .I2(n4105), .O(n4106));
  LUT3 #(.INIT(8'h96)) lut_n4107 (.I0(x522), .I1(x523), .I2(x524), .O(n4107));
  LUT5 #(.INIT(32'h96696996)) lut_n4108 (.I0(x513), .I1(x514), .I2(x515), .I3(n4102), .I4(n4103), .O(n4108));
  LUT5 #(.INIT(32'hFF969600)) lut_n4109 (.I0(x519), .I1(x520), .I2(x521), .I3(n4107), .I4(n4108), .O(n4109));
  LUT3 #(.INIT(8'h96)) lut_n4110 (.I0(x528), .I1(x529), .I2(x530), .O(n4110));
  LUT5 #(.INIT(32'h96696996)) lut_n4111 (.I0(x519), .I1(x520), .I2(x521), .I3(n4107), .I4(n4108), .O(n4111));
  LUT5 #(.INIT(32'hFF969600)) lut_n4112 (.I0(x525), .I1(x526), .I2(x527), .I3(n4110), .I4(n4111), .O(n4112));
  LUT3 #(.INIT(8'h96)) lut_n4113 (.I0(n4101), .I1(n4104), .I2(n4105), .O(n4113));
  LUT3 #(.INIT(8'hE8)) lut_n4114 (.I0(n4109), .I1(n4112), .I2(n4113), .O(n4114));
  LUT3 #(.INIT(8'h96)) lut_n4115 (.I0(n4086), .I1(n4094), .I2(n4095), .O(n4115));
  LUT3 #(.INIT(8'hE8)) lut_n4116 (.I0(n4106), .I1(n4114), .I2(n4115), .O(n4116));
  LUT3 #(.INIT(8'h96)) lut_n4117 (.I0(x534), .I1(x535), .I2(x536), .O(n4117));
  LUT5 #(.INIT(32'h96696996)) lut_n4118 (.I0(x525), .I1(x526), .I2(x527), .I3(n4110), .I4(n4111), .O(n4118));
  LUT5 #(.INIT(32'hFF969600)) lut_n4119 (.I0(x531), .I1(x532), .I2(x533), .I3(n4117), .I4(n4118), .O(n4119));
  LUT3 #(.INIT(8'h96)) lut_n4120 (.I0(x540), .I1(x541), .I2(x542), .O(n4120));
  LUT5 #(.INIT(32'h96696996)) lut_n4121 (.I0(x531), .I1(x532), .I2(x533), .I3(n4117), .I4(n4118), .O(n4121));
  LUT5 #(.INIT(32'hFF969600)) lut_n4122 (.I0(x537), .I1(x538), .I2(x539), .I3(n4120), .I4(n4121), .O(n4122));
  LUT3 #(.INIT(8'h96)) lut_n4123 (.I0(n4109), .I1(n4112), .I2(n4113), .O(n4123));
  LUT3 #(.INIT(8'hE8)) lut_n4124 (.I0(n4119), .I1(n4122), .I2(n4123), .O(n4124));
  LUT3 #(.INIT(8'h96)) lut_n4125 (.I0(x546), .I1(x547), .I2(x548), .O(n4125));
  LUT5 #(.INIT(32'h96696996)) lut_n4126 (.I0(x537), .I1(x538), .I2(x539), .I3(n4120), .I4(n4121), .O(n4126));
  LUT5 #(.INIT(32'hFF969600)) lut_n4127 (.I0(x543), .I1(x544), .I2(x545), .I3(n4125), .I4(n4126), .O(n4127));
  LUT3 #(.INIT(8'h96)) lut_n4128 (.I0(x552), .I1(x553), .I2(x554), .O(n4128));
  LUT5 #(.INIT(32'h96696996)) lut_n4129 (.I0(x543), .I1(x544), .I2(x545), .I3(n4125), .I4(n4126), .O(n4129));
  LUT5 #(.INIT(32'hFF969600)) lut_n4130 (.I0(x549), .I1(x550), .I2(x551), .I3(n4128), .I4(n4129), .O(n4130));
  LUT3 #(.INIT(8'h96)) lut_n4131 (.I0(n4119), .I1(n4122), .I2(n4123), .O(n4131));
  LUT3 #(.INIT(8'hE8)) lut_n4132 (.I0(n4127), .I1(n4130), .I2(n4131), .O(n4132));
  LUT3 #(.INIT(8'h96)) lut_n4133 (.I0(n4106), .I1(n4114), .I2(n4115), .O(n4133));
  LUT3 #(.INIT(8'hE8)) lut_n4134 (.I0(n4124), .I1(n4132), .I2(n4133), .O(n4134));
  LUT3 #(.INIT(8'h96)) lut_n4135 (.I0(n4078), .I1(n4096), .I2(n4097), .O(n4135));
  LUT3 #(.INIT(8'hE8)) lut_n4136 (.I0(n4116), .I1(n4134), .I2(n4135), .O(n4136));
  LUT3 #(.INIT(8'h96)) lut_n4137 (.I0(n4020), .I1(n4058), .I2(n4059), .O(n4137));
  LUT3 #(.INIT(8'hE8)) lut_n4138 (.I0(n4098), .I1(n4136), .I2(n4137), .O(n4138));
  LUT3 #(.INIT(8'h96)) lut_n4139 (.I0(n3902), .I1(n3980), .I2(n3981), .O(n4139));
  LUT3 #(.INIT(8'hE8)) lut_n4140 (.I0(n4060), .I1(n4138), .I2(n4139), .O(n4140));
  LUT3 #(.INIT(8'h96)) lut_n4141 (.I0(n3674), .I1(n3822), .I2(n3823), .O(n4141));
  LUT3 #(.INIT(8'hE8)) lut_n4142 (.I0(n3982), .I1(n4140), .I2(n4141), .O(n4142));
  LUT3 #(.INIT(8'h96)) lut_n4143 (.I0(n3436), .I1(n3594), .I2(n3595), .O(n4143));
  LUT3 #(.INIT(8'hE8)) lut_n4144 (.I0(n3824), .I1(n4142), .I2(n4143), .O(n4144));
  LUT3 #(.INIT(8'h96)) lut_n4145 (.I0(n2641), .I1(n2959), .I2(n3277), .O(n4145));
  LUT3 #(.INIT(8'hE8)) lut_n4146 (.I0(n3596), .I1(n4144), .I2(n4145), .O(n4146));
  LUT3 #(.INIT(8'h96)) lut_n4147 (.I0(x558), .I1(x559), .I2(x560), .O(n4147));
  LUT5 #(.INIT(32'h96696996)) lut_n4148 (.I0(x549), .I1(x550), .I2(x551), .I3(n4128), .I4(n4129), .O(n4148));
  LUT5 #(.INIT(32'hFF969600)) lut_n4149 (.I0(x555), .I1(x556), .I2(x557), .I3(n4147), .I4(n4148), .O(n4149));
  LUT3 #(.INIT(8'h96)) lut_n4150 (.I0(x564), .I1(x565), .I2(x566), .O(n4150));
  LUT5 #(.INIT(32'h96696996)) lut_n4151 (.I0(x555), .I1(x556), .I2(x557), .I3(n4147), .I4(n4148), .O(n4151));
  LUT5 #(.INIT(32'hFF969600)) lut_n4152 (.I0(x561), .I1(x562), .I2(x563), .I3(n4150), .I4(n4151), .O(n4152));
  LUT3 #(.INIT(8'h96)) lut_n4153 (.I0(n4127), .I1(n4130), .I2(n4131), .O(n4153));
  LUT3 #(.INIT(8'hE8)) lut_n4154 (.I0(n4149), .I1(n4152), .I2(n4153), .O(n4154));
  LUT3 #(.INIT(8'h96)) lut_n4155 (.I0(x570), .I1(x571), .I2(x572), .O(n4155));
  LUT5 #(.INIT(32'h96696996)) lut_n4156 (.I0(x561), .I1(x562), .I2(x563), .I3(n4150), .I4(n4151), .O(n4156));
  LUT5 #(.INIT(32'hFF969600)) lut_n4157 (.I0(x567), .I1(x568), .I2(x569), .I3(n4155), .I4(n4156), .O(n4157));
  LUT3 #(.INIT(8'h96)) lut_n4158 (.I0(x576), .I1(x577), .I2(x578), .O(n4158));
  LUT5 #(.INIT(32'h96696996)) lut_n4159 (.I0(x567), .I1(x568), .I2(x569), .I3(n4155), .I4(n4156), .O(n4159));
  LUT5 #(.INIT(32'hFF969600)) lut_n4160 (.I0(x573), .I1(x574), .I2(x575), .I3(n4158), .I4(n4159), .O(n4160));
  LUT3 #(.INIT(8'h96)) lut_n4161 (.I0(n4149), .I1(n4152), .I2(n4153), .O(n4161));
  LUT3 #(.INIT(8'hE8)) lut_n4162 (.I0(n4157), .I1(n4160), .I2(n4161), .O(n4162));
  LUT3 #(.INIT(8'h96)) lut_n4163 (.I0(n4124), .I1(n4132), .I2(n4133), .O(n4163));
  LUT3 #(.INIT(8'hE8)) lut_n4164 (.I0(n4154), .I1(n4162), .I2(n4163), .O(n4164));
  LUT3 #(.INIT(8'h96)) lut_n4165 (.I0(x582), .I1(x583), .I2(x584), .O(n4165));
  LUT5 #(.INIT(32'h96696996)) lut_n4166 (.I0(x573), .I1(x574), .I2(x575), .I3(n4158), .I4(n4159), .O(n4166));
  LUT5 #(.INIT(32'hFF969600)) lut_n4167 (.I0(x579), .I1(x580), .I2(x581), .I3(n4165), .I4(n4166), .O(n4167));
  LUT3 #(.INIT(8'h96)) lut_n4168 (.I0(x588), .I1(x589), .I2(x590), .O(n4168));
  LUT5 #(.INIT(32'h96696996)) lut_n4169 (.I0(x579), .I1(x580), .I2(x581), .I3(n4165), .I4(n4166), .O(n4169));
  LUT5 #(.INIT(32'hFF969600)) lut_n4170 (.I0(x585), .I1(x586), .I2(x587), .I3(n4168), .I4(n4169), .O(n4170));
  LUT3 #(.INIT(8'h96)) lut_n4171 (.I0(n4157), .I1(n4160), .I2(n4161), .O(n4171));
  LUT3 #(.INIT(8'hE8)) lut_n4172 (.I0(n4167), .I1(n4170), .I2(n4171), .O(n4172));
  LUT3 #(.INIT(8'h96)) lut_n4173 (.I0(x594), .I1(x595), .I2(x596), .O(n4173));
  LUT5 #(.INIT(32'h96696996)) lut_n4174 (.I0(x585), .I1(x586), .I2(x587), .I3(n4168), .I4(n4169), .O(n4174));
  LUT5 #(.INIT(32'hFF969600)) lut_n4175 (.I0(x591), .I1(x592), .I2(x593), .I3(n4173), .I4(n4174), .O(n4175));
  LUT3 #(.INIT(8'h96)) lut_n4176 (.I0(x600), .I1(x601), .I2(x602), .O(n4176));
  LUT5 #(.INIT(32'h96696996)) lut_n4177 (.I0(x591), .I1(x592), .I2(x593), .I3(n4173), .I4(n4174), .O(n4177));
  LUT5 #(.INIT(32'hFF969600)) lut_n4178 (.I0(x597), .I1(x598), .I2(x599), .I3(n4176), .I4(n4177), .O(n4178));
  LUT3 #(.INIT(8'h96)) lut_n4179 (.I0(n4167), .I1(n4170), .I2(n4171), .O(n4179));
  LUT3 #(.INIT(8'hE8)) lut_n4180 (.I0(n4175), .I1(n4178), .I2(n4179), .O(n4180));
  LUT3 #(.INIT(8'h96)) lut_n4181 (.I0(n4154), .I1(n4162), .I2(n4163), .O(n4181));
  LUT3 #(.INIT(8'hE8)) lut_n4182 (.I0(n4172), .I1(n4180), .I2(n4181), .O(n4182));
  LUT3 #(.INIT(8'h96)) lut_n4183 (.I0(n4116), .I1(n4134), .I2(n4135), .O(n4183));
  LUT3 #(.INIT(8'hE8)) lut_n4184 (.I0(n4164), .I1(n4182), .I2(n4183), .O(n4184));
  LUT3 #(.INIT(8'h96)) lut_n4185 (.I0(x606), .I1(x607), .I2(x608), .O(n4185));
  LUT5 #(.INIT(32'h96696996)) lut_n4186 (.I0(x597), .I1(x598), .I2(x599), .I3(n4176), .I4(n4177), .O(n4186));
  LUT5 #(.INIT(32'hFF969600)) lut_n4187 (.I0(x603), .I1(x604), .I2(x605), .I3(n4185), .I4(n4186), .O(n4187));
  LUT3 #(.INIT(8'h96)) lut_n4188 (.I0(x612), .I1(x613), .I2(x614), .O(n4188));
  LUT5 #(.INIT(32'h96696996)) lut_n4189 (.I0(x603), .I1(x604), .I2(x605), .I3(n4185), .I4(n4186), .O(n4189));
  LUT5 #(.INIT(32'hFF969600)) lut_n4190 (.I0(x609), .I1(x610), .I2(x611), .I3(n4188), .I4(n4189), .O(n4190));
  LUT3 #(.INIT(8'h96)) lut_n4191 (.I0(n4175), .I1(n4178), .I2(n4179), .O(n4191));
  LUT3 #(.INIT(8'hE8)) lut_n4192 (.I0(n4187), .I1(n4190), .I2(n4191), .O(n4192));
  LUT3 #(.INIT(8'h96)) lut_n4193 (.I0(x618), .I1(x619), .I2(x620), .O(n4193));
  LUT5 #(.INIT(32'h96696996)) lut_n4194 (.I0(x609), .I1(x610), .I2(x611), .I3(n4188), .I4(n4189), .O(n4194));
  LUT5 #(.INIT(32'hFF969600)) lut_n4195 (.I0(x615), .I1(x616), .I2(x617), .I3(n4193), .I4(n4194), .O(n4195));
  LUT3 #(.INIT(8'h96)) lut_n4196 (.I0(x624), .I1(x625), .I2(x626), .O(n4196));
  LUT5 #(.INIT(32'h96696996)) lut_n4197 (.I0(x615), .I1(x616), .I2(x617), .I3(n4193), .I4(n4194), .O(n4197));
  LUT5 #(.INIT(32'hFF969600)) lut_n4198 (.I0(x621), .I1(x622), .I2(x623), .I3(n4196), .I4(n4197), .O(n4198));
  LUT3 #(.INIT(8'h96)) lut_n4199 (.I0(n4187), .I1(n4190), .I2(n4191), .O(n4199));
  LUT3 #(.INIT(8'hE8)) lut_n4200 (.I0(n4195), .I1(n4198), .I2(n4199), .O(n4200));
  LUT3 #(.INIT(8'h96)) lut_n4201 (.I0(n4172), .I1(n4180), .I2(n4181), .O(n4201));
  LUT3 #(.INIT(8'hE8)) lut_n4202 (.I0(n4192), .I1(n4200), .I2(n4201), .O(n4202));
  LUT3 #(.INIT(8'h96)) lut_n4203 (.I0(x630), .I1(x631), .I2(x632), .O(n4203));
  LUT5 #(.INIT(32'h96696996)) lut_n4204 (.I0(x621), .I1(x622), .I2(x623), .I3(n4196), .I4(n4197), .O(n4204));
  LUT5 #(.INIT(32'hFF969600)) lut_n4205 (.I0(x627), .I1(x628), .I2(x629), .I3(n4203), .I4(n4204), .O(n4205));
  LUT3 #(.INIT(8'h96)) lut_n4206 (.I0(x636), .I1(x637), .I2(x638), .O(n4206));
  LUT5 #(.INIT(32'h96696996)) lut_n4207 (.I0(x627), .I1(x628), .I2(x629), .I3(n4203), .I4(n4204), .O(n4207));
  LUT5 #(.INIT(32'hFF969600)) lut_n4208 (.I0(x633), .I1(x634), .I2(x635), .I3(n4206), .I4(n4207), .O(n4208));
  LUT3 #(.INIT(8'h96)) lut_n4209 (.I0(n4195), .I1(n4198), .I2(n4199), .O(n4209));
  LUT3 #(.INIT(8'hE8)) lut_n4210 (.I0(n4205), .I1(n4208), .I2(n4209), .O(n4210));
  LUT3 #(.INIT(8'h96)) lut_n4211 (.I0(x642), .I1(x643), .I2(x644), .O(n4211));
  LUT5 #(.INIT(32'h96696996)) lut_n4212 (.I0(x633), .I1(x634), .I2(x635), .I3(n4206), .I4(n4207), .O(n4212));
  LUT5 #(.INIT(32'hFF969600)) lut_n4213 (.I0(x639), .I1(x640), .I2(x641), .I3(n4211), .I4(n4212), .O(n4213));
  LUT3 #(.INIT(8'h96)) lut_n4214 (.I0(x648), .I1(x649), .I2(x650), .O(n4214));
  LUT5 #(.INIT(32'h96696996)) lut_n4215 (.I0(x639), .I1(x640), .I2(x641), .I3(n4211), .I4(n4212), .O(n4215));
  LUT5 #(.INIT(32'hFF969600)) lut_n4216 (.I0(x645), .I1(x646), .I2(x647), .I3(n4214), .I4(n4215), .O(n4216));
  LUT3 #(.INIT(8'h96)) lut_n4217 (.I0(n4205), .I1(n4208), .I2(n4209), .O(n4217));
  LUT3 #(.INIT(8'hE8)) lut_n4218 (.I0(n4213), .I1(n4216), .I2(n4217), .O(n4218));
  LUT3 #(.INIT(8'h96)) lut_n4219 (.I0(n4192), .I1(n4200), .I2(n4201), .O(n4219));
  LUT3 #(.INIT(8'hE8)) lut_n4220 (.I0(n4210), .I1(n4218), .I2(n4219), .O(n4220));
  LUT3 #(.INIT(8'h96)) lut_n4221 (.I0(n4164), .I1(n4182), .I2(n4183), .O(n4221));
  LUT3 #(.INIT(8'hE8)) lut_n4222 (.I0(n4202), .I1(n4220), .I2(n4221), .O(n4222));
  LUT3 #(.INIT(8'h96)) lut_n4223 (.I0(n4098), .I1(n4136), .I2(n4137), .O(n4223));
  LUT3 #(.INIT(8'hE8)) lut_n4224 (.I0(n4184), .I1(n4222), .I2(n4223), .O(n4224));
  LUT3 #(.INIT(8'h96)) lut_n4225 (.I0(x654), .I1(x655), .I2(x656), .O(n4225));
  LUT5 #(.INIT(32'h96696996)) lut_n4226 (.I0(x645), .I1(x646), .I2(x647), .I3(n4214), .I4(n4215), .O(n4226));
  LUT5 #(.INIT(32'hFF969600)) lut_n4227 (.I0(x651), .I1(x652), .I2(x653), .I3(n4225), .I4(n4226), .O(n4227));
  LUT3 #(.INIT(8'h96)) lut_n4228 (.I0(x660), .I1(x661), .I2(x662), .O(n4228));
  LUT5 #(.INIT(32'h96696996)) lut_n4229 (.I0(x651), .I1(x652), .I2(x653), .I3(n4225), .I4(n4226), .O(n4229));
  LUT5 #(.INIT(32'hFF969600)) lut_n4230 (.I0(x657), .I1(x658), .I2(x659), .I3(n4228), .I4(n4229), .O(n4230));
  LUT3 #(.INIT(8'h96)) lut_n4231 (.I0(n4213), .I1(n4216), .I2(n4217), .O(n4231));
  LUT3 #(.INIT(8'hE8)) lut_n4232 (.I0(n4227), .I1(n4230), .I2(n4231), .O(n4232));
  LUT3 #(.INIT(8'h96)) lut_n4233 (.I0(x666), .I1(x667), .I2(x668), .O(n4233));
  LUT5 #(.INIT(32'h96696996)) lut_n4234 (.I0(x657), .I1(x658), .I2(x659), .I3(n4228), .I4(n4229), .O(n4234));
  LUT5 #(.INIT(32'hFF969600)) lut_n4235 (.I0(x663), .I1(x664), .I2(x665), .I3(n4233), .I4(n4234), .O(n4235));
  LUT3 #(.INIT(8'h96)) lut_n4236 (.I0(x672), .I1(x673), .I2(x674), .O(n4236));
  LUT5 #(.INIT(32'h96696996)) lut_n4237 (.I0(x663), .I1(x664), .I2(x665), .I3(n4233), .I4(n4234), .O(n4237));
  LUT5 #(.INIT(32'hFF969600)) lut_n4238 (.I0(x669), .I1(x670), .I2(x671), .I3(n4236), .I4(n4237), .O(n4238));
  LUT3 #(.INIT(8'h96)) lut_n4239 (.I0(n4227), .I1(n4230), .I2(n4231), .O(n4239));
  LUT3 #(.INIT(8'hE8)) lut_n4240 (.I0(n4235), .I1(n4238), .I2(n4239), .O(n4240));
  LUT3 #(.INIT(8'h96)) lut_n4241 (.I0(n4210), .I1(n4218), .I2(n4219), .O(n4241));
  LUT3 #(.INIT(8'hE8)) lut_n4242 (.I0(n4232), .I1(n4240), .I2(n4241), .O(n4242));
  LUT3 #(.INIT(8'h96)) lut_n4243 (.I0(x678), .I1(x679), .I2(x680), .O(n4243));
  LUT5 #(.INIT(32'h96696996)) lut_n4244 (.I0(x669), .I1(x670), .I2(x671), .I3(n4236), .I4(n4237), .O(n4244));
  LUT5 #(.INIT(32'hFF969600)) lut_n4245 (.I0(x675), .I1(x676), .I2(x677), .I3(n4243), .I4(n4244), .O(n4245));
  LUT3 #(.INIT(8'h96)) lut_n4246 (.I0(x684), .I1(x685), .I2(x686), .O(n4246));
  LUT5 #(.INIT(32'h96696996)) lut_n4247 (.I0(x675), .I1(x676), .I2(x677), .I3(n4243), .I4(n4244), .O(n4247));
  LUT5 #(.INIT(32'hFF969600)) lut_n4248 (.I0(x681), .I1(x682), .I2(x683), .I3(n4246), .I4(n4247), .O(n4248));
  LUT3 #(.INIT(8'h96)) lut_n4249 (.I0(n4235), .I1(n4238), .I2(n4239), .O(n4249));
  LUT3 #(.INIT(8'hE8)) lut_n4250 (.I0(n4245), .I1(n4248), .I2(n4249), .O(n4250));
  LUT3 #(.INIT(8'h96)) lut_n4251 (.I0(x690), .I1(x691), .I2(x692), .O(n4251));
  LUT5 #(.INIT(32'h96696996)) lut_n4252 (.I0(x681), .I1(x682), .I2(x683), .I3(n4246), .I4(n4247), .O(n4252));
  LUT5 #(.INIT(32'hFF969600)) lut_n4253 (.I0(x687), .I1(x688), .I2(x689), .I3(n4251), .I4(n4252), .O(n4253));
  LUT3 #(.INIT(8'h96)) lut_n4254 (.I0(x696), .I1(x697), .I2(x698), .O(n4254));
  LUT5 #(.INIT(32'h96696996)) lut_n4255 (.I0(x687), .I1(x688), .I2(x689), .I3(n4251), .I4(n4252), .O(n4255));
  LUT5 #(.INIT(32'hFF969600)) lut_n4256 (.I0(x693), .I1(x694), .I2(x695), .I3(n4254), .I4(n4255), .O(n4256));
  LUT3 #(.INIT(8'h96)) lut_n4257 (.I0(n4245), .I1(n4248), .I2(n4249), .O(n4257));
  LUT3 #(.INIT(8'hE8)) lut_n4258 (.I0(n4253), .I1(n4256), .I2(n4257), .O(n4258));
  LUT3 #(.INIT(8'h96)) lut_n4259 (.I0(n4232), .I1(n4240), .I2(n4241), .O(n4259));
  LUT3 #(.INIT(8'hE8)) lut_n4260 (.I0(n4250), .I1(n4258), .I2(n4259), .O(n4260));
  LUT3 #(.INIT(8'h96)) lut_n4261 (.I0(n4202), .I1(n4220), .I2(n4221), .O(n4261));
  LUT3 #(.INIT(8'hE8)) lut_n4262 (.I0(n4242), .I1(n4260), .I2(n4261), .O(n4262));
  LUT3 #(.INIT(8'h96)) lut_n4263 (.I0(x702), .I1(x703), .I2(x704), .O(n4263));
  LUT5 #(.INIT(32'h96696996)) lut_n4264 (.I0(x693), .I1(x694), .I2(x695), .I3(n4254), .I4(n4255), .O(n4264));
  LUT5 #(.INIT(32'hFF969600)) lut_n4265 (.I0(x699), .I1(x700), .I2(x701), .I3(n4263), .I4(n4264), .O(n4265));
  LUT3 #(.INIT(8'h96)) lut_n4266 (.I0(x708), .I1(x709), .I2(x710), .O(n4266));
  LUT5 #(.INIT(32'h96696996)) lut_n4267 (.I0(x699), .I1(x700), .I2(x701), .I3(n4263), .I4(n4264), .O(n4267));
  LUT5 #(.INIT(32'hFF969600)) lut_n4268 (.I0(x705), .I1(x706), .I2(x707), .I3(n4266), .I4(n4267), .O(n4268));
  LUT3 #(.INIT(8'h96)) lut_n4269 (.I0(n4253), .I1(n4256), .I2(n4257), .O(n4269));
  LUT3 #(.INIT(8'hE8)) lut_n4270 (.I0(n4265), .I1(n4268), .I2(n4269), .O(n4270));
  LUT3 #(.INIT(8'h96)) lut_n4271 (.I0(x714), .I1(x715), .I2(x716), .O(n4271));
  LUT5 #(.INIT(32'h96696996)) lut_n4272 (.I0(x705), .I1(x706), .I2(x707), .I3(n4266), .I4(n4267), .O(n4272));
  LUT5 #(.INIT(32'hFF969600)) lut_n4273 (.I0(x711), .I1(x712), .I2(x713), .I3(n4271), .I4(n4272), .O(n4273));
  LUT3 #(.INIT(8'h96)) lut_n4274 (.I0(x720), .I1(x721), .I2(x722), .O(n4274));
  LUT5 #(.INIT(32'h96696996)) lut_n4275 (.I0(x711), .I1(x712), .I2(x713), .I3(n4271), .I4(n4272), .O(n4275));
  LUT5 #(.INIT(32'hFF969600)) lut_n4276 (.I0(x717), .I1(x718), .I2(x719), .I3(n4274), .I4(n4275), .O(n4276));
  LUT3 #(.INIT(8'h96)) lut_n4277 (.I0(n4265), .I1(n4268), .I2(n4269), .O(n4277));
  LUT3 #(.INIT(8'hE8)) lut_n4278 (.I0(n4273), .I1(n4276), .I2(n4277), .O(n4278));
  LUT3 #(.INIT(8'h96)) lut_n4279 (.I0(n4250), .I1(n4258), .I2(n4259), .O(n4279));
  LUT3 #(.INIT(8'hE8)) lut_n4280 (.I0(n4270), .I1(n4278), .I2(n4279), .O(n4280));
  LUT3 #(.INIT(8'h96)) lut_n4281 (.I0(x726), .I1(x727), .I2(x728), .O(n4281));
  LUT5 #(.INIT(32'h96696996)) lut_n4282 (.I0(x717), .I1(x718), .I2(x719), .I3(n4274), .I4(n4275), .O(n4282));
  LUT5 #(.INIT(32'hFF969600)) lut_n4283 (.I0(x723), .I1(x724), .I2(x725), .I3(n4281), .I4(n4282), .O(n4283));
  LUT3 #(.INIT(8'h96)) lut_n4284 (.I0(x732), .I1(x733), .I2(x734), .O(n4284));
  LUT5 #(.INIT(32'h96696996)) lut_n4285 (.I0(x723), .I1(x724), .I2(x725), .I3(n4281), .I4(n4282), .O(n4285));
  LUT5 #(.INIT(32'hFF969600)) lut_n4286 (.I0(x729), .I1(x730), .I2(x731), .I3(n4284), .I4(n4285), .O(n4286));
  LUT3 #(.INIT(8'h96)) lut_n4287 (.I0(n4273), .I1(n4276), .I2(n4277), .O(n4287));
  LUT3 #(.INIT(8'hE8)) lut_n4288 (.I0(n4283), .I1(n4286), .I2(n4287), .O(n4288));
  LUT3 #(.INIT(8'h96)) lut_n4289 (.I0(x738), .I1(x739), .I2(x740), .O(n4289));
  LUT5 #(.INIT(32'h96696996)) lut_n4290 (.I0(x729), .I1(x730), .I2(x731), .I3(n4284), .I4(n4285), .O(n4290));
  LUT5 #(.INIT(32'hFF969600)) lut_n4291 (.I0(x735), .I1(x736), .I2(x737), .I3(n4289), .I4(n4290), .O(n4291));
  LUT3 #(.INIT(8'h96)) lut_n4292 (.I0(x744), .I1(x745), .I2(x746), .O(n4292));
  LUT5 #(.INIT(32'h96696996)) lut_n4293 (.I0(x735), .I1(x736), .I2(x737), .I3(n4289), .I4(n4290), .O(n4293));
  LUT5 #(.INIT(32'hFF969600)) lut_n4294 (.I0(x741), .I1(x742), .I2(x743), .I3(n4292), .I4(n4293), .O(n4294));
  LUT3 #(.INIT(8'h96)) lut_n4295 (.I0(n4283), .I1(n4286), .I2(n4287), .O(n4295));
  LUT3 #(.INIT(8'hE8)) lut_n4296 (.I0(n4291), .I1(n4294), .I2(n4295), .O(n4296));
  LUT3 #(.INIT(8'h96)) lut_n4297 (.I0(n4270), .I1(n4278), .I2(n4279), .O(n4297));
  LUT3 #(.INIT(8'hE8)) lut_n4298 (.I0(n4288), .I1(n4296), .I2(n4297), .O(n4298));
  LUT3 #(.INIT(8'h96)) lut_n4299 (.I0(n4242), .I1(n4260), .I2(n4261), .O(n4299));
  LUT3 #(.INIT(8'hE8)) lut_n4300 (.I0(n4280), .I1(n4298), .I2(n4299), .O(n4300));
  LUT3 #(.INIT(8'h96)) lut_n4301 (.I0(n4184), .I1(n4222), .I2(n4223), .O(n4301));
  LUT3 #(.INIT(8'hE8)) lut_n4302 (.I0(n4262), .I1(n4300), .I2(n4301), .O(n4302));
  LUT3 #(.INIT(8'h96)) lut_n4303 (.I0(n4060), .I1(n4138), .I2(n4139), .O(n4303));
  LUT3 #(.INIT(8'hE8)) lut_n4304 (.I0(n4224), .I1(n4302), .I2(n4303), .O(n4304));
  LUT3 #(.INIT(8'h96)) lut_n4305 (.I0(x750), .I1(x751), .I2(x752), .O(n4305));
  LUT5 #(.INIT(32'h96696996)) lut_n4306 (.I0(x741), .I1(x742), .I2(x743), .I3(n4292), .I4(n4293), .O(n4306));
  LUT5 #(.INIT(32'hFF969600)) lut_n4307 (.I0(x747), .I1(x748), .I2(x749), .I3(n4305), .I4(n4306), .O(n4307));
  LUT3 #(.INIT(8'h96)) lut_n4308 (.I0(x756), .I1(x757), .I2(x758), .O(n4308));
  LUT5 #(.INIT(32'h96696996)) lut_n4309 (.I0(x747), .I1(x748), .I2(x749), .I3(n4305), .I4(n4306), .O(n4309));
  LUT5 #(.INIT(32'hFF969600)) lut_n4310 (.I0(x753), .I1(x754), .I2(x755), .I3(n4308), .I4(n4309), .O(n4310));
  LUT3 #(.INIT(8'h96)) lut_n4311 (.I0(n4291), .I1(n4294), .I2(n4295), .O(n4311));
  LUT3 #(.INIT(8'hE8)) lut_n4312 (.I0(n4307), .I1(n4310), .I2(n4311), .O(n4312));
  LUT3 #(.INIT(8'h96)) lut_n4313 (.I0(x762), .I1(x763), .I2(x764), .O(n4313));
  LUT5 #(.INIT(32'h96696996)) lut_n4314 (.I0(x753), .I1(x754), .I2(x755), .I3(n4308), .I4(n4309), .O(n4314));
  LUT5 #(.INIT(32'hFF969600)) lut_n4315 (.I0(x759), .I1(x760), .I2(x761), .I3(n4313), .I4(n4314), .O(n4315));
  LUT3 #(.INIT(8'h96)) lut_n4316 (.I0(x768), .I1(x769), .I2(x770), .O(n4316));
  LUT5 #(.INIT(32'h96696996)) lut_n4317 (.I0(x759), .I1(x760), .I2(x761), .I3(n4313), .I4(n4314), .O(n4317));
  LUT5 #(.INIT(32'hFF969600)) lut_n4318 (.I0(x765), .I1(x766), .I2(x767), .I3(n4316), .I4(n4317), .O(n4318));
  LUT3 #(.INIT(8'h96)) lut_n4319 (.I0(n4307), .I1(n4310), .I2(n4311), .O(n4319));
  LUT3 #(.INIT(8'hE8)) lut_n4320 (.I0(n4315), .I1(n4318), .I2(n4319), .O(n4320));
  LUT3 #(.INIT(8'h96)) lut_n4321 (.I0(n4288), .I1(n4296), .I2(n4297), .O(n4321));
  LUT3 #(.INIT(8'hE8)) lut_n4322 (.I0(n4312), .I1(n4320), .I2(n4321), .O(n4322));
  LUT3 #(.INIT(8'h96)) lut_n4323 (.I0(x774), .I1(x775), .I2(x776), .O(n4323));
  LUT5 #(.INIT(32'h96696996)) lut_n4324 (.I0(x765), .I1(x766), .I2(x767), .I3(n4316), .I4(n4317), .O(n4324));
  LUT5 #(.INIT(32'hFF969600)) lut_n4325 (.I0(x771), .I1(x772), .I2(x773), .I3(n4323), .I4(n4324), .O(n4325));
  LUT3 #(.INIT(8'h96)) lut_n4326 (.I0(x780), .I1(x781), .I2(x782), .O(n4326));
  LUT5 #(.INIT(32'h96696996)) lut_n4327 (.I0(x771), .I1(x772), .I2(x773), .I3(n4323), .I4(n4324), .O(n4327));
  LUT5 #(.INIT(32'hFF969600)) lut_n4328 (.I0(x777), .I1(x778), .I2(x779), .I3(n4326), .I4(n4327), .O(n4328));
  LUT3 #(.INIT(8'h96)) lut_n4329 (.I0(n4315), .I1(n4318), .I2(n4319), .O(n4329));
  LUT3 #(.INIT(8'hE8)) lut_n4330 (.I0(n4325), .I1(n4328), .I2(n4329), .O(n4330));
  LUT3 #(.INIT(8'h96)) lut_n4331 (.I0(x786), .I1(x787), .I2(x788), .O(n4331));
  LUT5 #(.INIT(32'h96696996)) lut_n4332 (.I0(x777), .I1(x778), .I2(x779), .I3(n4326), .I4(n4327), .O(n4332));
  LUT5 #(.INIT(32'hFF969600)) lut_n4333 (.I0(x783), .I1(x784), .I2(x785), .I3(n4331), .I4(n4332), .O(n4333));
  LUT3 #(.INIT(8'h96)) lut_n4334 (.I0(x792), .I1(x793), .I2(x794), .O(n4334));
  LUT5 #(.INIT(32'h96696996)) lut_n4335 (.I0(x783), .I1(x784), .I2(x785), .I3(n4331), .I4(n4332), .O(n4335));
  LUT5 #(.INIT(32'hFF969600)) lut_n4336 (.I0(x789), .I1(x790), .I2(x791), .I3(n4334), .I4(n4335), .O(n4336));
  LUT3 #(.INIT(8'h96)) lut_n4337 (.I0(n4325), .I1(n4328), .I2(n4329), .O(n4337));
  LUT3 #(.INIT(8'hE8)) lut_n4338 (.I0(n4333), .I1(n4336), .I2(n4337), .O(n4338));
  LUT3 #(.INIT(8'h96)) lut_n4339 (.I0(n4312), .I1(n4320), .I2(n4321), .O(n4339));
  LUT3 #(.INIT(8'hE8)) lut_n4340 (.I0(n4330), .I1(n4338), .I2(n4339), .O(n4340));
  LUT3 #(.INIT(8'h96)) lut_n4341 (.I0(n4280), .I1(n4298), .I2(n4299), .O(n4341));
  LUT3 #(.INIT(8'hE8)) lut_n4342 (.I0(n4322), .I1(n4340), .I2(n4341), .O(n4342));
  LUT3 #(.INIT(8'h96)) lut_n4343 (.I0(x798), .I1(x799), .I2(x800), .O(n4343));
  LUT5 #(.INIT(32'h96696996)) lut_n4344 (.I0(x789), .I1(x790), .I2(x791), .I3(n4334), .I4(n4335), .O(n4344));
  LUT5 #(.INIT(32'hFF969600)) lut_n4345 (.I0(x795), .I1(x796), .I2(x797), .I3(n4343), .I4(n4344), .O(n4345));
  LUT3 #(.INIT(8'h96)) lut_n4346 (.I0(x804), .I1(x805), .I2(x806), .O(n4346));
  LUT5 #(.INIT(32'h96696996)) lut_n4347 (.I0(x795), .I1(x796), .I2(x797), .I3(n4343), .I4(n4344), .O(n4347));
  LUT5 #(.INIT(32'hFF969600)) lut_n4348 (.I0(x801), .I1(x802), .I2(x803), .I3(n4346), .I4(n4347), .O(n4348));
  LUT3 #(.INIT(8'h96)) lut_n4349 (.I0(n4333), .I1(n4336), .I2(n4337), .O(n4349));
  LUT3 #(.INIT(8'hE8)) lut_n4350 (.I0(n4345), .I1(n4348), .I2(n4349), .O(n4350));
  LUT3 #(.INIT(8'h96)) lut_n4351 (.I0(x810), .I1(x811), .I2(x812), .O(n4351));
  LUT5 #(.INIT(32'h96696996)) lut_n4352 (.I0(x801), .I1(x802), .I2(x803), .I3(n4346), .I4(n4347), .O(n4352));
  LUT5 #(.INIT(32'hFF969600)) lut_n4353 (.I0(x807), .I1(x808), .I2(x809), .I3(n4351), .I4(n4352), .O(n4353));
  LUT3 #(.INIT(8'h96)) lut_n4354 (.I0(x816), .I1(x817), .I2(x818), .O(n4354));
  LUT5 #(.INIT(32'h96696996)) lut_n4355 (.I0(x807), .I1(x808), .I2(x809), .I3(n4351), .I4(n4352), .O(n4355));
  LUT5 #(.INIT(32'hFF969600)) lut_n4356 (.I0(x813), .I1(x814), .I2(x815), .I3(n4354), .I4(n4355), .O(n4356));
  LUT3 #(.INIT(8'h96)) lut_n4357 (.I0(n4345), .I1(n4348), .I2(n4349), .O(n4357));
  LUT3 #(.INIT(8'hE8)) lut_n4358 (.I0(n4353), .I1(n4356), .I2(n4357), .O(n4358));
  LUT3 #(.INIT(8'h96)) lut_n4359 (.I0(n4330), .I1(n4338), .I2(n4339), .O(n4359));
  LUT3 #(.INIT(8'hE8)) lut_n4360 (.I0(n4350), .I1(n4358), .I2(n4359), .O(n4360));
  LUT3 #(.INIT(8'h96)) lut_n4361 (.I0(x822), .I1(x823), .I2(x824), .O(n4361));
  LUT5 #(.INIT(32'h96696996)) lut_n4362 (.I0(x813), .I1(x814), .I2(x815), .I3(n4354), .I4(n4355), .O(n4362));
  LUT5 #(.INIT(32'hFF969600)) lut_n4363 (.I0(x819), .I1(x820), .I2(x821), .I3(n4361), .I4(n4362), .O(n4363));
  LUT3 #(.INIT(8'h96)) lut_n4364 (.I0(x828), .I1(x829), .I2(x830), .O(n4364));
  LUT5 #(.INIT(32'h96696996)) lut_n4365 (.I0(x819), .I1(x820), .I2(x821), .I3(n4361), .I4(n4362), .O(n4365));
  LUT5 #(.INIT(32'hFF969600)) lut_n4366 (.I0(x825), .I1(x826), .I2(x827), .I3(n4364), .I4(n4365), .O(n4366));
  LUT3 #(.INIT(8'h96)) lut_n4367 (.I0(n4353), .I1(n4356), .I2(n4357), .O(n4367));
  LUT3 #(.INIT(8'hE8)) lut_n4368 (.I0(n4363), .I1(n4366), .I2(n4367), .O(n4368));
  LUT3 #(.INIT(8'h96)) lut_n4369 (.I0(x834), .I1(x835), .I2(x836), .O(n4369));
  LUT5 #(.INIT(32'h96696996)) lut_n4370 (.I0(x825), .I1(x826), .I2(x827), .I3(n4364), .I4(n4365), .O(n4370));
  LUT5 #(.INIT(32'hFF969600)) lut_n4371 (.I0(x831), .I1(x832), .I2(x833), .I3(n4369), .I4(n4370), .O(n4371));
  LUT3 #(.INIT(8'h96)) lut_n4372 (.I0(x840), .I1(x841), .I2(x842), .O(n4372));
  LUT5 #(.INIT(32'h96696996)) lut_n4373 (.I0(x831), .I1(x832), .I2(x833), .I3(n4369), .I4(n4370), .O(n4373));
  LUT5 #(.INIT(32'hFF969600)) lut_n4374 (.I0(x837), .I1(x838), .I2(x839), .I3(n4372), .I4(n4373), .O(n4374));
  LUT3 #(.INIT(8'h96)) lut_n4375 (.I0(n4363), .I1(n4366), .I2(n4367), .O(n4375));
  LUT3 #(.INIT(8'hE8)) lut_n4376 (.I0(n4371), .I1(n4374), .I2(n4375), .O(n4376));
  LUT3 #(.INIT(8'h96)) lut_n4377 (.I0(n4350), .I1(n4358), .I2(n4359), .O(n4377));
  LUT3 #(.INIT(8'hE8)) lut_n4378 (.I0(n4368), .I1(n4376), .I2(n4377), .O(n4378));
  LUT3 #(.INIT(8'h96)) lut_n4379 (.I0(n4322), .I1(n4340), .I2(n4341), .O(n4379));
  LUT3 #(.INIT(8'hE8)) lut_n4380 (.I0(n4360), .I1(n4378), .I2(n4379), .O(n4380));
  LUT3 #(.INIT(8'h96)) lut_n4381 (.I0(n4262), .I1(n4300), .I2(n4301), .O(n4381));
  LUT3 #(.INIT(8'hE8)) lut_n4382 (.I0(n4342), .I1(n4380), .I2(n4381), .O(n4382));
  LUT3 #(.INIT(8'h96)) lut_n4383 (.I0(x846), .I1(x847), .I2(x848), .O(n4383));
  LUT5 #(.INIT(32'h96696996)) lut_n4384 (.I0(x837), .I1(x838), .I2(x839), .I3(n4372), .I4(n4373), .O(n4384));
  LUT5 #(.INIT(32'hFF969600)) lut_n4385 (.I0(x843), .I1(x844), .I2(x845), .I3(n4383), .I4(n4384), .O(n4385));
  LUT3 #(.INIT(8'h96)) lut_n4386 (.I0(x852), .I1(x853), .I2(x854), .O(n4386));
  LUT5 #(.INIT(32'h96696996)) lut_n4387 (.I0(x843), .I1(x844), .I2(x845), .I3(n4383), .I4(n4384), .O(n4387));
  LUT5 #(.INIT(32'hFF969600)) lut_n4388 (.I0(x849), .I1(x850), .I2(x851), .I3(n4386), .I4(n4387), .O(n4388));
  LUT3 #(.INIT(8'h96)) lut_n4389 (.I0(n4371), .I1(n4374), .I2(n4375), .O(n4389));
  LUT3 #(.INIT(8'hE8)) lut_n4390 (.I0(n4385), .I1(n4388), .I2(n4389), .O(n4390));
  LUT3 #(.INIT(8'h96)) lut_n4391 (.I0(x858), .I1(x859), .I2(x860), .O(n4391));
  LUT5 #(.INIT(32'h96696996)) lut_n4392 (.I0(x849), .I1(x850), .I2(x851), .I3(n4386), .I4(n4387), .O(n4392));
  LUT5 #(.INIT(32'hFF969600)) lut_n4393 (.I0(x855), .I1(x856), .I2(x857), .I3(n4391), .I4(n4392), .O(n4393));
  LUT3 #(.INIT(8'h96)) lut_n4394 (.I0(x864), .I1(x865), .I2(x866), .O(n4394));
  LUT5 #(.INIT(32'h96696996)) lut_n4395 (.I0(x855), .I1(x856), .I2(x857), .I3(n4391), .I4(n4392), .O(n4395));
  LUT5 #(.INIT(32'hFF969600)) lut_n4396 (.I0(x861), .I1(x862), .I2(x863), .I3(n4394), .I4(n4395), .O(n4396));
  LUT3 #(.INIT(8'h96)) lut_n4397 (.I0(n4385), .I1(n4388), .I2(n4389), .O(n4397));
  LUT3 #(.INIT(8'hE8)) lut_n4398 (.I0(n4393), .I1(n4396), .I2(n4397), .O(n4398));
  LUT3 #(.INIT(8'h96)) lut_n4399 (.I0(n4368), .I1(n4376), .I2(n4377), .O(n4399));
  LUT3 #(.INIT(8'hE8)) lut_n4400 (.I0(n4390), .I1(n4398), .I2(n4399), .O(n4400));
  LUT3 #(.INIT(8'h96)) lut_n4401 (.I0(x870), .I1(x871), .I2(x872), .O(n4401));
  LUT5 #(.INIT(32'h96696996)) lut_n4402 (.I0(x861), .I1(x862), .I2(x863), .I3(n4394), .I4(n4395), .O(n4402));
  LUT5 #(.INIT(32'hFF969600)) lut_n4403 (.I0(x867), .I1(x868), .I2(x869), .I3(n4401), .I4(n4402), .O(n4403));
  LUT3 #(.INIT(8'h96)) lut_n4404 (.I0(x876), .I1(x877), .I2(x878), .O(n4404));
  LUT5 #(.INIT(32'h96696996)) lut_n4405 (.I0(x867), .I1(x868), .I2(x869), .I3(n4401), .I4(n4402), .O(n4405));
  LUT5 #(.INIT(32'hFF969600)) lut_n4406 (.I0(x873), .I1(x874), .I2(x875), .I3(n4404), .I4(n4405), .O(n4406));
  LUT3 #(.INIT(8'h96)) lut_n4407 (.I0(n4393), .I1(n4396), .I2(n4397), .O(n4407));
  LUT3 #(.INIT(8'hE8)) lut_n4408 (.I0(n4403), .I1(n4406), .I2(n4407), .O(n4408));
  LUT3 #(.INIT(8'h96)) lut_n4409 (.I0(x882), .I1(x883), .I2(x884), .O(n4409));
  LUT5 #(.INIT(32'h96696996)) lut_n4410 (.I0(x873), .I1(x874), .I2(x875), .I3(n4404), .I4(n4405), .O(n4410));
  LUT5 #(.INIT(32'hFF969600)) lut_n4411 (.I0(x879), .I1(x880), .I2(x881), .I3(n4409), .I4(n4410), .O(n4411));
  LUT3 #(.INIT(8'h96)) lut_n4412 (.I0(x888), .I1(x889), .I2(x890), .O(n4412));
  LUT5 #(.INIT(32'h96696996)) lut_n4413 (.I0(x879), .I1(x880), .I2(x881), .I3(n4409), .I4(n4410), .O(n4413));
  LUT5 #(.INIT(32'hFF969600)) lut_n4414 (.I0(x885), .I1(x886), .I2(x887), .I3(n4412), .I4(n4413), .O(n4414));
  LUT3 #(.INIT(8'h96)) lut_n4415 (.I0(n4403), .I1(n4406), .I2(n4407), .O(n4415));
  LUT3 #(.INIT(8'hE8)) lut_n4416 (.I0(n4411), .I1(n4414), .I2(n4415), .O(n4416));
  LUT3 #(.INIT(8'h96)) lut_n4417 (.I0(n4390), .I1(n4398), .I2(n4399), .O(n4417));
  LUT3 #(.INIT(8'hE8)) lut_n4418 (.I0(n4408), .I1(n4416), .I2(n4417), .O(n4418));
  LUT3 #(.INIT(8'h96)) lut_n4419 (.I0(n4360), .I1(n4378), .I2(n4379), .O(n4419));
  LUT3 #(.INIT(8'hE8)) lut_n4420 (.I0(n4400), .I1(n4418), .I2(n4419), .O(n4420));
  LUT3 #(.INIT(8'h96)) lut_n4421 (.I0(x894), .I1(x895), .I2(x896), .O(n4421));
  LUT5 #(.INIT(32'h96696996)) lut_n4422 (.I0(x885), .I1(x886), .I2(x887), .I3(n4412), .I4(n4413), .O(n4422));
  LUT5 #(.INIT(32'hFF969600)) lut_n4423 (.I0(x891), .I1(x892), .I2(x893), .I3(n4421), .I4(n4422), .O(n4423));
  LUT3 #(.INIT(8'h96)) lut_n4424 (.I0(x900), .I1(x901), .I2(x902), .O(n4424));
  LUT5 #(.INIT(32'h96696996)) lut_n4425 (.I0(x891), .I1(x892), .I2(x893), .I3(n4421), .I4(n4422), .O(n4425));
  LUT5 #(.INIT(32'hFF969600)) lut_n4426 (.I0(x897), .I1(x898), .I2(x899), .I3(n4424), .I4(n4425), .O(n4426));
  LUT3 #(.INIT(8'h96)) lut_n4427 (.I0(n4411), .I1(n4414), .I2(n4415), .O(n4427));
  LUT3 #(.INIT(8'hE8)) lut_n4428 (.I0(n4423), .I1(n4426), .I2(n4427), .O(n4428));
  LUT3 #(.INIT(8'h96)) lut_n4429 (.I0(x906), .I1(x907), .I2(x908), .O(n4429));
  LUT5 #(.INIT(32'h96696996)) lut_n4430 (.I0(x897), .I1(x898), .I2(x899), .I3(n4424), .I4(n4425), .O(n4430));
  LUT5 #(.INIT(32'hFF969600)) lut_n4431 (.I0(x903), .I1(x904), .I2(x905), .I3(n4429), .I4(n4430), .O(n4431));
  LUT3 #(.INIT(8'h96)) lut_n4432 (.I0(x912), .I1(x913), .I2(x914), .O(n4432));
  LUT5 #(.INIT(32'h96696996)) lut_n4433 (.I0(x903), .I1(x904), .I2(x905), .I3(n4429), .I4(n4430), .O(n4433));
  LUT5 #(.INIT(32'hFF969600)) lut_n4434 (.I0(x909), .I1(x910), .I2(x911), .I3(n4432), .I4(n4433), .O(n4434));
  LUT3 #(.INIT(8'h96)) lut_n4435 (.I0(n4423), .I1(n4426), .I2(n4427), .O(n4435));
  LUT3 #(.INIT(8'hE8)) lut_n4436 (.I0(n4431), .I1(n4434), .I2(n4435), .O(n4436));
  LUT3 #(.INIT(8'h96)) lut_n4437 (.I0(n4408), .I1(n4416), .I2(n4417), .O(n4437));
  LUT3 #(.INIT(8'hE8)) lut_n4438 (.I0(n4428), .I1(n4436), .I2(n4437), .O(n4438));
  LUT3 #(.INIT(8'h96)) lut_n4439 (.I0(x918), .I1(x919), .I2(x920), .O(n4439));
  LUT5 #(.INIT(32'h96696996)) lut_n4440 (.I0(x909), .I1(x910), .I2(x911), .I3(n4432), .I4(n4433), .O(n4440));
  LUT5 #(.INIT(32'hFF969600)) lut_n4441 (.I0(x915), .I1(x916), .I2(x917), .I3(n4439), .I4(n4440), .O(n4441));
  LUT3 #(.INIT(8'h96)) lut_n4442 (.I0(x924), .I1(x925), .I2(x926), .O(n4442));
  LUT5 #(.INIT(32'h96696996)) lut_n4443 (.I0(x915), .I1(x916), .I2(x917), .I3(n4439), .I4(n4440), .O(n4443));
  LUT5 #(.INIT(32'hFF969600)) lut_n4444 (.I0(x921), .I1(x922), .I2(x923), .I3(n4442), .I4(n4443), .O(n4444));
  LUT3 #(.INIT(8'h96)) lut_n4445 (.I0(n4431), .I1(n4434), .I2(n4435), .O(n4445));
  LUT3 #(.INIT(8'hE8)) lut_n4446 (.I0(n4441), .I1(n4444), .I2(n4445), .O(n4446));
  LUT3 #(.INIT(8'h96)) lut_n4447 (.I0(x930), .I1(x931), .I2(x932), .O(n4447));
  LUT5 #(.INIT(32'h96696996)) lut_n4448 (.I0(x921), .I1(x922), .I2(x923), .I3(n4442), .I4(n4443), .O(n4448));
  LUT5 #(.INIT(32'hFF969600)) lut_n4449 (.I0(x927), .I1(x928), .I2(x929), .I3(n4447), .I4(n4448), .O(n4449));
  LUT3 #(.INIT(8'h96)) lut_n4450 (.I0(x936), .I1(x937), .I2(x938), .O(n4450));
  LUT5 #(.INIT(32'h96696996)) lut_n4451 (.I0(x927), .I1(x928), .I2(x929), .I3(n4447), .I4(n4448), .O(n4451));
  LUT5 #(.INIT(32'hFF969600)) lut_n4452 (.I0(x933), .I1(x934), .I2(x935), .I3(n4450), .I4(n4451), .O(n4452));
  LUT3 #(.INIT(8'h96)) lut_n4453 (.I0(n4441), .I1(n4444), .I2(n4445), .O(n4453));
  LUT3 #(.INIT(8'hE8)) lut_n4454 (.I0(n4449), .I1(n4452), .I2(n4453), .O(n4454));
  LUT3 #(.INIT(8'h96)) lut_n4455 (.I0(n4428), .I1(n4436), .I2(n4437), .O(n4455));
  LUT3 #(.INIT(8'hE8)) lut_n4456 (.I0(n4446), .I1(n4454), .I2(n4455), .O(n4456));
  LUT3 #(.INIT(8'h96)) lut_n4457 (.I0(n4400), .I1(n4418), .I2(n4419), .O(n4457));
  LUT3 #(.INIT(8'hE8)) lut_n4458 (.I0(n4438), .I1(n4456), .I2(n4457), .O(n4458));
  LUT3 #(.INIT(8'h96)) lut_n4459 (.I0(n4342), .I1(n4380), .I2(n4381), .O(n4459));
  LUT3 #(.INIT(8'hE8)) lut_n4460 (.I0(n4420), .I1(n4458), .I2(n4459), .O(n4460));
  LUT3 #(.INIT(8'h96)) lut_n4461 (.I0(n4224), .I1(n4302), .I2(n4303), .O(n4461));
  LUT3 #(.INIT(8'hE8)) lut_n4462 (.I0(n4382), .I1(n4460), .I2(n4461), .O(n4462));
  LUT3 #(.INIT(8'h96)) lut_n4463 (.I0(n3982), .I1(n4140), .I2(n4141), .O(n4463));
  LUT3 #(.INIT(8'hE8)) lut_n4464 (.I0(n4304), .I1(n4462), .I2(n4463), .O(n4464));
  LUT3 #(.INIT(8'h96)) lut_n4465 (.I0(x942), .I1(x943), .I2(x944), .O(n4465));
  LUT5 #(.INIT(32'h96696996)) lut_n4466 (.I0(x933), .I1(x934), .I2(x935), .I3(n4450), .I4(n4451), .O(n4466));
  LUT5 #(.INIT(32'hFF969600)) lut_n4467 (.I0(x939), .I1(x940), .I2(x941), .I3(n4465), .I4(n4466), .O(n4467));
  LUT3 #(.INIT(8'h96)) lut_n4468 (.I0(x948), .I1(x949), .I2(x950), .O(n4468));
  LUT5 #(.INIT(32'h96696996)) lut_n4469 (.I0(x939), .I1(x940), .I2(x941), .I3(n4465), .I4(n4466), .O(n4469));
  LUT5 #(.INIT(32'hFF969600)) lut_n4470 (.I0(x945), .I1(x946), .I2(x947), .I3(n4468), .I4(n4469), .O(n4470));
  LUT3 #(.INIT(8'h96)) lut_n4471 (.I0(n4449), .I1(n4452), .I2(n4453), .O(n4471));
  LUT3 #(.INIT(8'hE8)) lut_n4472 (.I0(n4467), .I1(n4470), .I2(n4471), .O(n4472));
  LUT3 #(.INIT(8'h96)) lut_n4473 (.I0(x954), .I1(x955), .I2(x956), .O(n4473));
  LUT5 #(.INIT(32'h96696996)) lut_n4474 (.I0(x945), .I1(x946), .I2(x947), .I3(n4468), .I4(n4469), .O(n4474));
  LUT5 #(.INIT(32'hFF969600)) lut_n4475 (.I0(x951), .I1(x952), .I2(x953), .I3(n4473), .I4(n4474), .O(n4475));
  LUT3 #(.INIT(8'h96)) lut_n4476 (.I0(x960), .I1(x961), .I2(x962), .O(n4476));
  LUT5 #(.INIT(32'h96696996)) lut_n4477 (.I0(x951), .I1(x952), .I2(x953), .I3(n4473), .I4(n4474), .O(n4477));
  LUT5 #(.INIT(32'hFF969600)) lut_n4478 (.I0(x957), .I1(x958), .I2(x959), .I3(n4476), .I4(n4477), .O(n4478));
  LUT3 #(.INIT(8'h96)) lut_n4479 (.I0(n4467), .I1(n4470), .I2(n4471), .O(n4479));
  LUT3 #(.INIT(8'hE8)) lut_n4480 (.I0(n4475), .I1(n4478), .I2(n4479), .O(n4480));
  LUT3 #(.INIT(8'h96)) lut_n4481 (.I0(n4446), .I1(n4454), .I2(n4455), .O(n4481));
  LUT3 #(.INIT(8'hE8)) lut_n4482 (.I0(n4472), .I1(n4480), .I2(n4481), .O(n4482));
  LUT3 #(.INIT(8'h96)) lut_n4483 (.I0(x966), .I1(x967), .I2(x968), .O(n4483));
  LUT5 #(.INIT(32'h96696996)) lut_n4484 (.I0(x957), .I1(x958), .I2(x959), .I3(n4476), .I4(n4477), .O(n4484));
  LUT5 #(.INIT(32'hFF969600)) lut_n4485 (.I0(x963), .I1(x964), .I2(x965), .I3(n4483), .I4(n4484), .O(n4485));
  LUT3 #(.INIT(8'h96)) lut_n4486 (.I0(x972), .I1(x973), .I2(x974), .O(n4486));
  LUT5 #(.INIT(32'h96696996)) lut_n4487 (.I0(x963), .I1(x964), .I2(x965), .I3(n4483), .I4(n4484), .O(n4487));
  LUT5 #(.INIT(32'hFF969600)) lut_n4488 (.I0(x969), .I1(x970), .I2(x971), .I3(n4486), .I4(n4487), .O(n4488));
  LUT3 #(.INIT(8'h96)) lut_n4489 (.I0(n4475), .I1(n4478), .I2(n4479), .O(n4489));
  LUT3 #(.INIT(8'hE8)) lut_n4490 (.I0(n4485), .I1(n4488), .I2(n4489), .O(n4490));
  LUT3 #(.INIT(8'h96)) lut_n4491 (.I0(x978), .I1(x979), .I2(x980), .O(n4491));
  LUT5 #(.INIT(32'h96696996)) lut_n4492 (.I0(x969), .I1(x970), .I2(x971), .I3(n4486), .I4(n4487), .O(n4492));
  LUT5 #(.INIT(32'hFF969600)) lut_n4493 (.I0(x975), .I1(x976), .I2(x977), .I3(n4491), .I4(n4492), .O(n4493));
  LUT3 #(.INIT(8'h96)) lut_n4494 (.I0(x984), .I1(x985), .I2(x986), .O(n4494));
  LUT5 #(.INIT(32'h96696996)) lut_n4495 (.I0(x975), .I1(x976), .I2(x977), .I3(n4491), .I4(n4492), .O(n4495));
  LUT5 #(.INIT(32'hFF969600)) lut_n4496 (.I0(x981), .I1(x982), .I2(x983), .I3(n4494), .I4(n4495), .O(n4496));
  LUT3 #(.INIT(8'h96)) lut_n4497 (.I0(n4485), .I1(n4488), .I2(n4489), .O(n4497));
  LUT3 #(.INIT(8'hE8)) lut_n4498 (.I0(n4493), .I1(n4496), .I2(n4497), .O(n4498));
  LUT3 #(.INIT(8'h96)) lut_n4499 (.I0(n4472), .I1(n4480), .I2(n4481), .O(n4499));
  LUT3 #(.INIT(8'hE8)) lut_n4500 (.I0(n4490), .I1(n4498), .I2(n4499), .O(n4500));
  LUT3 #(.INIT(8'h96)) lut_n4501 (.I0(n4438), .I1(n4456), .I2(n4457), .O(n4501));
  LUT3 #(.INIT(8'hE8)) lut_n4502 (.I0(n4482), .I1(n4500), .I2(n4501), .O(n4502));
  LUT3 #(.INIT(8'h96)) lut_n4503 (.I0(x990), .I1(x991), .I2(x992), .O(n4503));
  LUT5 #(.INIT(32'h96696996)) lut_n4504 (.I0(x981), .I1(x982), .I2(x983), .I3(n4494), .I4(n4495), .O(n4504));
  LUT5 #(.INIT(32'hFF969600)) lut_n4505 (.I0(x987), .I1(x988), .I2(x989), .I3(n4503), .I4(n4504), .O(n4505));
  LUT3 #(.INIT(8'h96)) lut_n4506 (.I0(x996), .I1(x997), .I2(x998), .O(n4506));
  LUT5 #(.INIT(32'h96696996)) lut_n4507 (.I0(x987), .I1(x988), .I2(x989), .I3(n4503), .I4(n4504), .O(n4507));
  LUT5 #(.INIT(32'hFF969600)) lut_n4508 (.I0(x993), .I1(x994), .I2(x995), .I3(n4506), .I4(n4507), .O(n4508));
  LUT3 #(.INIT(8'h96)) lut_n4509 (.I0(n4493), .I1(n4496), .I2(n4497), .O(n4509));
  LUT3 #(.INIT(8'hE8)) lut_n4510 (.I0(n4505), .I1(n4508), .I2(n4509), .O(n4510));
  LUT3 #(.INIT(8'h96)) lut_n4511 (.I0(x1002), .I1(x1003), .I2(x1004), .O(n4511));
  LUT5 #(.INIT(32'h96696996)) lut_n4512 (.I0(x993), .I1(x994), .I2(x995), .I3(n4506), .I4(n4507), .O(n4512));
  LUT5 #(.INIT(32'hFF969600)) lut_n4513 (.I0(x999), .I1(x1000), .I2(x1001), .I3(n4511), .I4(n4512), .O(n4513));
  LUT3 #(.INIT(8'h96)) lut_n4514 (.I0(x1008), .I1(x1009), .I2(x1010), .O(n4514));
  LUT5 #(.INIT(32'h96696996)) lut_n4515 (.I0(x999), .I1(x1000), .I2(x1001), .I3(n4511), .I4(n4512), .O(n4515));
  LUT5 #(.INIT(32'hFF969600)) lut_n4516 (.I0(x1005), .I1(x1006), .I2(x1007), .I3(n4514), .I4(n4515), .O(n4516));
  LUT3 #(.INIT(8'h96)) lut_n4517 (.I0(n4505), .I1(n4508), .I2(n4509), .O(n4517));
  LUT3 #(.INIT(8'hE8)) lut_n4518 (.I0(n4513), .I1(n4516), .I2(n4517), .O(n4518));
  LUT3 #(.INIT(8'h96)) lut_n4519 (.I0(n4490), .I1(n4498), .I2(n4499), .O(n4519));
  LUT3 #(.INIT(8'hE8)) lut_n4520 (.I0(n4510), .I1(n4518), .I2(n4519), .O(n4520));
  LUT3 #(.INIT(8'h96)) lut_n4521 (.I0(x1014), .I1(x1015), .I2(x1016), .O(n4521));
  LUT5 #(.INIT(32'h96696996)) lut_n4522 (.I0(x1005), .I1(x1006), .I2(x1007), .I3(n4514), .I4(n4515), .O(n4522));
  LUT5 #(.INIT(32'hFF969600)) lut_n4523 (.I0(x1011), .I1(x1012), .I2(x1013), .I3(n4521), .I4(n4522), .O(n4523));
  LUT3 #(.INIT(8'h96)) lut_n4524 (.I0(x1020), .I1(x1021), .I2(x1022), .O(n4524));
  LUT5 #(.INIT(32'h96696996)) lut_n4525 (.I0(x1011), .I1(x1012), .I2(x1013), .I3(n4521), .I4(n4522), .O(n4525));
  LUT5 #(.INIT(32'hFF969600)) lut_n4526 (.I0(x1017), .I1(x1018), .I2(x1019), .I3(n4524), .I4(n4525), .O(n4526));
  LUT3 #(.INIT(8'h96)) lut_n4527 (.I0(n4513), .I1(n4516), .I2(n4517), .O(n4527));
  LUT3 #(.INIT(8'hE8)) lut_n4528 (.I0(n4523), .I1(n4526), .I2(n4527), .O(n4528));
  LUT3 #(.INIT(8'h96)) lut_n4529 (.I0(x1026), .I1(x1027), .I2(x1028), .O(n4529));
  LUT5 #(.INIT(32'h96696996)) lut_n4530 (.I0(x1017), .I1(x1018), .I2(x1019), .I3(n4524), .I4(n4525), .O(n4530));
  LUT5 #(.INIT(32'hFF969600)) lut_n4531 (.I0(x1023), .I1(x1024), .I2(x1025), .I3(n4529), .I4(n4530), .O(n4531));
  LUT3 #(.INIT(8'h96)) lut_n4532 (.I0(x1032), .I1(x1033), .I2(x1034), .O(n4532));
  LUT5 #(.INIT(32'h96696996)) lut_n4533 (.I0(x1023), .I1(x1024), .I2(x1025), .I3(n4529), .I4(n4530), .O(n4533));
  LUT5 #(.INIT(32'hFF969600)) lut_n4534 (.I0(x1029), .I1(x1030), .I2(x1031), .I3(n4532), .I4(n4533), .O(n4534));
  LUT3 #(.INIT(8'h96)) lut_n4535 (.I0(n4523), .I1(n4526), .I2(n4527), .O(n4535));
  LUT3 #(.INIT(8'hE8)) lut_n4536 (.I0(n4531), .I1(n4534), .I2(n4535), .O(n4536));
  LUT3 #(.INIT(8'h96)) lut_n4537 (.I0(n4510), .I1(n4518), .I2(n4519), .O(n4537));
  LUT3 #(.INIT(8'hE8)) lut_n4538 (.I0(n4528), .I1(n4536), .I2(n4537), .O(n4538));
  LUT3 #(.INIT(8'h96)) lut_n4539 (.I0(n4482), .I1(n4500), .I2(n4501), .O(n4539));
  LUT3 #(.INIT(8'hE8)) lut_n4540 (.I0(n4520), .I1(n4538), .I2(n4539), .O(n4540));
  LUT3 #(.INIT(8'h96)) lut_n4541 (.I0(n4420), .I1(n4458), .I2(n4459), .O(n4541));
  LUT3 #(.INIT(8'hE8)) lut_n4542 (.I0(n4502), .I1(n4540), .I2(n4541), .O(n4542));
  LUT3 #(.INIT(8'h96)) lut_n4543 (.I0(x1038), .I1(x1039), .I2(x1040), .O(n4543));
  LUT5 #(.INIT(32'h96696996)) lut_n4544 (.I0(x1029), .I1(x1030), .I2(x1031), .I3(n4532), .I4(n4533), .O(n4544));
  LUT5 #(.INIT(32'hFF969600)) lut_n4545 (.I0(x1035), .I1(x1036), .I2(x1037), .I3(n4543), .I4(n4544), .O(n4545));
  LUT3 #(.INIT(8'h96)) lut_n4546 (.I0(x1044), .I1(x1045), .I2(x1046), .O(n4546));
  LUT5 #(.INIT(32'h96696996)) lut_n4547 (.I0(x1035), .I1(x1036), .I2(x1037), .I3(n4543), .I4(n4544), .O(n4547));
  LUT5 #(.INIT(32'hFF969600)) lut_n4548 (.I0(x1041), .I1(x1042), .I2(x1043), .I3(n4546), .I4(n4547), .O(n4548));
  LUT3 #(.INIT(8'h96)) lut_n4549 (.I0(n4531), .I1(n4534), .I2(n4535), .O(n4549));
  LUT3 #(.INIT(8'hE8)) lut_n4550 (.I0(n4545), .I1(n4548), .I2(n4549), .O(n4550));
  LUT3 #(.INIT(8'h96)) lut_n4551 (.I0(x1050), .I1(x1051), .I2(x1052), .O(n4551));
  LUT5 #(.INIT(32'h96696996)) lut_n4552 (.I0(x1041), .I1(x1042), .I2(x1043), .I3(n4546), .I4(n4547), .O(n4552));
  LUT5 #(.INIT(32'hFF969600)) lut_n4553 (.I0(x1047), .I1(x1048), .I2(x1049), .I3(n4551), .I4(n4552), .O(n4553));
  LUT3 #(.INIT(8'h96)) lut_n4554 (.I0(x1056), .I1(x1057), .I2(x1058), .O(n4554));
  LUT5 #(.INIT(32'h96696996)) lut_n4555 (.I0(x1047), .I1(x1048), .I2(x1049), .I3(n4551), .I4(n4552), .O(n4555));
  LUT5 #(.INIT(32'hFF969600)) lut_n4556 (.I0(x1053), .I1(x1054), .I2(x1055), .I3(n4554), .I4(n4555), .O(n4556));
  LUT3 #(.INIT(8'h96)) lut_n4557 (.I0(n4545), .I1(n4548), .I2(n4549), .O(n4557));
  LUT3 #(.INIT(8'hE8)) lut_n4558 (.I0(n4553), .I1(n4556), .I2(n4557), .O(n4558));
  LUT3 #(.INIT(8'h96)) lut_n4559 (.I0(n4528), .I1(n4536), .I2(n4537), .O(n4559));
  LUT3 #(.INIT(8'hE8)) lut_n4560 (.I0(n4550), .I1(n4558), .I2(n4559), .O(n4560));
  LUT3 #(.INIT(8'h96)) lut_n4561 (.I0(x1062), .I1(x1063), .I2(x1064), .O(n4561));
  LUT5 #(.INIT(32'h96696996)) lut_n4562 (.I0(x1053), .I1(x1054), .I2(x1055), .I3(n4554), .I4(n4555), .O(n4562));
  LUT5 #(.INIT(32'hFF969600)) lut_n4563 (.I0(x1059), .I1(x1060), .I2(x1061), .I3(n4561), .I4(n4562), .O(n4563));
  LUT3 #(.INIT(8'h96)) lut_n4564 (.I0(x1068), .I1(x1069), .I2(x1070), .O(n4564));
  LUT5 #(.INIT(32'h96696996)) lut_n4565 (.I0(x1059), .I1(x1060), .I2(x1061), .I3(n4561), .I4(n4562), .O(n4565));
  LUT5 #(.INIT(32'hFF969600)) lut_n4566 (.I0(x1065), .I1(x1066), .I2(x1067), .I3(n4564), .I4(n4565), .O(n4566));
  LUT3 #(.INIT(8'h96)) lut_n4567 (.I0(n4553), .I1(n4556), .I2(n4557), .O(n4567));
  LUT3 #(.INIT(8'hE8)) lut_n4568 (.I0(n4563), .I1(n4566), .I2(n4567), .O(n4568));
  LUT3 #(.INIT(8'h96)) lut_n4569 (.I0(x1074), .I1(x1075), .I2(x1076), .O(n4569));
  LUT5 #(.INIT(32'h96696996)) lut_n4570 (.I0(x1065), .I1(x1066), .I2(x1067), .I3(n4564), .I4(n4565), .O(n4570));
  LUT5 #(.INIT(32'hFF969600)) lut_n4571 (.I0(x1071), .I1(x1072), .I2(x1073), .I3(n4569), .I4(n4570), .O(n4571));
  LUT3 #(.INIT(8'h96)) lut_n4572 (.I0(x1080), .I1(x1081), .I2(x1082), .O(n4572));
  LUT5 #(.INIT(32'h96696996)) lut_n4573 (.I0(x1071), .I1(x1072), .I2(x1073), .I3(n4569), .I4(n4570), .O(n4573));
  LUT5 #(.INIT(32'hFF969600)) lut_n4574 (.I0(x1077), .I1(x1078), .I2(x1079), .I3(n4572), .I4(n4573), .O(n4574));
  LUT3 #(.INIT(8'h96)) lut_n4575 (.I0(n4563), .I1(n4566), .I2(n4567), .O(n4575));
  LUT3 #(.INIT(8'hE8)) lut_n4576 (.I0(n4571), .I1(n4574), .I2(n4575), .O(n4576));
  LUT3 #(.INIT(8'h96)) lut_n4577 (.I0(n4550), .I1(n4558), .I2(n4559), .O(n4577));
  LUT3 #(.INIT(8'hE8)) lut_n4578 (.I0(n4568), .I1(n4576), .I2(n4577), .O(n4578));
  LUT3 #(.INIT(8'h96)) lut_n4579 (.I0(n4520), .I1(n4538), .I2(n4539), .O(n4579));
  LUT3 #(.INIT(8'hE8)) lut_n4580 (.I0(n4560), .I1(n4578), .I2(n4579), .O(n4580));
  LUT3 #(.INIT(8'h96)) lut_n4581 (.I0(x1086), .I1(x1087), .I2(x1088), .O(n4581));
  LUT5 #(.INIT(32'h96696996)) lut_n4582 (.I0(x1077), .I1(x1078), .I2(x1079), .I3(n4572), .I4(n4573), .O(n4582));
  LUT5 #(.INIT(32'hFF969600)) lut_n4583 (.I0(x1083), .I1(x1084), .I2(x1085), .I3(n4581), .I4(n4582), .O(n4583));
  LUT3 #(.INIT(8'h96)) lut_n4584 (.I0(x1092), .I1(x1093), .I2(x1094), .O(n4584));
  LUT5 #(.INIT(32'h96696996)) lut_n4585 (.I0(x1083), .I1(x1084), .I2(x1085), .I3(n4581), .I4(n4582), .O(n4585));
  LUT5 #(.INIT(32'hFF969600)) lut_n4586 (.I0(x1089), .I1(x1090), .I2(x1091), .I3(n4584), .I4(n4585), .O(n4586));
  LUT3 #(.INIT(8'h96)) lut_n4587 (.I0(n4571), .I1(n4574), .I2(n4575), .O(n4587));
  LUT3 #(.INIT(8'hE8)) lut_n4588 (.I0(n4583), .I1(n4586), .I2(n4587), .O(n4588));
  LUT3 #(.INIT(8'h96)) lut_n4589 (.I0(x1098), .I1(x1099), .I2(x1100), .O(n4589));
  LUT5 #(.INIT(32'h96696996)) lut_n4590 (.I0(x1089), .I1(x1090), .I2(x1091), .I3(n4584), .I4(n4585), .O(n4590));
  LUT5 #(.INIT(32'hFF969600)) lut_n4591 (.I0(x1095), .I1(x1096), .I2(x1097), .I3(n4589), .I4(n4590), .O(n4591));
  LUT3 #(.INIT(8'h96)) lut_n4592 (.I0(x1104), .I1(x1105), .I2(x1106), .O(n4592));
  LUT5 #(.INIT(32'h96696996)) lut_n4593 (.I0(x1095), .I1(x1096), .I2(x1097), .I3(n4589), .I4(n4590), .O(n4593));
  LUT5 #(.INIT(32'hFF969600)) lut_n4594 (.I0(x1101), .I1(x1102), .I2(x1103), .I3(n4592), .I4(n4593), .O(n4594));
  LUT3 #(.INIT(8'h96)) lut_n4595 (.I0(n4583), .I1(n4586), .I2(n4587), .O(n4595));
  LUT3 #(.INIT(8'hE8)) lut_n4596 (.I0(n4591), .I1(n4594), .I2(n4595), .O(n4596));
  LUT3 #(.INIT(8'h96)) lut_n4597 (.I0(n4568), .I1(n4576), .I2(n4577), .O(n4597));
  LUT3 #(.INIT(8'hE8)) lut_n4598 (.I0(n4588), .I1(n4596), .I2(n4597), .O(n4598));
  LUT3 #(.INIT(8'h96)) lut_n4599 (.I0(x1110), .I1(x1111), .I2(x1112), .O(n4599));
  LUT5 #(.INIT(32'h96696996)) lut_n4600 (.I0(x1101), .I1(x1102), .I2(x1103), .I3(n4592), .I4(n4593), .O(n4600));
  LUT5 #(.INIT(32'hFF969600)) lut_n4601 (.I0(x1107), .I1(x1108), .I2(x1109), .I3(n4599), .I4(n4600), .O(n4601));
  LUT3 #(.INIT(8'h96)) lut_n4602 (.I0(x1116), .I1(x1117), .I2(x1118), .O(n4602));
  LUT5 #(.INIT(32'h96696996)) lut_n4603 (.I0(x1107), .I1(x1108), .I2(x1109), .I3(n4599), .I4(n4600), .O(n4603));
  LUT5 #(.INIT(32'hFF969600)) lut_n4604 (.I0(x1113), .I1(x1114), .I2(x1115), .I3(n4602), .I4(n4603), .O(n4604));
  LUT3 #(.INIT(8'h96)) lut_n4605 (.I0(n4591), .I1(n4594), .I2(n4595), .O(n4605));
  LUT3 #(.INIT(8'hE8)) lut_n4606 (.I0(n4601), .I1(n4604), .I2(n4605), .O(n4606));
  LUT3 #(.INIT(8'h96)) lut_n4607 (.I0(x1122), .I1(x1123), .I2(x1124), .O(n4607));
  LUT5 #(.INIT(32'h96696996)) lut_n4608 (.I0(x1113), .I1(x1114), .I2(x1115), .I3(n4602), .I4(n4603), .O(n4608));
  LUT5 #(.INIT(32'hFF969600)) lut_n4609 (.I0(x1119), .I1(x1120), .I2(x1121), .I3(n4607), .I4(n4608), .O(n4609));
  LUT3 #(.INIT(8'h96)) lut_n4610 (.I0(x1128), .I1(x1129), .I2(x1130), .O(n4610));
  LUT5 #(.INIT(32'h96696996)) lut_n4611 (.I0(x1119), .I1(x1120), .I2(x1121), .I3(n4607), .I4(n4608), .O(n4611));
  LUT5 #(.INIT(32'hFF969600)) lut_n4612 (.I0(x1125), .I1(x1126), .I2(x1127), .I3(n4610), .I4(n4611), .O(n4612));
  LUT3 #(.INIT(8'h96)) lut_n4613 (.I0(n4601), .I1(n4604), .I2(n4605), .O(n4613));
  LUT3 #(.INIT(8'hE8)) lut_n4614 (.I0(n4609), .I1(n4612), .I2(n4613), .O(n4614));
  LUT3 #(.INIT(8'h96)) lut_n4615 (.I0(n4588), .I1(n4596), .I2(n4597), .O(n4615));
  LUT3 #(.INIT(8'hE8)) lut_n4616 (.I0(n4606), .I1(n4614), .I2(n4615), .O(n4616));
  LUT3 #(.INIT(8'h96)) lut_n4617 (.I0(n4560), .I1(n4578), .I2(n4579), .O(n4617));
  LUT3 #(.INIT(8'hE8)) lut_n4618 (.I0(n4598), .I1(n4616), .I2(n4617), .O(n4618));
  LUT3 #(.INIT(8'h96)) lut_n4619 (.I0(n4502), .I1(n4540), .I2(n4541), .O(n4619));
  LUT3 #(.INIT(8'hE8)) lut_n4620 (.I0(n4580), .I1(n4618), .I2(n4619), .O(n4620));
  LUT3 #(.INIT(8'h96)) lut_n4621 (.I0(n4382), .I1(n4460), .I2(n4461), .O(n4621));
  LUT3 #(.INIT(8'hE8)) lut_n4622 (.I0(n4542), .I1(n4620), .I2(n4621), .O(n4622));
  LUT3 #(.INIT(8'h96)) lut_n4623 (.I0(x1134), .I1(x1135), .I2(x1136), .O(n4623));
  LUT5 #(.INIT(32'h96696996)) lut_n4624 (.I0(x1125), .I1(x1126), .I2(x1127), .I3(n4610), .I4(n4611), .O(n4624));
  LUT5 #(.INIT(32'hFF969600)) lut_n4625 (.I0(x1131), .I1(x1132), .I2(x1133), .I3(n4623), .I4(n4624), .O(n4625));
  LUT3 #(.INIT(8'h96)) lut_n4626 (.I0(x1140), .I1(x1141), .I2(x1142), .O(n4626));
  LUT5 #(.INIT(32'h96696996)) lut_n4627 (.I0(x1131), .I1(x1132), .I2(x1133), .I3(n4623), .I4(n4624), .O(n4627));
  LUT5 #(.INIT(32'hFF969600)) lut_n4628 (.I0(x1137), .I1(x1138), .I2(x1139), .I3(n4626), .I4(n4627), .O(n4628));
  LUT3 #(.INIT(8'h96)) lut_n4629 (.I0(n4609), .I1(n4612), .I2(n4613), .O(n4629));
  LUT3 #(.INIT(8'hE8)) lut_n4630 (.I0(n4625), .I1(n4628), .I2(n4629), .O(n4630));
  LUT3 #(.INIT(8'h96)) lut_n4631 (.I0(x1146), .I1(x1147), .I2(x1148), .O(n4631));
  LUT5 #(.INIT(32'h96696996)) lut_n4632 (.I0(x1137), .I1(x1138), .I2(x1139), .I3(n4626), .I4(n4627), .O(n4632));
  LUT5 #(.INIT(32'hFF969600)) lut_n4633 (.I0(x1143), .I1(x1144), .I2(x1145), .I3(n4631), .I4(n4632), .O(n4633));
  LUT3 #(.INIT(8'h96)) lut_n4634 (.I0(x1152), .I1(x1153), .I2(x1154), .O(n4634));
  LUT5 #(.INIT(32'h96696996)) lut_n4635 (.I0(x1143), .I1(x1144), .I2(x1145), .I3(n4631), .I4(n4632), .O(n4635));
  LUT5 #(.INIT(32'hFF969600)) lut_n4636 (.I0(x1149), .I1(x1150), .I2(x1151), .I3(n4634), .I4(n4635), .O(n4636));
  LUT3 #(.INIT(8'h96)) lut_n4637 (.I0(n4625), .I1(n4628), .I2(n4629), .O(n4637));
  LUT3 #(.INIT(8'hE8)) lut_n4638 (.I0(n4633), .I1(n4636), .I2(n4637), .O(n4638));
  LUT3 #(.INIT(8'h96)) lut_n4639 (.I0(n4606), .I1(n4614), .I2(n4615), .O(n4639));
  LUT3 #(.INIT(8'hE8)) lut_n4640 (.I0(n4630), .I1(n4638), .I2(n4639), .O(n4640));
  LUT3 #(.INIT(8'h96)) lut_n4641 (.I0(x1158), .I1(x1159), .I2(x1160), .O(n4641));
  LUT5 #(.INIT(32'h96696996)) lut_n4642 (.I0(x1149), .I1(x1150), .I2(x1151), .I3(n4634), .I4(n4635), .O(n4642));
  LUT5 #(.INIT(32'hFF969600)) lut_n4643 (.I0(x1155), .I1(x1156), .I2(x1157), .I3(n4641), .I4(n4642), .O(n4643));
  LUT3 #(.INIT(8'h96)) lut_n4644 (.I0(x1164), .I1(x1165), .I2(x1166), .O(n4644));
  LUT5 #(.INIT(32'h96696996)) lut_n4645 (.I0(x1155), .I1(x1156), .I2(x1157), .I3(n4641), .I4(n4642), .O(n4645));
  LUT5 #(.INIT(32'hFF969600)) lut_n4646 (.I0(x1161), .I1(x1162), .I2(x1163), .I3(n4644), .I4(n4645), .O(n4646));
  LUT3 #(.INIT(8'h96)) lut_n4647 (.I0(n4633), .I1(n4636), .I2(n4637), .O(n4647));
  LUT3 #(.INIT(8'hE8)) lut_n4648 (.I0(n4643), .I1(n4646), .I2(n4647), .O(n4648));
  LUT3 #(.INIT(8'h96)) lut_n4649 (.I0(x1170), .I1(x1171), .I2(x1172), .O(n4649));
  LUT5 #(.INIT(32'h96696996)) lut_n4650 (.I0(x1161), .I1(x1162), .I2(x1163), .I3(n4644), .I4(n4645), .O(n4650));
  LUT5 #(.INIT(32'hFF969600)) lut_n4651 (.I0(x1167), .I1(x1168), .I2(x1169), .I3(n4649), .I4(n4650), .O(n4651));
  LUT3 #(.INIT(8'h96)) lut_n4652 (.I0(x1176), .I1(x1177), .I2(x1178), .O(n4652));
  LUT5 #(.INIT(32'h96696996)) lut_n4653 (.I0(x1167), .I1(x1168), .I2(x1169), .I3(n4649), .I4(n4650), .O(n4653));
  LUT5 #(.INIT(32'hFF969600)) lut_n4654 (.I0(x1173), .I1(x1174), .I2(x1175), .I3(n4652), .I4(n4653), .O(n4654));
  LUT3 #(.INIT(8'h96)) lut_n4655 (.I0(n4643), .I1(n4646), .I2(n4647), .O(n4655));
  LUT3 #(.INIT(8'hE8)) lut_n4656 (.I0(n4651), .I1(n4654), .I2(n4655), .O(n4656));
  LUT3 #(.INIT(8'h96)) lut_n4657 (.I0(n4630), .I1(n4638), .I2(n4639), .O(n4657));
  LUT3 #(.INIT(8'hE8)) lut_n4658 (.I0(n4648), .I1(n4656), .I2(n4657), .O(n4658));
  LUT3 #(.INIT(8'h96)) lut_n4659 (.I0(n4598), .I1(n4616), .I2(n4617), .O(n4659));
  LUT3 #(.INIT(8'hE8)) lut_n4660 (.I0(n4640), .I1(n4658), .I2(n4659), .O(n4660));
  LUT3 #(.INIT(8'h96)) lut_n4661 (.I0(x1182), .I1(x1183), .I2(x1184), .O(n4661));
  LUT5 #(.INIT(32'h96696996)) lut_n4662 (.I0(x1173), .I1(x1174), .I2(x1175), .I3(n4652), .I4(n4653), .O(n4662));
  LUT5 #(.INIT(32'hFF969600)) lut_n4663 (.I0(x1179), .I1(x1180), .I2(x1181), .I3(n4661), .I4(n4662), .O(n4663));
  LUT3 #(.INIT(8'h96)) lut_n4664 (.I0(x1188), .I1(x1189), .I2(x1190), .O(n4664));
  LUT5 #(.INIT(32'h96696996)) lut_n4665 (.I0(x1179), .I1(x1180), .I2(x1181), .I3(n4661), .I4(n4662), .O(n4665));
  LUT5 #(.INIT(32'hFF969600)) lut_n4666 (.I0(x1185), .I1(x1186), .I2(x1187), .I3(n4664), .I4(n4665), .O(n4666));
  LUT3 #(.INIT(8'h96)) lut_n4667 (.I0(n4651), .I1(n4654), .I2(n4655), .O(n4667));
  LUT3 #(.INIT(8'hE8)) lut_n4668 (.I0(n4663), .I1(n4666), .I2(n4667), .O(n4668));
  LUT3 #(.INIT(8'h96)) lut_n4669 (.I0(x1194), .I1(x1195), .I2(x1196), .O(n4669));
  LUT5 #(.INIT(32'h96696996)) lut_n4670 (.I0(x1185), .I1(x1186), .I2(x1187), .I3(n4664), .I4(n4665), .O(n4670));
  LUT5 #(.INIT(32'hFF969600)) lut_n4671 (.I0(x1191), .I1(x1192), .I2(x1193), .I3(n4669), .I4(n4670), .O(n4671));
  LUT3 #(.INIT(8'h96)) lut_n4672 (.I0(x1200), .I1(x1201), .I2(x1202), .O(n4672));
  LUT5 #(.INIT(32'h96696996)) lut_n4673 (.I0(x1191), .I1(x1192), .I2(x1193), .I3(n4669), .I4(n4670), .O(n4673));
  LUT5 #(.INIT(32'hFF969600)) lut_n4674 (.I0(x1197), .I1(x1198), .I2(x1199), .I3(n4672), .I4(n4673), .O(n4674));
  LUT3 #(.INIT(8'h96)) lut_n4675 (.I0(n4663), .I1(n4666), .I2(n4667), .O(n4675));
  LUT3 #(.INIT(8'hE8)) lut_n4676 (.I0(n4671), .I1(n4674), .I2(n4675), .O(n4676));
  LUT3 #(.INIT(8'h96)) lut_n4677 (.I0(n4648), .I1(n4656), .I2(n4657), .O(n4677));
  LUT3 #(.INIT(8'hE8)) lut_n4678 (.I0(n4668), .I1(n4676), .I2(n4677), .O(n4678));
  LUT3 #(.INIT(8'h96)) lut_n4679 (.I0(x1206), .I1(x1207), .I2(x1208), .O(n4679));
  LUT5 #(.INIT(32'h96696996)) lut_n4680 (.I0(x1197), .I1(x1198), .I2(x1199), .I3(n4672), .I4(n4673), .O(n4680));
  LUT5 #(.INIT(32'hFF969600)) lut_n4681 (.I0(x1203), .I1(x1204), .I2(x1205), .I3(n4679), .I4(n4680), .O(n4681));
  LUT3 #(.INIT(8'h96)) lut_n4682 (.I0(x1212), .I1(x1213), .I2(x1214), .O(n4682));
  LUT5 #(.INIT(32'h96696996)) lut_n4683 (.I0(x1203), .I1(x1204), .I2(x1205), .I3(n4679), .I4(n4680), .O(n4683));
  LUT5 #(.INIT(32'hFF969600)) lut_n4684 (.I0(x1209), .I1(x1210), .I2(x1211), .I3(n4682), .I4(n4683), .O(n4684));
  LUT3 #(.INIT(8'h96)) lut_n4685 (.I0(n4671), .I1(n4674), .I2(n4675), .O(n4685));
  LUT3 #(.INIT(8'hE8)) lut_n4686 (.I0(n4681), .I1(n4684), .I2(n4685), .O(n4686));
  LUT3 #(.INIT(8'h96)) lut_n4687 (.I0(x1218), .I1(x1219), .I2(x1220), .O(n4687));
  LUT5 #(.INIT(32'h96696996)) lut_n4688 (.I0(x1209), .I1(x1210), .I2(x1211), .I3(n4682), .I4(n4683), .O(n4688));
  LUT5 #(.INIT(32'hFF969600)) lut_n4689 (.I0(x1215), .I1(x1216), .I2(x1217), .I3(n4687), .I4(n4688), .O(n4689));
  LUT3 #(.INIT(8'h96)) lut_n4690 (.I0(x1224), .I1(x1225), .I2(x1226), .O(n4690));
  LUT5 #(.INIT(32'h96696996)) lut_n4691 (.I0(x1215), .I1(x1216), .I2(x1217), .I3(n4687), .I4(n4688), .O(n4691));
  LUT5 #(.INIT(32'hFF969600)) lut_n4692 (.I0(x1221), .I1(x1222), .I2(x1223), .I3(n4690), .I4(n4691), .O(n4692));
  LUT3 #(.INIT(8'h96)) lut_n4693 (.I0(n4681), .I1(n4684), .I2(n4685), .O(n4693));
  LUT3 #(.INIT(8'hE8)) lut_n4694 (.I0(n4689), .I1(n4692), .I2(n4693), .O(n4694));
  LUT3 #(.INIT(8'h96)) lut_n4695 (.I0(n4668), .I1(n4676), .I2(n4677), .O(n4695));
  LUT3 #(.INIT(8'hE8)) lut_n4696 (.I0(n4686), .I1(n4694), .I2(n4695), .O(n4696));
  LUT3 #(.INIT(8'h96)) lut_n4697 (.I0(n4640), .I1(n4658), .I2(n4659), .O(n4697));
  LUT3 #(.INIT(8'hE8)) lut_n4698 (.I0(n4678), .I1(n4696), .I2(n4697), .O(n4698));
  LUT3 #(.INIT(8'h96)) lut_n4699 (.I0(n4580), .I1(n4618), .I2(n4619), .O(n4699));
  LUT3 #(.INIT(8'hE8)) lut_n4700 (.I0(n4660), .I1(n4698), .I2(n4699), .O(n4700));
  LUT3 #(.INIT(8'h96)) lut_n4701 (.I0(x1230), .I1(x1231), .I2(x1232), .O(n4701));
  LUT5 #(.INIT(32'h96696996)) lut_n4702 (.I0(x1221), .I1(x1222), .I2(x1223), .I3(n4690), .I4(n4691), .O(n4702));
  LUT5 #(.INIT(32'hFF969600)) lut_n4703 (.I0(x1227), .I1(x1228), .I2(x1229), .I3(n4701), .I4(n4702), .O(n4703));
  LUT3 #(.INIT(8'h96)) lut_n4704 (.I0(x1236), .I1(x1237), .I2(x1238), .O(n4704));
  LUT5 #(.INIT(32'h96696996)) lut_n4705 (.I0(x1227), .I1(x1228), .I2(x1229), .I3(n4701), .I4(n4702), .O(n4705));
  LUT5 #(.INIT(32'hFF969600)) lut_n4706 (.I0(x1233), .I1(x1234), .I2(x1235), .I3(n4704), .I4(n4705), .O(n4706));
  LUT3 #(.INIT(8'h96)) lut_n4707 (.I0(n4689), .I1(n4692), .I2(n4693), .O(n4707));
  LUT3 #(.INIT(8'hE8)) lut_n4708 (.I0(n4703), .I1(n4706), .I2(n4707), .O(n4708));
  LUT3 #(.INIT(8'h96)) lut_n4709 (.I0(x1242), .I1(x1243), .I2(x1244), .O(n4709));
  LUT5 #(.INIT(32'h96696996)) lut_n4710 (.I0(x1233), .I1(x1234), .I2(x1235), .I3(n4704), .I4(n4705), .O(n4710));
  LUT5 #(.INIT(32'hFF969600)) lut_n4711 (.I0(x1239), .I1(x1240), .I2(x1241), .I3(n4709), .I4(n4710), .O(n4711));
  LUT3 #(.INIT(8'h96)) lut_n4712 (.I0(x1248), .I1(x1249), .I2(x1250), .O(n4712));
  LUT5 #(.INIT(32'h96696996)) lut_n4713 (.I0(x1239), .I1(x1240), .I2(x1241), .I3(n4709), .I4(n4710), .O(n4713));
  LUT5 #(.INIT(32'hFF969600)) lut_n4714 (.I0(x1245), .I1(x1246), .I2(x1247), .I3(n4712), .I4(n4713), .O(n4714));
  LUT3 #(.INIT(8'h96)) lut_n4715 (.I0(n4703), .I1(n4706), .I2(n4707), .O(n4715));
  LUT3 #(.INIT(8'hE8)) lut_n4716 (.I0(n4711), .I1(n4714), .I2(n4715), .O(n4716));
  LUT3 #(.INIT(8'h96)) lut_n4717 (.I0(n4686), .I1(n4694), .I2(n4695), .O(n4717));
  LUT3 #(.INIT(8'hE8)) lut_n4718 (.I0(n4708), .I1(n4716), .I2(n4717), .O(n4718));
  LUT3 #(.INIT(8'h96)) lut_n4719 (.I0(x1254), .I1(x1255), .I2(x1256), .O(n4719));
  LUT5 #(.INIT(32'h96696996)) lut_n4720 (.I0(x1245), .I1(x1246), .I2(x1247), .I3(n4712), .I4(n4713), .O(n4720));
  LUT5 #(.INIT(32'hFF969600)) lut_n4721 (.I0(x1251), .I1(x1252), .I2(x1253), .I3(n4719), .I4(n4720), .O(n4721));
  LUT3 #(.INIT(8'h96)) lut_n4722 (.I0(x1260), .I1(x1261), .I2(x1262), .O(n4722));
  LUT5 #(.INIT(32'h96696996)) lut_n4723 (.I0(x1251), .I1(x1252), .I2(x1253), .I3(n4719), .I4(n4720), .O(n4723));
  LUT5 #(.INIT(32'hFF969600)) lut_n4724 (.I0(x1257), .I1(x1258), .I2(x1259), .I3(n4722), .I4(n4723), .O(n4724));
  LUT3 #(.INIT(8'h96)) lut_n4725 (.I0(n4711), .I1(n4714), .I2(n4715), .O(n4725));
  LUT3 #(.INIT(8'hE8)) lut_n4726 (.I0(n4721), .I1(n4724), .I2(n4725), .O(n4726));
  LUT3 #(.INIT(8'h96)) lut_n4727 (.I0(x1266), .I1(x1267), .I2(x1268), .O(n4727));
  LUT5 #(.INIT(32'h96696996)) lut_n4728 (.I0(x1257), .I1(x1258), .I2(x1259), .I3(n4722), .I4(n4723), .O(n4728));
  LUT5 #(.INIT(32'hFF969600)) lut_n4729 (.I0(x1263), .I1(x1264), .I2(x1265), .I3(n4727), .I4(n4728), .O(n4729));
  LUT3 #(.INIT(8'h96)) lut_n4730 (.I0(x1272), .I1(x1273), .I2(x1274), .O(n4730));
  LUT5 #(.INIT(32'h96696996)) lut_n4731 (.I0(x1263), .I1(x1264), .I2(x1265), .I3(n4727), .I4(n4728), .O(n4731));
  LUT5 #(.INIT(32'hFF969600)) lut_n4732 (.I0(x1269), .I1(x1270), .I2(x1271), .I3(n4730), .I4(n4731), .O(n4732));
  LUT3 #(.INIT(8'h96)) lut_n4733 (.I0(n4721), .I1(n4724), .I2(n4725), .O(n4733));
  LUT3 #(.INIT(8'hE8)) lut_n4734 (.I0(n4729), .I1(n4732), .I2(n4733), .O(n4734));
  LUT3 #(.INIT(8'h96)) lut_n4735 (.I0(n4708), .I1(n4716), .I2(n4717), .O(n4735));
  LUT3 #(.INIT(8'hE8)) lut_n4736 (.I0(n4726), .I1(n4734), .I2(n4735), .O(n4736));
  LUT3 #(.INIT(8'h96)) lut_n4737 (.I0(n4678), .I1(n4696), .I2(n4697), .O(n4737));
  LUT3 #(.INIT(8'hE8)) lut_n4738 (.I0(n4718), .I1(n4736), .I2(n4737), .O(n4738));
  LUT3 #(.INIT(8'h96)) lut_n4739 (.I0(x1278), .I1(x1279), .I2(x1280), .O(n4739));
  LUT5 #(.INIT(32'h96696996)) lut_n4740 (.I0(x1269), .I1(x1270), .I2(x1271), .I3(n4730), .I4(n4731), .O(n4740));
  LUT5 #(.INIT(32'hFF969600)) lut_n4741 (.I0(x1275), .I1(x1276), .I2(x1277), .I3(n4739), .I4(n4740), .O(n4741));
  LUT3 #(.INIT(8'h96)) lut_n4742 (.I0(x1284), .I1(x1285), .I2(x1286), .O(n4742));
  LUT5 #(.INIT(32'h96696996)) lut_n4743 (.I0(x1275), .I1(x1276), .I2(x1277), .I3(n4739), .I4(n4740), .O(n4743));
  LUT5 #(.INIT(32'hFF969600)) lut_n4744 (.I0(x1281), .I1(x1282), .I2(x1283), .I3(n4742), .I4(n4743), .O(n4744));
  LUT3 #(.INIT(8'h96)) lut_n4745 (.I0(n4729), .I1(n4732), .I2(n4733), .O(n4745));
  LUT3 #(.INIT(8'hE8)) lut_n4746 (.I0(n4741), .I1(n4744), .I2(n4745), .O(n4746));
  LUT3 #(.INIT(8'h96)) lut_n4747 (.I0(x1290), .I1(x1291), .I2(x1292), .O(n4747));
  LUT5 #(.INIT(32'h96696996)) lut_n4748 (.I0(x1281), .I1(x1282), .I2(x1283), .I3(n4742), .I4(n4743), .O(n4748));
  LUT5 #(.INIT(32'hFF969600)) lut_n4749 (.I0(x1287), .I1(x1288), .I2(x1289), .I3(n4747), .I4(n4748), .O(n4749));
  LUT3 #(.INIT(8'h96)) lut_n4750 (.I0(x1296), .I1(x1297), .I2(x1298), .O(n4750));
  LUT5 #(.INIT(32'h96696996)) lut_n4751 (.I0(x1287), .I1(x1288), .I2(x1289), .I3(n4747), .I4(n4748), .O(n4751));
  LUT5 #(.INIT(32'hFF969600)) lut_n4752 (.I0(x1293), .I1(x1294), .I2(x1295), .I3(n4750), .I4(n4751), .O(n4752));
  LUT3 #(.INIT(8'h96)) lut_n4753 (.I0(n4741), .I1(n4744), .I2(n4745), .O(n4753));
  LUT3 #(.INIT(8'hE8)) lut_n4754 (.I0(n4749), .I1(n4752), .I2(n4753), .O(n4754));
  LUT3 #(.INIT(8'h96)) lut_n4755 (.I0(n4726), .I1(n4734), .I2(n4735), .O(n4755));
  LUT3 #(.INIT(8'hE8)) lut_n4756 (.I0(n4746), .I1(n4754), .I2(n4755), .O(n4756));
  LUT3 #(.INIT(8'h96)) lut_n4757 (.I0(x1302), .I1(x1303), .I2(x1304), .O(n4757));
  LUT5 #(.INIT(32'h96696996)) lut_n4758 (.I0(x1293), .I1(x1294), .I2(x1295), .I3(n4750), .I4(n4751), .O(n4758));
  LUT5 #(.INIT(32'hFF969600)) lut_n4759 (.I0(x1299), .I1(x1300), .I2(x1301), .I3(n4757), .I4(n4758), .O(n4759));
  LUT3 #(.INIT(8'h96)) lut_n4760 (.I0(x1308), .I1(x1309), .I2(x1310), .O(n4760));
  LUT5 #(.INIT(32'h96696996)) lut_n4761 (.I0(x1299), .I1(x1300), .I2(x1301), .I3(n4757), .I4(n4758), .O(n4761));
  LUT5 #(.INIT(32'hFF969600)) lut_n4762 (.I0(x1305), .I1(x1306), .I2(x1307), .I3(n4760), .I4(n4761), .O(n4762));
  LUT3 #(.INIT(8'h96)) lut_n4763 (.I0(n4749), .I1(n4752), .I2(n4753), .O(n4763));
  LUT3 #(.INIT(8'hE8)) lut_n4764 (.I0(n4759), .I1(n4762), .I2(n4763), .O(n4764));
  LUT3 #(.INIT(8'h96)) lut_n4765 (.I0(x1314), .I1(x1315), .I2(x1316), .O(n4765));
  LUT5 #(.INIT(32'h96696996)) lut_n4766 (.I0(x1305), .I1(x1306), .I2(x1307), .I3(n4760), .I4(n4761), .O(n4766));
  LUT5 #(.INIT(32'hFF969600)) lut_n4767 (.I0(x1311), .I1(x1312), .I2(x1313), .I3(n4765), .I4(n4766), .O(n4767));
  LUT3 #(.INIT(8'h96)) lut_n4768 (.I0(x1320), .I1(x1321), .I2(x1322), .O(n4768));
  LUT5 #(.INIT(32'h96696996)) lut_n4769 (.I0(x1311), .I1(x1312), .I2(x1313), .I3(n4765), .I4(n4766), .O(n4769));
  LUT5 #(.INIT(32'hFF969600)) lut_n4770 (.I0(x1317), .I1(x1318), .I2(x1319), .I3(n4768), .I4(n4769), .O(n4770));
  LUT3 #(.INIT(8'h96)) lut_n4771 (.I0(n4759), .I1(n4762), .I2(n4763), .O(n4771));
  LUT3 #(.INIT(8'hE8)) lut_n4772 (.I0(n4767), .I1(n4770), .I2(n4771), .O(n4772));
  LUT3 #(.INIT(8'h96)) lut_n4773 (.I0(n4746), .I1(n4754), .I2(n4755), .O(n4773));
  LUT3 #(.INIT(8'hE8)) lut_n4774 (.I0(n4764), .I1(n4772), .I2(n4773), .O(n4774));
  LUT3 #(.INIT(8'h96)) lut_n4775 (.I0(n4718), .I1(n4736), .I2(n4737), .O(n4775));
  LUT3 #(.INIT(8'hE8)) lut_n4776 (.I0(n4756), .I1(n4774), .I2(n4775), .O(n4776));
  LUT3 #(.INIT(8'h96)) lut_n4777 (.I0(n4660), .I1(n4698), .I2(n4699), .O(n4777));
  LUT3 #(.INIT(8'hE8)) lut_n4778 (.I0(n4738), .I1(n4776), .I2(n4777), .O(n4778));
  LUT3 #(.INIT(8'h96)) lut_n4779 (.I0(n4542), .I1(n4620), .I2(n4621), .O(n4779));
  LUT3 #(.INIT(8'hE8)) lut_n4780 (.I0(n4700), .I1(n4778), .I2(n4779), .O(n4780));
  LUT3 #(.INIT(8'h96)) lut_n4781 (.I0(n4304), .I1(n4462), .I2(n4463), .O(n4781));
  LUT3 #(.INIT(8'hE8)) lut_n4782 (.I0(n4622), .I1(n4780), .I2(n4781), .O(n4782));
  LUT3 #(.INIT(8'h96)) lut_n4783 (.I0(n3824), .I1(n4142), .I2(n4143), .O(n4783));
  LUT3 #(.INIT(8'hE8)) lut_n4784 (.I0(n4464), .I1(n4782), .I2(n4783), .O(n4784));
  LUT3 #(.INIT(8'h96)) lut_n4785 (.I0(x1326), .I1(x1327), .I2(x1328), .O(n4785));
  LUT5 #(.INIT(32'h96696996)) lut_n4786 (.I0(x1317), .I1(x1318), .I2(x1319), .I3(n4768), .I4(n4769), .O(n4786));
  LUT5 #(.INIT(32'hFF969600)) lut_n4787 (.I0(x1323), .I1(x1324), .I2(x1325), .I3(n4785), .I4(n4786), .O(n4787));
  LUT3 #(.INIT(8'h96)) lut_n4788 (.I0(x1332), .I1(x1333), .I2(x1334), .O(n4788));
  LUT5 #(.INIT(32'h96696996)) lut_n4789 (.I0(x1323), .I1(x1324), .I2(x1325), .I3(n4785), .I4(n4786), .O(n4789));
  LUT5 #(.INIT(32'hFF969600)) lut_n4790 (.I0(x1329), .I1(x1330), .I2(x1331), .I3(n4788), .I4(n4789), .O(n4790));
  LUT3 #(.INIT(8'h96)) lut_n4791 (.I0(n4767), .I1(n4770), .I2(n4771), .O(n4791));
  LUT3 #(.INIT(8'hE8)) lut_n4792 (.I0(n4787), .I1(n4790), .I2(n4791), .O(n4792));
  LUT3 #(.INIT(8'h96)) lut_n4793 (.I0(x1338), .I1(x1339), .I2(x1340), .O(n4793));
  LUT5 #(.INIT(32'h96696996)) lut_n4794 (.I0(x1329), .I1(x1330), .I2(x1331), .I3(n4788), .I4(n4789), .O(n4794));
  LUT5 #(.INIT(32'hFF969600)) lut_n4795 (.I0(x1335), .I1(x1336), .I2(x1337), .I3(n4793), .I4(n4794), .O(n4795));
  LUT3 #(.INIT(8'h96)) lut_n4796 (.I0(x1344), .I1(x1345), .I2(x1346), .O(n4796));
  LUT5 #(.INIT(32'h96696996)) lut_n4797 (.I0(x1335), .I1(x1336), .I2(x1337), .I3(n4793), .I4(n4794), .O(n4797));
  LUT5 #(.INIT(32'hFF969600)) lut_n4798 (.I0(x1341), .I1(x1342), .I2(x1343), .I3(n4796), .I4(n4797), .O(n4798));
  LUT3 #(.INIT(8'h96)) lut_n4799 (.I0(n4787), .I1(n4790), .I2(n4791), .O(n4799));
  LUT3 #(.INIT(8'hE8)) lut_n4800 (.I0(n4795), .I1(n4798), .I2(n4799), .O(n4800));
  LUT3 #(.INIT(8'h96)) lut_n4801 (.I0(n4764), .I1(n4772), .I2(n4773), .O(n4801));
  LUT3 #(.INIT(8'hE8)) lut_n4802 (.I0(n4792), .I1(n4800), .I2(n4801), .O(n4802));
  LUT3 #(.INIT(8'h96)) lut_n4803 (.I0(x1350), .I1(x1351), .I2(x1352), .O(n4803));
  LUT5 #(.INIT(32'h96696996)) lut_n4804 (.I0(x1341), .I1(x1342), .I2(x1343), .I3(n4796), .I4(n4797), .O(n4804));
  LUT5 #(.INIT(32'hFF969600)) lut_n4805 (.I0(x1347), .I1(x1348), .I2(x1349), .I3(n4803), .I4(n4804), .O(n4805));
  LUT3 #(.INIT(8'h96)) lut_n4806 (.I0(x1356), .I1(x1357), .I2(x1358), .O(n4806));
  LUT5 #(.INIT(32'h96696996)) lut_n4807 (.I0(x1347), .I1(x1348), .I2(x1349), .I3(n4803), .I4(n4804), .O(n4807));
  LUT5 #(.INIT(32'hFF969600)) lut_n4808 (.I0(x1353), .I1(x1354), .I2(x1355), .I3(n4806), .I4(n4807), .O(n4808));
  LUT3 #(.INIT(8'h96)) lut_n4809 (.I0(n4795), .I1(n4798), .I2(n4799), .O(n4809));
  LUT3 #(.INIT(8'hE8)) lut_n4810 (.I0(n4805), .I1(n4808), .I2(n4809), .O(n4810));
  LUT3 #(.INIT(8'h96)) lut_n4811 (.I0(x1362), .I1(x1363), .I2(x1364), .O(n4811));
  LUT5 #(.INIT(32'h96696996)) lut_n4812 (.I0(x1353), .I1(x1354), .I2(x1355), .I3(n4806), .I4(n4807), .O(n4812));
  LUT5 #(.INIT(32'hFF969600)) lut_n4813 (.I0(x1359), .I1(x1360), .I2(x1361), .I3(n4811), .I4(n4812), .O(n4813));
  LUT3 #(.INIT(8'h96)) lut_n4814 (.I0(x1368), .I1(x1369), .I2(x1370), .O(n4814));
  LUT5 #(.INIT(32'h96696996)) lut_n4815 (.I0(x1359), .I1(x1360), .I2(x1361), .I3(n4811), .I4(n4812), .O(n4815));
  LUT5 #(.INIT(32'hFF969600)) lut_n4816 (.I0(x1365), .I1(x1366), .I2(x1367), .I3(n4814), .I4(n4815), .O(n4816));
  LUT3 #(.INIT(8'h96)) lut_n4817 (.I0(n4805), .I1(n4808), .I2(n4809), .O(n4817));
  LUT3 #(.INIT(8'hE8)) lut_n4818 (.I0(n4813), .I1(n4816), .I2(n4817), .O(n4818));
  LUT3 #(.INIT(8'h96)) lut_n4819 (.I0(n4792), .I1(n4800), .I2(n4801), .O(n4819));
  LUT3 #(.INIT(8'hE8)) lut_n4820 (.I0(n4810), .I1(n4818), .I2(n4819), .O(n4820));
  LUT3 #(.INIT(8'h96)) lut_n4821 (.I0(n4756), .I1(n4774), .I2(n4775), .O(n4821));
  LUT3 #(.INIT(8'hE8)) lut_n4822 (.I0(n4802), .I1(n4820), .I2(n4821), .O(n4822));
  LUT3 #(.INIT(8'h96)) lut_n4823 (.I0(x1374), .I1(x1375), .I2(x1376), .O(n4823));
  LUT5 #(.INIT(32'h96696996)) lut_n4824 (.I0(x1365), .I1(x1366), .I2(x1367), .I3(n4814), .I4(n4815), .O(n4824));
  LUT5 #(.INIT(32'hFF969600)) lut_n4825 (.I0(x1371), .I1(x1372), .I2(x1373), .I3(n4823), .I4(n4824), .O(n4825));
  LUT3 #(.INIT(8'h96)) lut_n4826 (.I0(x1380), .I1(x1381), .I2(x1382), .O(n4826));
  LUT5 #(.INIT(32'h96696996)) lut_n4827 (.I0(x1371), .I1(x1372), .I2(x1373), .I3(n4823), .I4(n4824), .O(n4827));
  LUT5 #(.INIT(32'hFF969600)) lut_n4828 (.I0(x1377), .I1(x1378), .I2(x1379), .I3(n4826), .I4(n4827), .O(n4828));
  LUT3 #(.INIT(8'h96)) lut_n4829 (.I0(n4813), .I1(n4816), .I2(n4817), .O(n4829));
  LUT3 #(.INIT(8'hE8)) lut_n4830 (.I0(n4825), .I1(n4828), .I2(n4829), .O(n4830));
  LUT3 #(.INIT(8'h96)) lut_n4831 (.I0(x1386), .I1(x1387), .I2(x1388), .O(n4831));
  LUT5 #(.INIT(32'h96696996)) lut_n4832 (.I0(x1377), .I1(x1378), .I2(x1379), .I3(n4826), .I4(n4827), .O(n4832));
  LUT5 #(.INIT(32'hFF969600)) lut_n4833 (.I0(x1383), .I1(x1384), .I2(x1385), .I3(n4831), .I4(n4832), .O(n4833));
  LUT3 #(.INIT(8'h96)) lut_n4834 (.I0(x1392), .I1(x1393), .I2(x1394), .O(n4834));
  LUT5 #(.INIT(32'h96696996)) lut_n4835 (.I0(x1383), .I1(x1384), .I2(x1385), .I3(n4831), .I4(n4832), .O(n4835));
  LUT5 #(.INIT(32'hFF969600)) lut_n4836 (.I0(x1389), .I1(x1390), .I2(x1391), .I3(n4834), .I4(n4835), .O(n4836));
  LUT3 #(.INIT(8'h96)) lut_n4837 (.I0(n4825), .I1(n4828), .I2(n4829), .O(n4837));
  LUT3 #(.INIT(8'hE8)) lut_n4838 (.I0(n4833), .I1(n4836), .I2(n4837), .O(n4838));
  LUT3 #(.INIT(8'h96)) lut_n4839 (.I0(n4810), .I1(n4818), .I2(n4819), .O(n4839));
  LUT3 #(.INIT(8'hE8)) lut_n4840 (.I0(n4830), .I1(n4838), .I2(n4839), .O(n4840));
  LUT3 #(.INIT(8'h96)) lut_n4841 (.I0(x1398), .I1(x1399), .I2(x1400), .O(n4841));
  LUT5 #(.INIT(32'h96696996)) lut_n4842 (.I0(x1389), .I1(x1390), .I2(x1391), .I3(n4834), .I4(n4835), .O(n4842));
  LUT5 #(.INIT(32'hFF969600)) lut_n4843 (.I0(x1395), .I1(x1396), .I2(x1397), .I3(n4841), .I4(n4842), .O(n4843));
  LUT3 #(.INIT(8'h96)) lut_n4844 (.I0(x1404), .I1(x1405), .I2(x1406), .O(n4844));
  LUT5 #(.INIT(32'h96696996)) lut_n4845 (.I0(x1395), .I1(x1396), .I2(x1397), .I3(n4841), .I4(n4842), .O(n4845));
  LUT5 #(.INIT(32'hFF969600)) lut_n4846 (.I0(x1401), .I1(x1402), .I2(x1403), .I3(n4844), .I4(n4845), .O(n4846));
  LUT3 #(.INIT(8'h96)) lut_n4847 (.I0(n4833), .I1(n4836), .I2(n4837), .O(n4847));
  LUT3 #(.INIT(8'hE8)) lut_n4848 (.I0(n4843), .I1(n4846), .I2(n4847), .O(n4848));
  LUT3 #(.INIT(8'h96)) lut_n4849 (.I0(x1410), .I1(x1411), .I2(x1412), .O(n4849));
  LUT5 #(.INIT(32'h96696996)) lut_n4850 (.I0(x1401), .I1(x1402), .I2(x1403), .I3(n4844), .I4(n4845), .O(n4850));
  LUT5 #(.INIT(32'hFF969600)) lut_n4851 (.I0(x1407), .I1(x1408), .I2(x1409), .I3(n4849), .I4(n4850), .O(n4851));
  LUT3 #(.INIT(8'h96)) lut_n4852 (.I0(x1416), .I1(x1417), .I2(x1418), .O(n4852));
  LUT5 #(.INIT(32'h96696996)) lut_n4853 (.I0(x1407), .I1(x1408), .I2(x1409), .I3(n4849), .I4(n4850), .O(n4853));
  LUT5 #(.INIT(32'hFF969600)) lut_n4854 (.I0(x1413), .I1(x1414), .I2(x1415), .I3(n4852), .I4(n4853), .O(n4854));
  LUT3 #(.INIT(8'h96)) lut_n4855 (.I0(n4843), .I1(n4846), .I2(n4847), .O(n4855));
  LUT3 #(.INIT(8'hE8)) lut_n4856 (.I0(n4851), .I1(n4854), .I2(n4855), .O(n4856));
  LUT3 #(.INIT(8'h96)) lut_n4857 (.I0(n4830), .I1(n4838), .I2(n4839), .O(n4857));
  LUT3 #(.INIT(8'hE8)) lut_n4858 (.I0(n4848), .I1(n4856), .I2(n4857), .O(n4858));
  LUT3 #(.INIT(8'h96)) lut_n4859 (.I0(n4802), .I1(n4820), .I2(n4821), .O(n4859));
  LUT3 #(.INIT(8'hE8)) lut_n4860 (.I0(n4840), .I1(n4858), .I2(n4859), .O(n4860));
  LUT3 #(.INIT(8'h96)) lut_n4861 (.I0(n4738), .I1(n4776), .I2(n4777), .O(n4861));
  LUT3 #(.INIT(8'hE8)) lut_n4862 (.I0(n4822), .I1(n4860), .I2(n4861), .O(n4862));
  LUT3 #(.INIT(8'h96)) lut_n4863 (.I0(x1422), .I1(x1423), .I2(x1424), .O(n4863));
  LUT5 #(.INIT(32'h96696996)) lut_n4864 (.I0(x1413), .I1(x1414), .I2(x1415), .I3(n4852), .I4(n4853), .O(n4864));
  LUT5 #(.INIT(32'hFF969600)) lut_n4865 (.I0(x1419), .I1(x1420), .I2(x1421), .I3(n4863), .I4(n4864), .O(n4865));
  LUT3 #(.INIT(8'h96)) lut_n4866 (.I0(x1428), .I1(x1429), .I2(x1430), .O(n4866));
  LUT5 #(.INIT(32'h96696996)) lut_n4867 (.I0(x1419), .I1(x1420), .I2(x1421), .I3(n4863), .I4(n4864), .O(n4867));
  LUT5 #(.INIT(32'hFF969600)) lut_n4868 (.I0(x1425), .I1(x1426), .I2(x1427), .I3(n4866), .I4(n4867), .O(n4868));
  LUT3 #(.INIT(8'h96)) lut_n4869 (.I0(n4851), .I1(n4854), .I2(n4855), .O(n4869));
  LUT3 #(.INIT(8'hE8)) lut_n4870 (.I0(n4865), .I1(n4868), .I2(n4869), .O(n4870));
  LUT3 #(.INIT(8'h96)) lut_n4871 (.I0(x1434), .I1(x1435), .I2(x1436), .O(n4871));
  LUT5 #(.INIT(32'h96696996)) lut_n4872 (.I0(x1425), .I1(x1426), .I2(x1427), .I3(n4866), .I4(n4867), .O(n4872));
  LUT5 #(.INIT(32'hFF969600)) lut_n4873 (.I0(x1431), .I1(x1432), .I2(x1433), .I3(n4871), .I4(n4872), .O(n4873));
  LUT3 #(.INIT(8'h96)) lut_n4874 (.I0(x1440), .I1(x1441), .I2(x1442), .O(n4874));
  LUT5 #(.INIT(32'h96696996)) lut_n4875 (.I0(x1431), .I1(x1432), .I2(x1433), .I3(n4871), .I4(n4872), .O(n4875));
  LUT5 #(.INIT(32'hFF969600)) lut_n4876 (.I0(x1437), .I1(x1438), .I2(x1439), .I3(n4874), .I4(n4875), .O(n4876));
  LUT3 #(.INIT(8'h96)) lut_n4877 (.I0(n4865), .I1(n4868), .I2(n4869), .O(n4877));
  LUT3 #(.INIT(8'hE8)) lut_n4878 (.I0(n4873), .I1(n4876), .I2(n4877), .O(n4878));
  LUT3 #(.INIT(8'h96)) lut_n4879 (.I0(n4848), .I1(n4856), .I2(n4857), .O(n4879));
  LUT3 #(.INIT(8'hE8)) lut_n4880 (.I0(n4870), .I1(n4878), .I2(n4879), .O(n4880));
  LUT3 #(.INIT(8'h96)) lut_n4881 (.I0(x1446), .I1(x1447), .I2(x1448), .O(n4881));
  LUT5 #(.INIT(32'h96696996)) lut_n4882 (.I0(x1437), .I1(x1438), .I2(x1439), .I3(n4874), .I4(n4875), .O(n4882));
  LUT5 #(.INIT(32'hFF969600)) lut_n4883 (.I0(x1443), .I1(x1444), .I2(x1445), .I3(n4881), .I4(n4882), .O(n4883));
  LUT3 #(.INIT(8'h96)) lut_n4884 (.I0(x1452), .I1(x1453), .I2(x1454), .O(n4884));
  LUT5 #(.INIT(32'h96696996)) lut_n4885 (.I0(x1443), .I1(x1444), .I2(x1445), .I3(n4881), .I4(n4882), .O(n4885));
  LUT5 #(.INIT(32'hFF969600)) lut_n4886 (.I0(x1449), .I1(x1450), .I2(x1451), .I3(n4884), .I4(n4885), .O(n4886));
  LUT3 #(.INIT(8'h96)) lut_n4887 (.I0(n4873), .I1(n4876), .I2(n4877), .O(n4887));
  LUT3 #(.INIT(8'hE8)) lut_n4888 (.I0(n4883), .I1(n4886), .I2(n4887), .O(n4888));
  LUT3 #(.INIT(8'h96)) lut_n4889 (.I0(x1458), .I1(x1459), .I2(x1460), .O(n4889));
  LUT5 #(.INIT(32'h96696996)) lut_n4890 (.I0(x1449), .I1(x1450), .I2(x1451), .I3(n4884), .I4(n4885), .O(n4890));
  LUT5 #(.INIT(32'hFF969600)) lut_n4891 (.I0(x1455), .I1(x1456), .I2(x1457), .I3(n4889), .I4(n4890), .O(n4891));
  LUT3 #(.INIT(8'h96)) lut_n4892 (.I0(x1464), .I1(x1465), .I2(x1466), .O(n4892));
  LUT5 #(.INIT(32'h96696996)) lut_n4893 (.I0(x1455), .I1(x1456), .I2(x1457), .I3(n4889), .I4(n4890), .O(n4893));
  LUT5 #(.INIT(32'hFF969600)) lut_n4894 (.I0(x1461), .I1(x1462), .I2(x1463), .I3(n4892), .I4(n4893), .O(n4894));
  LUT3 #(.INIT(8'h96)) lut_n4895 (.I0(n4883), .I1(n4886), .I2(n4887), .O(n4895));
  LUT3 #(.INIT(8'hE8)) lut_n4896 (.I0(n4891), .I1(n4894), .I2(n4895), .O(n4896));
  LUT3 #(.INIT(8'h96)) lut_n4897 (.I0(n4870), .I1(n4878), .I2(n4879), .O(n4897));
  LUT3 #(.INIT(8'hE8)) lut_n4898 (.I0(n4888), .I1(n4896), .I2(n4897), .O(n4898));
  LUT3 #(.INIT(8'h96)) lut_n4899 (.I0(n4840), .I1(n4858), .I2(n4859), .O(n4899));
  LUT3 #(.INIT(8'hE8)) lut_n4900 (.I0(n4880), .I1(n4898), .I2(n4899), .O(n4900));
  LUT3 #(.INIT(8'h96)) lut_n4901 (.I0(x1470), .I1(x1471), .I2(x1472), .O(n4901));
  LUT5 #(.INIT(32'h96696996)) lut_n4902 (.I0(x1461), .I1(x1462), .I2(x1463), .I3(n4892), .I4(n4893), .O(n4902));
  LUT5 #(.INIT(32'hFF969600)) lut_n4903 (.I0(x1467), .I1(x1468), .I2(x1469), .I3(n4901), .I4(n4902), .O(n4903));
  LUT3 #(.INIT(8'h96)) lut_n4904 (.I0(x1476), .I1(x1477), .I2(x1478), .O(n4904));
  LUT5 #(.INIT(32'h96696996)) lut_n4905 (.I0(x1467), .I1(x1468), .I2(x1469), .I3(n4901), .I4(n4902), .O(n4905));
  LUT5 #(.INIT(32'hFF969600)) lut_n4906 (.I0(x1473), .I1(x1474), .I2(x1475), .I3(n4904), .I4(n4905), .O(n4906));
  LUT3 #(.INIT(8'h96)) lut_n4907 (.I0(n4891), .I1(n4894), .I2(n4895), .O(n4907));
  LUT3 #(.INIT(8'hE8)) lut_n4908 (.I0(n4903), .I1(n4906), .I2(n4907), .O(n4908));
  LUT3 #(.INIT(8'h96)) lut_n4909 (.I0(x1482), .I1(x1483), .I2(x1484), .O(n4909));
  LUT5 #(.INIT(32'h96696996)) lut_n4910 (.I0(x1473), .I1(x1474), .I2(x1475), .I3(n4904), .I4(n4905), .O(n4910));
  LUT5 #(.INIT(32'hFF969600)) lut_n4911 (.I0(x1479), .I1(x1480), .I2(x1481), .I3(n4909), .I4(n4910), .O(n4911));
  LUT3 #(.INIT(8'h96)) lut_n4912 (.I0(x1488), .I1(x1489), .I2(x1490), .O(n4912));
  LUT5 #(.INIT(32'h96696996)) lut_n4913 (.I0(x1479), .I1(x1480), .I2(x1481), .I3(n4909), .I4(n4910), .O(n4913));
  LUT5 #(.INIT(32'hFF969600)) lut_n4914 (.I0(x1485), .I1(x1486), .I2(x1487), .I3(n4912), .I4(n4913), .O(n4914));
  LUT3 #(.INIT(8'h96)) lut_n4915 (.I0(n4903), .I1(n4906), .I2(n4907), .O(n4915));
  LUT3 #(.INIT(8'hE8)) lut_n4916 (.I0(n4911), .I1(n4914), .I2(n4915), .O(n4916));
  LUT3 #(.INIT(8'h96)) lut_n4917 (.I0(n4888), .I1(n4896), .I2(n4897), .O(n4917));
  LUT3 #(.INIT(8'hE8)) lut_n4918 (.I0(n4908), .I1(n4916), .I2(n4917), .O(n4918));
  LUT3 #(.INIT(8'h96)) lut_n4919 (.I0(x1494), .I1(x1495), .I2(x1496), .O(n4919));
  LUT5 #(.INIT(32'h96696996)) lut_n4920 (.I0(x1485), .I1(x1486), .I2(x1487), .I3(n4912), .I4(n4913), .O(n4920));
  LUT5 #(.INIT(32'hFF969600)) lut_n4921 (.I0(x1491), .I1(x1492), .I2(x1493), .I3(n4919), .I4(n4920), .O(n4921));
  LUT3 #(.INIT(8'h96)) lut_n4922 (.I0(x1500), .I1(x1501), .I2(x1502), .O(n4922));
  LUT5 #(.INIT(32'h96696996)) lut_n4923 (.I0(x1491), .I1(x1492), .I2(x1493), .I3(n4919), .I4(n4920), .O(n4923));
  LUT5 #(.INIT(32'hFF969600)) lut_n4924 (.I0(x1497), .I1(x1498), .I2(x1499), .I3(n4922), .I4(n4923), .O(n4924));
  LUT3 #(.INIT(8'h96)) lut_n4925 (.I0(n4911), .I1(n4914), .I2(n4915), .O(n4925));
  LUT3 #(.INIT(8'hE8)) lut_n4926 (.I0(n4921), .I1(n4924), .I2(n4925), .O(n4926));
  LUT3 #(.INIT(8'h96)) lut_n4927 (.I0(x1506), .I1(x1507), .I2(x1508), .O(n4927));
  LUT5 #(.INIT(32'h96696996)) lut_n4928 (.I0(x1497), .I1(x1498), .I2(x1499), .I3(n4922), .I4(n4923), .O(n4928));
  LUT5 #(.INIT(32'hFF969600)) lut_n4929 (.I0(x1503), .I1(x1504), .I2(x1505), .I3(n4927), .I4(n4928), .O(n4929));
  LUT3 #(.INIT(8'h96)) lut_n4930 (.I0(x1512), .I1(x1513), .I2(x1514), .O(n4930));
  LUT5 #(.INIT(32'h96696996)) lut_n4931 (.I0(x1503), .I1(x1504), .I2(x1505), .I3(n4927), .I4(n4928), .O(n4931));
  LUT5 #(.INIT(32'hFF969600)) lut_n4932 (.I0(x1509), .I1(x1510), .I2(x1511), .I3(n4930), .I4(n4931), .O(n4932));
  LUT3 #(.INIT(8'h96)) lut_n4933 (.I0(n4921), .I1(n4924), .I2(n4925), .O(n4933));
  LUT3 #(.INIT(8'hE8)) lut_n4934 (.I0(n4929), .I1(n4932), .I2(n4933), .O(n4934));
  LUT3 #(.INIT(8'h96)) lut_n4935 (.I0(n4908), .I1(n4916), .I2(n4917), .O(n4935));
  LUT3 #(.INIT(8'hE8)) lut_n4936 (.I0(n4926), .I1(n4934), .I2(n4935), .O(n4936));
  LUT3 #(.INIT(8'h96)) lut_n4937 (.I0(n4880), .I1(n4898), .I2(n4899), .O(n4937));
  LUT3 #(.INIT(8'hE8)) lut_n4938 (.I0(n4918), .I1(n4936), .I2(n4937), .O(n4938));
  LUT3 #(.INIT(8'h96)) lut_n4939 (.I0(n4822), .I1(n4860), .I2(n4861), .O(n4939));
  LUT3 #(.INIT(8'hE8)) lut_n4940 (.I0(n4900), .I1(n4938), .I2(n4939), .O(n4940));
  LUT3 #(.INIT(8'h96)) lut_n4941 (.I0(n4700), .I1(n4778), .I2(n4779), .O(n4941));
  LUT3 #(.INIT(8'hE8)) lut_n4942 (.I0(n4862), .I1(n4940), .I2(n4941), .O(n4942));
  LUT3 #(.INIT(8'h96)) lut_n4943 (.I0(x1518), .I1(x1519), .I2(x1520), .O(n4943));
  LUT5 #(.INIT(32'h96696996)) lut_n4944 (.I0(x1509), .I1(x1510), .I2(x1511), .I3(n4930), .I4(n4931), .O(n4944));
  LUT5 #(.INIT(32'hFF969600)) lut_n4945 (.I0(x1515), .I1(x1516), .I2(x1517), .I3(n4943), .I4(n4944), .O(n4945));
  LUT3 #(.INIT(8'h96)) lut_n4946 (.I0(x1524), .I1(x1525), .I2(x1526), .O(n4946));
  LUT5 #(.INIT(32'h96696996)) lut_n4947 (.I0(x1515), .I1(x1516), .I2(x1517), .I3(n4943), .I4(n4944), .O(n4947));
  LUT5 #(.INIT(32'hFF969600)) lut_n4948 (.I0(x1521), .I1(x1522), .I2(x1523), .I3(n4946), .I4(n4947), .O(n4948));
  LUT3 #(.INIT(8'h96)) lut_n4949 (.I0(n4929), .I1(n4932), .I2(n4933), .O(n4949));
  LUT3 #(.INIT(8'hE8)) lut_n4950 (.I0(n4945), .I1(n4948), .I2(n4949), .O(n4950));
  LUT3 #(.INIT(8'h96)) lut_n4951 (.I0(x1530), .I1(x1531), .I2(x1532), .O(n4951));
  LUT5 #(.INIT(32'h96696996)) lut_n4952 (.I0(x1521), .I1(x1522), .I2(x1523), .I3(n4946), .I4(n4947), .O(n4952));
  LUT5 #(.INIT(32'hFF969600)) lut_n4953 (.I0(x1527), .I1(x1528), .I2(x1529), .I3(n4951), .I4(n4952), .O(n4953));
  LUT3 #(.INIT(8'h96)) lut_n4954 (.I0(x1536), .I1(x1537), .I2(x1538), .O(n4954));
  LUT5 #(.INIT(32'h96696996)) lut_n4955 (.I0(x1527), .I1(x1528), .I2(x1529), .I3(n4951), .I4(n4952), .O(n4955));
  LUT5 #(.INIT(32'hFF969600)) lut_n4956 (.I0(x1533), .I1(x1534), .I2(x1535), .I3(n4954), .I4(n4955), .O(n4956));
  LUT3 #(.INIT(8'h96)) lut_n4957 (.I0(n4945), .I1(n4948), .I2(n4949), .O(n4957));
  LUT3 #(.INIT(8'hE8)) lut_n4958 (.I0(n4953), .I1(n4956), .I2(n4957), .O(n4958));
  LUT3 #(.INIT(8'h96)) lut_n4959 (.I0(n4926), .I1(n4934), .I2(n4935), .O(n4959));
  LUT3 #(.INIT(8'hE8)) lut_n4960 (.I0(n4950), .I1(n4958), .I2(n4959), .O(n4960));
  LUT3 #(.INIT(8'h96)) lut_n4961 (.I0(x1542), .I1(x1543), .I2(x1544), .O(n4961));
  LUT5 #(.INIT(32'h96696996)) lut_n4962 (.I0(x1533), .I1(x1534), .I2(x1535), .I3(n4954), .I4(n4955), .O(n4962));
  LUT5 #(.INIT(32'hFF969600)) lut_n4963 (.I0(x1539), .I1(x1540), .I2(x1541), .I3(n4961), .I4(n4962), .O(n4963));
  LUT3 #(.INIT(8'h96)) lut_n4964 (.I0(x1548), .I1(x1549), .I2(x1550), .O(n4964));
  LUT5 #(.INIT(32'h96696996)) lut_n4965 (.I0(x1539), .I1(x1540), .I2(x1541), .I3(n4961), .I4(n4962), .O(n4965));
  LUT5 #(.INIT(32'hFF969600)) lut_n4966 (.I0(x1545), .I1(x1546), .I2(x1547), .I3(n4964), .I4(n4965), .O(n4966));
  LUT3 #(.INIT(8'h96)) lut_n4967 (.I0(n4953), .I1(n4956), .I2(n4957), .O(n4967));
  LUT3 #(.INIT(8'hE8)) lut_n4968 (.I0(n4963), .I1(n4966), .I2(n4967), .O(n4968));
  LUT3 #(.INIT(8'h96)) lut_n4969 (.I0(x1554), .I1(x1555), .I2(x1556), .O(n4969));
  LUT5 #(.INIT(32'h96696996)) lut_n4970 (.I0(x1545), .I1(x1546), .I2(x1547), .I3(n4964), .I4(n4965), .O(n4970));
  LUT5 #(.INIT(32'hFF969600)) lut_n4971 (.I0(x1551), .I1(x1552), .I2(x1553), .I3(n4969), .I4(n4970), .O(n4971));
  LUT3 #(.INIT(8'h96)) lut_n4972 (.I0(x1560), .I1(x1561), .I2(x1562), .O(n4972));
  LUT5 #(.INIT(32'h96696996)) lut_n4973 (.I0(x1551), .I1(x1552), .I2(x1553), .I3(n4969), .I4(n4970), .O(n4973));
  LUT5 #(.INIT(32'hFF969600)) lut_n4974 (.I0(x1557), .I1(x1558), .I2(x1559), .I3(n4972), .I4(n4973), .O(n4974));
  LUT3 #(.INIT(8'h96)) lut_n4975 (.I0(n4963), .I1(n4966), .I2(n4967), .O(n4975));
  LUT3 #(.INIT(8'hE8)) lut_n4976 (.I0(n4971), .I1(n4974), .I2(n4975), .O(n4976));
  LUT3 #(.INIT(8'h96)) lut_n4977 (.I0(n4950), .I1(n4958), .I2(n4959), .O(n4977));
  LUT3 #(.INIT(8'hE8)) lut_n4978 (.I0(n4968), .I1(n4976), .I2(n4977), .O(n4978));
  LUT3 #(.INIT(8'h96)) lut_n4979 (.I0(n4918), .I1(n4936), .I2(n4937), .O(n4979));
  LUT3 #(.INIT(8'hE8)) lut_n4980 (.I0(n4960), .I1(n4978), .I2(n4979), .O(n4980));
  LUT3 #(.INIT(8'h96)) lut_n4981 (.I0(x1566), .I1(x1567), .I2(x1568), .O(n4981));
  LUT5 #(.INIT(32'h96696996)) lut_n4982 (.I0(x1557), .I1(x1558), .I2(x1559), .I3(n4972), .I4(n4973), .O(n4982));
  LUT5 #(.INIT(32'hFF969600)) lut_n4983 (.I0(x1563), .I1(x1564), .I2(x1565), .I3(n4981), .I4(n4982), .O(n4983));
  LUT3 #(.INIT(8'h96)) lut_n4984 (.I0(x1572), .I1(x1573), .I2(x1574), .O(n4984));
  LUT5 #(.INIT(32'h96696996)) lut_n4985 (.I0(x1563), .I1(x1564), .I2(x1565), .I3(n4981), .I4(n4982), .O(n4985));
  LUT5 #(.INIT(32'hFF969600)) lut_n4986 (.I0(x1569), .I1(x1570), .I2(x1571), .I3(n4984), .I4(n4985), .O(n4986));
  LUT3 #(.INIT(8'h96)) lut_n4987 (.I0(n4971), .I1(n4974), .I2(n4975), .O(n4987));
  LUT3 #(.INIT(8'hE8)) lut_n4988 (.I0(n4983), .I1(n4986), .I2(n4987), .O(n4988));
  LUT3 #(.INIT(8'h96)) lut_n4989 (.I0(x1578), .I1(x1579), .I2(x1580), .O(n4989));
  LUT5 #(.INIT(32'h96696996)) lut_n4990 (.I0(x1569), .I1(x1570), .I2(x1571), .I3(n4984), .I4(n4985), .O(n4990));
  LUT5 #(.INIT(32'hFF969600)) lut_n4991 (.I0(x1575), .I1(x1576), .I2(x1577), .I3(n4989), .I4(n4990), .O(n4991));
  LUT3 #(.INIT(8'h96)) lut_n4992 (.I0(x1584), .I1(x1585), .I2(x1586), .O(n4992));
  LUT5 #(.INIT(32'h96696996)) lut_n4993 (.I0(x1575), .I1(x1576), .I2(x1577), .I3(n4989), .I4(n4990), .O(n4993));
  LUT5 #(.INIT(32'hFF969600)) lut_n4994 (.I0(x1581), .I1(x1582), .I2(x1583), .I3(n4992), .I4(n4993), .O(n4994));
  LUT3 #(.INIT(8'h96)) lut_n4995 (.I0(n4983), .I1(n4986), .I2(n4987), .O(n4995));
  LUT3 #(.INIT(8'hE8)) lut_n4996 (.I0(n4991), .I1(n4994), .I2(n4995), .O(n4996));
  LUT3 #(.INIT(8'h96)) lut_n4997 (.I0(n4968), .I1(n4976), .I2(n4977), .O(n4997));
  LUT3 #(.INIT(8'hE8)) lut_n4998 (.I0(n4988), .I1(n4996), .I2(n4997), .O(n4998));
  LUT3 #(.INIT(8'h96)) lut_n4999 (.I0(x1590), .I1(x1591), .I2(x1592), .O(n4999));
  LUT5 #(.INIT(32'h96696996)) lut_n5000 (.I0(x1581), .I1(x1582), .I2(x1583), .I3(n4992), .I4(n4993), .O(n5000));
  LUT5 #(.INIT(32'hFF969600)) lut_n5001 (.I0(x1587), .I1(x1588), .I2(x1589), .I3(n4999), .I4(n5000), .O(n5001));
  LUT3 #(.INIT(8'h96)) lut_n5002 (.I0(x1596), .I1(x1597), .I2(x1598), .O(n5002));
  LUT5 #(.INIT(32'h96696996)) lut_n5003 (.I0(x1587), .I1(x1588), .I2(x1589), .I3(n4999), .I4(n5000), .O(n5003));
  LUT5 #(.INIT(32'hFF969600)) lut_n5004 (.I0(x1593), .I1(x1594), .I2(x1595), .I3(n5002), .I4(n5003), .O(n5004));
  LUT3 #(.INIT(8'h96)) lut_n5005 (.I0(n4991), .I1(n4994), .I2(n4995), .O(n5005));
  LUT3 #(.INIT(8'hE8)) lut_n5006 (.I0(n5001), .I1(n5004), .I2(n5005), .O(n5006));
  LUT3 #(.INIT(8'h96)) lut_n5007 (.I0(x1602), .I1(x1603), .I2(x1604), .O(n5007));
  LUT5 #(.INIT(32'h96696996)) lut_n5008 (.I0(x1593), .I1(x1594), .I2(x1595), .I3(n5002), .I4(n5003), .O(n5008));
  LUT5 #(.INIT(32'hFF969600)) lut_n5009 (.I0(x1599), .I1(x1600), .I2(x1601), .I3(n5007), .I4(n5008), .O(n5009));
  LUT3 #(.INIT(8'h96)) lut_n5010 (.I0(x1608), .I1(x1609), .I2(x1610), .O(n5010));
  LUT5 #(.INIT(32'h96696996)) lut_n5011 (.I0(x1599), .I1(x1600), .I2(x1601), .I3(n5007), .I4(n5008), .O(n5011));
  LUT5 #(.INIT(32'hFF969600)) lut_n5012 (.I0(x1605), .I1(x1606), .I2(x1607), .I3(n5010), .I4(n5011), .O(n5012));
  LUT3 #(.INIT(8'h96)) lut_n5013 (.I0(n5001), .I1(n5004), .I2(n5005), .O(n5013));
  LUT3 #(.INIT(8'hE8)) lut_n5014 (.I0(n5009), .I1(n5012), .I2(n5013), .O(n5014));
  LUT3 #(.INIT(8'h96)) lut_n5015 (.I0(n4988), .I1(n4996), .I2(n4997), .O(n5015));
  LUT3 #(.INIT(8'hE8)) lut_n5016 (.I0(n5006), .I1(n5014), .I2(n5015), .O(n5016));
  LUT3 #(.INIT(8'h96)) lut_n5017 (.I0(n4960), .I1(n4978), .I2(n4979), .O(n5017));
  LUT3 #(.INIT(8'hE8)) lut_n5018 (.I0(n4998), .I1(n5016), .I2(n5017), .O(n5018));
  LUT3 #(.INIT(8'h96)) lut_n5019 (.I0(n4900), .I1(n4938), .I2(n4939), .O(n5019));
  LUT3 #(.INIT(8'hE8)) lut_n5020 (.I0(n4980), .I1(n5018), .I2(n5019), .O(n5020));
  LUT3 #(.INIT(8'h96)) lut_n5021 (.I0(x1614), .I1(x1615), .I2(x1616), .O(n5021));
  LUT5 #(.INIT(32'h96696996)) lut_n5022 (.I0(x1605), .I1(x1606), .I2(x1607), .I3(n5010), .I4(n5011), .O(n5022));
  LUT5 #(.INIT(32'hFF969600)) lut_n5023 (.I0(x1611), .I1(x1612), .I2(x1613), .I3(n5021), .I4(n5022), .O(n5023));
  LUT3 #(.INIT(8'h96)) lut_n5024 (.I0(x1620), .I1(x1621), .I2(x1622), .O(n5024));
  LUT5 #(.INIT(32'h96696996)) lut_n5025 (.I0(x1611), .I1(x1612), .I2(x1613), .I3(n5021), .I4(n5022), .O(n5025));
  LUT5 #(.INIT(32'hFF969600)) lut_n5026 (.I0(x1617), .I1(x1618), .I2(x1619), .I3(n5024), .I4(n5025), .O(n5026));
  LUT3 #(.INIT(8'h96)) lut_n5027 (.I0(n5009), .I1(n5012), .I2(n5013), .O(n5027));
  LUT3 #(.INIT(8'hE8)) lut_n5028 (.I0(n5023), .I1(n5026), .I2(n5027), .O(n5028));
  LUT3 #(.INIT(8'h96)) lut_n5029 (.I0(x1626), .I1(x1627), .I2(x1628), .O(n5029));
  LUT5 #(.INIT(32'h96696996)) lut_n5030 (.I0(x1617), .I1(x1618), .I2(x1619), .I3(n5024), .I4(n5025), .O(n5030));
  LUT5 #(.INIT(32'hFF969600)) lut_n5031 (.I0(x1623), .I1(x1624), .I2(x1625), .I3(n5029), .I4(n5030), .O(n5031));
  LUT3 #(.INIT(8'h96)) lut_n5032 (.I0(x1632), .I1(x1633), .I2(x1634), .O(n5032));
  LUT5 #(.INIT(32'h96696996)) lut_n5033 (.I0(x1623), .I1(x1624), .I2(x1625), .I3(n5029), .I4(n5030), .O(n5033));
  LUT5 #(.INIT(32'hFF969600)) lut_n5034 (.I0(x1629), .I1(x1630), .I2(x1631), .I3(n5032), .I4(n5033), .O(n5034));
  LUT3 #(.INIT(8'h96)) lut_n5035 (.I0(n5023), .I1(n5026), .I2(n5027), .O(n5035));
  LUT3 #(.INIT(8'hE8)) lut_n5036 (.I0(n5031), .I1(n5034), .I2(n5035), .O(n5036));
  LUT3 #(.INIT(8'h96)) lut_n5037 (.I0(n5006), .I1(n5014), .I2(n5015), .O(n5037));
  LUT3 #(.INIT(8'hE8)) lut_n5038 (.I0(n5028), .I1(n5036), .I2(n5037), .O(n5038));
  LUT3 #(.INIT(8'h96)) lut_n5039 (.I0(x1638), .I1(x1639), .I2(x1640), .O(n5039));
  LUT5 #(.INIT(32'h96696996)) lut_n5040 (.I0(x1629), .I1(x1630), .I2(x1631), .I3(n5032), .I4(n5033), .O(n5040));
  LUT5 #(.INIT(32'hFF969600)) lut_n5041 (.I0(x1635), .I1(x1636), .I2(x1637), .I3(n5039), .I4(n5040), .O(n5041));
  LUT3 #(.INIT(8'h96)) lut_n5042 (.I0(x1644), .I1(x1645), .I2(x1646), .O(n5042));
  LUT5 #(.INIT(32'h96696996)) lut_n5043 (.I0(x1635), .I1(x1636), .I2(x1637), .I3(n5039), .I4(n5040), .O(n5043));
  LUT5 #(.INIT(32'hFF969600)) lut_n5044 (.I0(x1641), .I1(x1642), .I2(x1643), .I3(n5042), .I4(n5043), .O(n5044));
  LUT3 #(.INIT(8'h96)) lut_n5045 (.I0(n5031), .I1(n5034), .I2(n5035), .O(n5045));
  LUT3 #(.INIT(8'hE8)) lut_n5046 (.I0(n5041), .I1(n5044), .I2(n5045), .O(n5046));
  LUT3 #(.INIT(8'h96)) lut_n5047 (.I0(x1650), .I1(x1651), .I2(x1652), .O(n5047));
  LUT5 #(.INIT(32'h96696996)) lut_n5048 (.I0(x1641), .I1(x1642), .I2(x1643), .I3(n5042), .I4(n5043), .O(n5048));
  LUT5 #(.INIT(32'hFF969600)) lut_n5049 (.I0(x1647), .I1(x1648), .I2(x1649), .I3(n5047), .I4(n5048), .O(n5049));
  LUT3 #(.INIT(8'h96)) lut_n5050 (.I0(x1656), .I1(x1657), .I2(x1658), .O(n5050));
  LUT5 #(.INIT(32'h96696996)) lut_n5051 (.I0(x1647), .I1(x1648), .I2(x1649), .I3(n5047), .I4(n5048), .O(n5051));
  LUT5 #(.INIT(32'hFF969600)) lut_n5052 (.I0(x1653), .I1(x1654), .I2(x1655), .I3(n5050), .I4(n5051), .O(n5052));
  LUT3 #(.INIT(8'h96)) lut_n5053 (.I0(n5041), .I1(n5044), .I2(n5045), .O(n5053));
  LUT3 #(.INIT(8'hE8)) lut_n5054 (.I0(n5049), .I1(n5052), .I2(n5053), .O(n5054));
  LUT3 #(.INIT(8'h96)) lut_n5055 (.I0(n5028), .I1(n5036), .I2(n5037), .O(n5055));
  LUT3 #(.INIT(8'hE8)) lut_n5056 (.I0(n5046), .I1(n5054), .I2(n5055), .O(n5056));
  LUT3 #(.INIT(8'h96)) lut_n5057 (.I0(n4998), .I1(n5016), .I2(n5017), .O(n5057));
  LUT3 #(.INIT(8'hE8)) lut_n5058 (.I0(n5038), .I1(n5056), .I2(n5057), .O(n5058));
  LUT3 #(.INIT(8'h96)) lut_n5059 (.I0(x1662), .I1(x1663), .I2(x1664), .O(n5059));
  LUT5 #(.INIT(32'h96696996)) lut_n5060 (.I0(x1653), .I1(x1654), .I2(x1655), .I3(n5050), .I4(n5051), .O(n5060));
  LUT5 #(.INIT(32'hFF969600)) lut_n5061 (.I0(x1659), .I1(x1660), .I2(x1661), .I3(n5059), .I4(n5060), .O(n5061));
  LUT3 #(.INIT(8'h96)) lut_n5062 (.I0(x1668), .I1(x1669), .I2(x1670), .O(n5062));
  LUT5 #(.INIT(32'h96696996)) lut_n5063 (.I0(x1659), .I1(x1660), .I2(x1661), .I3(n5059), .I4(n5060), .O(n5063));
  LUT5 #(.INIT(32'hFF969600)) lut_n5064 (.I0(x1665), .I1(x1666), .I2(x1667), .I3(n5062), .I4(n5063), .O(n5064));
  LUT3 #(.INIT(8'h96)) lut_n5065 (.I0(n5049), .I1(n5052), .I2(n5053), .O(n5065));
  LUT3 #(.INIT(8'hE8)) lut_n5066 (.I0(n5061), .I1(n5064), .I2(n5065), .O(n5066));
  LUT3 #(.INIT(8'h96)) lut_n5067 (.I0(x1674), .I1(x1675), .I2(x1676), .O(n5067));
  LUT5 #(.INIT(32'h96696996)) lut_n5068 (.I0(x1665), .I1(x1666), .I2(x1667), .I3(n5062), .I4(n5063), .O(n5068));
  LUT5 #(.INIT(32'hFF969600)) lut_n5069 (.I0(x1671), .I1(x1672), .I2(x1673), .I3(n5067), .I4(n5068), .O(n5069));
  LUT3 #(.INIT(8'h96)) lut_n5070 (.I0(x1680), .I1(x1681), .I2(x1682), .O(n5070));
  LUT5 #(.INIT(32'h96696996)) lut_n5071 (.I0(x1671), .I1(x1672), .I2(x1673), .I3(n5067), .I4(n5068), .O(n5071));
  LUT5 #(.INIT(32'hFF969600)) lut_n5072 (.I0(x1677), .I1(x1678), .I2(x1679), .I3(n5070), .I4(n5071), .O(n5072));
  LUT3 #(.INIT(8'h96)) lut_n5073 (.I0(n5061), .I1(n5064), .I2(n5065), .O(n5073));
  LUT3 #(.INIT(8'hE8)) lut_n5074 (.I0(n5069), .I1(n5072), .I2(n5073), .O(n5074));
  LUT3 #(.INIT(8'h96)) lut_n5075 (.I0(n5046), .I1(n5054), .I2(n5055), .O(n5075));
  LUT3 #(.INIT(8'hE8)) lut_n5076 (.I0(n5066), .I1(n5074), .I2(n5075), .O(n5076));
  LUT3 #(.INIT(8'h96)) lut_n5077 (.I0(x1686), .I1(x1687), .I2(x1688), .O(n5077));
  LUT5 #(.INIT(32'h96696996)) lut_n5078 (.I0(x1677), .I1(x1678), .I2(x1679), .I3(n5070), .I4(n5071), .O(n5078));
  LUT5 #(.INIT(32'hFF969600)) lut_n5079 (.I0(x1683), .I1(x1684), .I2(x1685), .I3(n5077), .I4(n5078), .O(n5079));
  LUT3 #(.INIT(8'h96)) lut_n5080 (.I0(x1692), .I1(x1693), .I2(x1694), .O(n5080));
  LUT5 #(.INIT(32'h96696996)) lut_n5081 (.I0(x1683), .I1(x1684), .I2(x1685), .I3(n5077), .I4(n5078), .O(n5081));
  LUT5 #(.INIT(32'hFF969600)) lut_n5082 (.I0(x1689), .I1(x1690), .I2(x1691), .I3(n5080), .I4(n5081), .O(n5082));
  LUT3 #(.INIT(8'h96)) lut_n5083 (.I0(n5069), .I1(n5072), .I2(n5073), .O(n5083));
  LUT3 #(.INIT(8'hE8)) lut_n5084 (.I0(n5079), .I1(n5082), .I2(n5083), .O(n5084));
  LUT3 #(.INIT(8'h96)) lut_n5085 (.I0(x1698), .I1(x1699), .I2(x1700), .O(n5085));
  LUT5 #(.INIT(32'h96696996)) lut_n5086 (.I0(x1689), .I1(x1690), .I2(x1691), .I3(n5080), .I4(n5081), .O(n5086));
  LUT5 #(.INIT(32'hFF969600)) lut_n5087 (.I0(x1695), .I1(x1696), .I2(x1697), .I3(n5085), .I4(n5086), .O(n5087));
  LUT3 #(.INIT(8'h96)) lut_n5088 (.I0(x1704), .I1(x1705), .I2(x1706), .O(n5088));
  LUT5 #(.INIT(32'h96696996)) lut_n5089 (.I0(x1695), .I1(x1696), .I2(x1697), .I3(n5085), .I4(n5086), .O(n5089));
  LUT5 #(.INIT(32'hFF969600)) lut_n5090 (.I0(x1701), .I1(x1702), .I2(x1703), .I3(n5088), .I4(n5089), .O(n5090));
  LUT3 #(.INIT(8'h96)) lut_n5091 (.I0(n5079), .I1(n5082), .I2(n5083), .O(n5091));
  LUT3 #(.INIT(8'hE8)) lut_n5092 (.I0(n5087), .I1(n5090), .I2(n5091), .O(n5092));
  LUT3 #(.INIT(8'h96)) lut_n5093 (.I0(n5066), .I1(n5074), .I2(n5075), .O(n5093));
  LUT3 #(.INIT(8'hE8)) lut_n5094 (.I0(n5084), .I1(n5092), .I2(n5093), .O(n5094));
  LUT3 #(.INIT(8'h96)) lut_n5095 (.I0(n5038), .I1(n5056), .I2(n5057), .O(n5095));
  LUT3 #(.INIT(8'hE8)) lut_n5096 (.I0(n5076), .I1(n5094), .I2(n5095), .O(n5096));
  LUT3 #(.INIT(8'h96)) lut_n5097 (.I0(n4980), .I1(n5018), .I2(n5019), .O(n5097));
  LUT3 #(.INIT(8'hE8)) lut_n5098 (.I0(n5058), .I1(n5096), .I2(n5097), .O(n5098));
  LUT3 #(.INIT(8'h96)) lut_n5099 (.I0(n4862), .I1(n4940), .I2(n4941), .O(n5099));
  LUT3 #(.INIT(8'hE8)) lut_n5100 (.I0(n5020), .I1(n5098), .I2(n5099), .O(n5100));
  LUT3 #(.INIT(8'h96)) lut_n5101 (.I0(n4622), .I1(n4780), .I2(n4781), .O(n5101));
  LUT3 #(.INIT(8'h96)) lut_n5102 (.I0(x1710), .I1(x1711), .I2(x1712), .O(n5102));
  LUT5 #(.INIT(32'h96696996)) lut_n5103 (.I0(x1701), .I1(x1702), .I2(x1703), .I3(n5088), .I4(n5089), .O(n5103));
  LUT5 #(.INIT(32'hFF969600)) lut_n5104 (.I0(x1707), .I1(x1708), .I2(x1709), .I3(n5102), .I4(n5103), .O(n5104));
  LUT3 #(.INIT(8'h96)) lut_n5105 (.I0(x1716), .I1(x1717), .I2(x1718), .O(n5105));
  LUT5 #(.INIT(32'h96696996)) lut_n5106 (.I0(x1707), .I1(x1708), .I2(x1709), .I3(n5102), .I4(n5103), .O(n5106));
  LUT5 #(.INIT(32'hFF969600)) lut_n5107 (.I0(x1713), .I1(x1714), .I2(x1715), .I3(n5105), .I4(n5106), .O(n5107));
  LUT3 #(.INIT(8'h96)) lut_n5108 (.I0(n5087), .I1(n5090), .I2(n5091), .O(n5108));
  LUT3 #(.INIT(8'hE8)) lut_n5109 (.I0(n5104), .I1(n5107), .I2(n5108), .O(n5109));
  LUT3 #(.INIT(8'h96)) lut_n5110 (.I0(x1722), .I1(x1723), .I2(x1724), .O(n5110));
  LUT5 #(.INIT(32'h96696996)) lut_n5111 (.I0(x1713), .I1(x1714), .I2(x1715), .I3(n5105), .I4(n5106), .O(n5111));
  LUT5 #(.INIT(32'hFF969600)) lut_n5112 (.I0(x1719), .I1(x1720), .I2(x1721), .I3(n5110), .I4(n5111), .O(n5112));
  LUT3 #(.INIT(8'h96)) lut_n5113 (.I0(x1728), .I1(x1729), .I2(x1730), .O(n5113));
  LUT5 #(.INIT(32'h96696996)) lut_n5114 (.I0(x1719), .I1(x1720), .I2(x1721), .I3(n5110), .I4(n5111), .O(n5114));
  LUT5 #(.INIT(32'hFF969600)) lut_n5115 (.I0(x1725), .I1(x1726), .I2(x1727), .I3(n5113), .I4(n5114), .O(n5115));
  LUT3 #(.INIT(8'h96)) lut_n5116 (.I0(n5104), .I1(n5107), .I2(n5108), .O(n5116));
  LUT3 #(.INIT(8'hE8)) lut_n5117 (.I0(n5112), .I1(n5115), .I2(n5116), .O(n5117));
  LUT3 #(.INIT(8'h96)) lut_n5118 (.I0(n5084), .I1(n5092), .I2(n5093), .O(n5118));
  LUT3 #(.INIT(8'hE8)) lut_n5119 (.I0(n5109), .I1(n5117), .I2(n5118), .O(n5119));
  LUT3 #(.INIT(8'h96)) lut_n5120 (.I0(x1734), .I1(x1735), .I2(x1736), .O(n5120));
  LUT5 #(.INIT(32'h96696996)) lut_n5121 (.I0(x1725), .I1(x1726), .I2(x1727), .I3(n5113), .I4(n5114), .O(n5121));
  LUT5 #(.INIT(32'hFF969600)) lut_n5122 (.I0(x1731), .I1(x1732), .I2(x1733), .I3(n5120), .I4(n5121), .O(n5122));
  LUT3 #(.INIT(8'h96)) lut_n5123 (.I0(x1740), .I1(x1741), .I2(x1742), .O(n5123));
  LUT5 #(.INIT(32'h96696996)) lut_n5124 (.I0(x1731), .I1(x1732), .I2(x1733), .I3(n5120), .I4(n5121), .O(n5124));
  LUT5 #(.INIT(32'hFF969600)) lut_n5125 (.I0(x1737), .I1(x1738), .I2(x1739), .I3(n5123), .I4(n5124), .O(n5125));
  LUT3 #(.INIT(8'h96)) lut_n5126 (.I0(n5112), .I1(n5115), .I2(n5116), .O(n5126));
  LUT3 #(.INIT(8'hE8)) lut_n5127 (.I0(n5122), .I1(n5125), .I2(n5126), .O(n5127));
  LUT3 #(.INIT(8'h96)) lut_n5128 (.I0(x1746), .I1(x1747), .I2(x1748), .O(n5128));
  LUT5 #(.INIT(32'h96696996)) lut_n5129 (.I0(x1737), .I1(x1738), .I2(x1739), .I3(n5123), .I4(n5124), .O(n5129));
  LUT5 #(.INIT(32'hFF969600)) lut_n5130 (.I0(x1743), .I1(x1744), .I2(x1745), .I3(n5128), .I4(n5129), .O(n5130));
  LUT3 #(.INIT(8'h96)) lut_n5131 (.I0(x1752), .I1(x1753), .I2(x1754), .O(n5131));
  LUT5 #(.INIT(32'h96696996)) lut_n5132 (.I0(x1743), .I1(x1744), .I2(x1745), .I3(n5128), .I4(n5129), .O(n5132));
  LUT5 #(.INIT(32'hFF969600)) lut_n5133 (.I0(x1749), .I1(x1750), .I2(x1751), .I3(n5131), .I4(n5132), .O(n5133));
  LUT3 #(.INIT(8'h96)) lut_n5134 (.I0(n5122), .I1(n5125), .I2(n5126), .O(n5134));
  LUT3 #(.INIT(8'hE8)) lut_n5135 (.I0(n5130), .I1(n5133), .I2(n5134), .O(n5135));
  LUT3 #(.INIT(8'h96)) lut_n5136 (.I0(n5109), .I1(n5117), .I2(n5118), .O(n5136));
  LUT3 #(.INIT(8'hE8)) lut_n5137 (.I0(n5127), .I1(n5135), .I2(n5136), .O(n5137));
  LUT3 #(.INIT(8'h96)) lut_n5138 (.I0(n5076), .I1(n5094), .I2(n5095), .O(n5138));
  LUT3 #(.INIT(8'hE8)) lut_n5139 (.I0(n5119), .I1(n5137), .I2(n5138), .O(n5139));
  LUT3 #(.INIT(8'h96)) lut_n5140 (.I0(x1758), .I1(x1759), .I2(x1760), .O(n5140));
  LUT5 #(.INIT(32'h96696996)) lut_n5141 (.I0(x1749), .I1(x1750), .I2(x1751), .I3(n5131), .I4(n5132), .O(n5141));
  LUT5 #(.INIT(32'hFF969600)) lut_n5142 (.I0(x1755), .I1(x1756), .I2(x1757), .I3(n5140), .I4(n5141), .O(n5142));
  LUT3 #(.INIT(8'h96)) lut_n5143 (.I0(x1764), .I1(x1765), .I2(x1766), .O(n5143));
  LUT5 #(.INIT(32'h96696996)) lut_n5144 (.I0(x1755), .I1(x1756), .I2(x1757), .I3(n5140), .I4(n5141), .O(n5144));
  LUT5 #(.INIT(32'hFF969600)) lut_n5145 (.I0(x1761), .I1(x1762), .I2(x1763), .I3(n5143), .I4(n5144), .O(n5145));
  LUT3 #(.INIT(8'h96)) lut_n5146 (.I0(n5130), .I1(n5133), .I2(n5134), .O(n5146));
  LUT3 #(.INIT(8'hE8)) lut_n5147 (.I0(n5142), .I1(n5145), .I2(n5146), .O(n5147));
  LUT3 #(.INIT(8'h96)) lut_n5148 (.I0(x1770), .I1(x1771), .I2(x1772), .O(n5148));
  LUT5 #(.INIT(32'h96696996)) lut_n5149 (.I0(x1761), .I1(x1762), .I2(x1763), .I3(n5143), .I4(n5144), .O(n5149));
  LUT5 #(.INIT(32'hFF969600)) lut_n5150 (.I0(x1767), .I1(x1768), .I2(x1769), .I3(n5148), .I4(n5149), .O(n5150));
  LUT3 #(.INIT(8'h96)) lut_n5151 (.I0(x1776), .I1(x1777), .I2(x1778), .O(n5151));
  LUT5 #(.INIT(32'h96696996)) lut_n5152 (.I0(x1767), .I1(x1768), .I2(x1769), .I3(n5148), .I4(n5149), .O(n5152));
  LUT5 #(.INIT(32'hFF969600)) lut_n5153 (.I0(x1773), .I1(x1774), .I2(x1775), .I3(n5151), .I4(n5152), .O(n5153));
  LUT3 #(.INIT(8'h96)) lut_n5154 (.I0(n5142), .I1(n5145), .I2(n5146), .O(n5154));
  LUT3 #(.INIT(8'hE8)) lut_n5155 (.I0(n5150), .I1(n5153), .I2(n5154), .O(n5155));
  LUT3 #(.INIT(8'h96)) lut_n5156 (.I0(n5127), .I1(n5135), .I2(n5136), .O(n5156));
  LUT3 #(.INIT(8'hE8)) lut_n5157 (.I0(n5147), .I1(n5155), .I2(n5156), .O(n5157));
  LUT3 #(.INIT(8'h96)) lut_n5158 (.I0(x1782), .I1(x1783), .I2(x1784), .O(n5158));
  LUT5 #(.INIT(32'h96696996)) lut_n5159 (.I0(x1773), .I1(x1774), .I2(x1775), .I3(n5151), .I4(n5152), .O(n5159));
  LUT5 #(.INIT(32'hFF969600)) lut_n5160 (.I0(x1779), .I1(x1780), .I2(x1781), .I3(n5158), .I4(n5159), .O(n5160));
  LUT3 #(.INIT(8'h96)) lut_n5161 (.I0(x1788), .I1(x1789), .I2(x1790), .O(n5161));
  LUT5 #(.INIT(32'h96696996)) lut_n5162 (.I0(x1779), .I1(x1780), .I2(x1781), .I3(n5158), .I4(n5159), .O(n5162));
  LUT5 #(.INIT(32'hFF969600)) lut_n5163 (.I0(x1785), .I1(x1786), .I2(x1787), .I3(n5161), .I4(n5162), .O(n5163));
  LUT3 #(.INIT(8'h96)) lut_n5164 (.I0(n5150), .I1(n5153), .I2(n5154), .O(n5164));
  LUT3 #(.INIT(8'hE8)) lut_n5165 (.I0(n5160), .I1(n5163), .I2(n5164), .O(n5165));
  LUT3 #(.INIT(8'h96)) lut_n5166 (.I0(x1794), .I1(x1795), .I2(x1796), .O(n5166));
  LUT5 #(.INIT(32'h96696996)) lut_n5167 (.I0(x1785), .I1(x1786), .I2(x1787), .I3(n5161), .I4(n5162), .O(n5167));
  LUT5 #(.INIT(32'hFF969600)) lut_n5168 (.I0(x1791), .I1(x1792), .I2(x1793), .I3(n5166), .I4(n5167), .O(n5168));
  LUT3 #(.INIT(8'h96)) lut_n5169 (.I0(x1800), .I1(x1801), .I2(x1802), .O(n5169));
  LUT5 #(.INIT(32'h96696996)) lut_n5170 (.I0(x1791), .I1(x1792), .I2(x1793), .I3(n5166), .I4(n5167), .O(n5170));
  LUT5 #(.INIT(32'hFF969600)) lut_n5171 (.I0(x1797), .I1(x1798), .I2(x1799), .I3(n5169), .I4(n5170), .O(n5171));
  LUT3 #(.INIT(8'h96)) lut_n5172 (.I0(n5160), .I1(n5163), .I2(n5164), .O(n5172));
  LUT3 #(.INIT(8'hE8)) lut_n5173 (.I0(n5168), .I1(n5171), .I2(n5172), .O(n5173));
  LUT3 #(.INIT(8'h96)) lut_n5174 (.I0(n5147), .I1(n5155), .I2(n5156), .O(n5174));
  LUT3 #(.INIT(8'hE8)) lut_n5175 (.I0(n5165), .I1(n5173), .I2(n5174), .O(n5175));
  LUT3 #(.INIT(8'h96)) lut_n5176 (.I0(n5119), .I1(n5137), .I2(n5138), .O(n5176));
  LUT3 #(.INIT(8'hE8)) lut_n5177 (.I0(n5157), .I1(n5175), .I2(n5176), .O(n5177));
  LUT3 #(.INIT(8'h96)) lut_n5178 (.I0(n5058), .I1(n5096), .I2(n5097), .O(n5178));
  LUT3 #(.INIT(8'hE8)) lut_n5179 (.I0(n5139), .I1(n5177), .I2(n5178), .O(n5179));
  LUT3 #(.INIT(8'h96)) lut_n5180 (.I0(x1806), .I1(x1807), .I2(x1808), .O(n5180));
  LUT5 #(.INIT(32'h96696996)) lut_n5181 (.I0(x1797), .I1(x1798), .I2(x1799), .I3(n5169), .I4(n5170), .O(n5181));
  LUT5 #(.INIT(32'hFF969600)) lut_n5182 (.I0(x1803), .I1(x1804), .I2(x1805), .I3(n5180), .I4(n5181), .O(n5182));
  LUT3 #(.INIT(8'h96)) lut_n5183 (.I0(x1812), .I1(x1813), .I2(x1814), .O(n5183));
  LUT5 #(.INIT(32'h96696996)) lut_n5184 (.I0(x1803), .I1(x1804), .I2(x1805), .I3(n5180), .I4(n5181), .O(n5184));
  LUT5 #(.INIT(32'hFF969600)) lut_n5185 (.I0(x1809), .I1(x1810), .I2(x1811), .I3(n5183), .I4(n5184), .O(n5185));
  LUT3 #(.INIT(8'h96)) lut_n5186 (.I0(n5168), .I1(n5171), .I2(n5172), .O(n5186));
  LUT3 #(.INIT(8'hE8)) lut_n5187 (.I0(n5182), .I1(n5185), .I2(n5186), .O(n5187));
  LUT3 #(.INIT(8'h96)) lut_n5188 (.I0(x1818), .I1(x1819), .I2(x1820), .O(n5188));
  LUT5 #(.INIT(32'h96696996)) lut_n5189 (.I0(x1809), .I1(x1810), .I2(x1811), .I3(n5183), .I4(n5184), .O(n5189));
  LUT5 #(.INIT(32'hFF969600)) lut_n5190 (.I0(x1815), .I1(x1816), .I2(x1817), .I3(n5188), .I4(n5189), .O(n5190));
  LUT3 #(.INIT(8'h96)) lut_n5191 (.I0(x1824), .I1(x1825), .I2(x1826), .O(n5191));
  LUT5 #(.INIT(32'h96696996)) lut_n5192 (.I0(x1815), .I1(x1816), .I2(x1817), .I3(n5188), .I4(n5189), .O(n5192));
  LUT5 #(.INIT(32'hFF969600)) lut_n5193 (.I0(x1821), .I1(x1822), .I2(x1823), .I3(n5191), .I4(n5192), .O(n5193));
  LUT3 #(.INIT(8'h96)) lut_n5194 (.I0(n5182), .I1(n5185), .I2(n5186), .O(n5194));
  LUT3 #(.INIT(8'hE8)) lut_n5195 (.I0(n5190), .I1(n5193), .I2(n5194), .O(n5195));
  LUT3 #(.INIT(8'h96)) lut_n5196 (.I0(n5165), .I1(n5173), .I2(n5174), .O(n5196));
  LUT3 #(.INIT(8'hE8)) lut_n5197 (.I0(n5187), .I1(n5195), .I2(n5196), .O(n5197));
  LUT3 #(.INIT(8'h96)) lut_n5198 (.I0(x1830), .I1(x1831), .I2(x1832), .O(n5198));
  LUT5 #(.INIT(32'h96696996)) lut_n5199 (.I0(x1821), .I1(x1822), .I2(x1823), .I3(n5191), .I4(n5192), .O(n5199));
  LUT5 #(.INIT(32'hFF969600)) lut_n5200 (.I0(x1827), .I1(x1828), .I2(x1829), .I3(n5198), .I4(n5199), .O(n5200));
  LUT3 #(.INIT(8'h96)) lut_n5201 (.I0(x1836), .I1(x1837), .I2(x1838), .O(n5201));
  LUT5 #(.INIT(32'h96696996)) lut_n5202 (.I0(x1827), .I1(x1828), .I2(x1829), .I3(n5198), .I4(n5199), .O(n5202));
  LUT5 #(.INIT(32'hFF969600)) lut_n5203 (.I0(x1833), .I1(x1834), .I2(x1835), .I3(n5201), .I4(n5202), .O(n5203));
  LUT3 #(.INIT(8'h96)) lut_n5204 (.I0(n5190), .I1(n5193), .I2(n5194), .O(n5204));
  LUT3 #(.INIT(8'hE8)) lut_n5205 (.I0(n5200), .I1(n5203), .I2(n5204), .O(n5205));
  LUT3 #(.INIT(8'h96)) lut_n5206 (.I0(x1842), .I1(x1843), .I2(x1844), .O(n5206));
  LUT5 #(.INIT(32'h96696996)) lut_n5207 (.I0(x1833), .I1(x1834), .I2(x1835), .I3(n5201), .I4(n5202), .O(n5207));
  LUT5 #(.INIT(32'hFF969600)) lut_n5208 (.I0(x1839), .I1(x1840), .I2(x1841), .I3(n5206), .I4(n5207), .O(n5208));
  LUT3 #(.INIT(8'h96)) lut_n5209 (.I0(x1848), .I1(x1849), .I2(x1850), .O(n5209));
  LUT5 #(.INIT(32'h96696996)) lut_n5210 (.I0(x1839), .I1(x1840), .I2(x1841), .I3(n5206), .I4(n5207), .O(n5210));
  LUT5 #(.INIT(32'hFF969600)) lut_n5211 (.I0(x1845), .I1(x1846), .I2(x1847), .I3(n5209), .I4(n5210), .O(n5211));
  LUT3 #(.INIT(8'h96)) lut_n5212 (.I0(n5200), .I1(n5203), .I2(n5204), .O(n5212));
  LUT3 #(.INIT(8'hE8)) lut_n5213 (.I0(n5208), .I1(n5211), .I2(n5212), .O(n5213));
  LUT3 #(.INIT(8'h96)) lut_n5214 (.I0(n5187), .I1(n5195), .I2(n5196), .O(n5214));
  LUT3 #(.INIT(8'hE8)) lut_n5215 (.I0(n5205), .I1(n5213), .I2(n5214), .O(n5215));
  LUT3 #(.INIT(8'h96)) lut_n5216 (.I0(n5157), .I1(n5175), .I2(n5176), .O(n5216));
  LUT3 #(.INIT(8'hE8)) lut_n5217 (.I0(n5197), .I1(n5215), .I2(n5216), .O(n5217));
  LUT3 #(.INIT(8'h96)) lut_n5218 (.I0(x1854), .I1(x1855), .I2(x1856), .O(n5218));
  LUT5 #(.INIT(32'h96696996)) lut_n5219 (.I0(x1845), .I1(x1846), .I2(x1847), .I3(n5209), .I4(n5210), .O(n5219));
  LUT5 #(.INIT(32'hFF969600)) lut_n5220 (.I0(x1851), .I1(x1852), .I2(x1853), .I3(n5218), .I4(n5219), .O(n5220));
  LUT3 #(.INIT(8'h96)) lut_n5221 (.I0(x1860), .I1(x1861), .I2(x1862), .O(n5221));
  LUT5 #(.INIT(32'h96696996)) lut_n5222 (.I0(x1851), .I1(x1852), .I2(x1853), .I3(n5218), .I4(n5219), .O(n5222));
  LUT5 #(.INIT(32'hFF969600)) lut_n5223 (.I0(x1857), .I1(x1858), .I2(x1859), .I3(n5221), .I4(n5222), .O(n5223));
  LUT3 #(.INIT(8'h96)) lut_n5224 (.I0(n5208), .I1(n5211), .I2(n5212), .O(n5224));
  LUT3 #(.INIT(8'hE8)) lut_n5225 (.I0(n5220), .I1(n5223), .I2(n5224), .O(n5225));
  LUT3 #(.INIT(8'h96)) lut_n5226 (.I0(x1866), .I1(x1867), .I2(x1868), .O(n5226));
  LUT5 #(.INIT(32'h96696996)) lut_n5227 (.I0(x1857), .I1(x1858), .I2(x1859), .I3(n5221), .I4(n5222), .O(n5227));
  LUT5 #(.INIT(32'hFF969600)) lut_n5228 (.I0(x1863), .I1(x1864), .I2(x1865), .I3(n5226), .I4(n5227), .O(n5228));
  LUT3 #(.INIT(8'h96)) lut_n5229 (.I0(x1872), .I1(x1873), .I2(x1874), .O(n5229));
  LUT5 #(.INIT(32'h96696996)) lut_n5230 (.I0(x1863), .I1(x1864), .I2(x1865), .I3(n5226), .I4(n5227), .O(n5230));
  LUT5 #(.INIT(32'hFF969600)) lut_n5231 (.I0(x1869), .I1(x1870), .I2(x1871), .I3(n5229), .I4(n5230), .O(n5231));
  LUT3 #(.INIT(8'h96)) lut_n5232 (.I0(n5220), .I1(n5223), .I2(n5224), .O(n5232));
  LUT3 #(.INIT(8'hE8)) lut_n5233 (.I0(n5228), .I1(n5231), .I2(n5232), .O(n5233));
  LUT3 #(.INIT(8'h96)) lut_n5234 (.I0(n5205), .I1(n5213), .I2(n5214), .O(n5234));
  LUT3 #(.INIT(8'hE8)) lut_n5235 (.I0(n5225), .I1(n5233), .I2(n5234), .O(n5235));
  LUT3 #(.INIT(8'h96)) lut_n5236 (.I0(x1878), .I1(x1879), .I2(x1880), .O(n5236));
  LUT5 #(.INIT(32'h96696996)) lut_n5237 (.I0(x1869), .I1(x1870), .I2(x1871), .I3(n5229), .I4(n5230), .O(n5237));
  LUT5 #(.INIT(32'hFF969600)) lut_n5238 (.I0(x1875), .I1(x1876), .I2(x1877), .I3(n5236), .I4(n5237), .O(n5238));
  LUT3 #(.INIT(8'h96)) lut_n5239 (.I0(x1884), .I1(x1885), .I2(x1886), .O(n5239));
  LUT5 #(.INIT(32'h96696996)) lut_n5240 (.I0(x1875), .I1(x1876), .I2(x1877), .I3(n5236), .I4(n5237), .O(n5240));
  LUT5 #(.INIT(32'hFF969600)) lut_n5241 (.I0(x1881), .I1(x1882), .I2(x1883), .I3(n5239), .I4(n5240), .O(n5241));
  LUT3 #(.INIT(8'h96)) lut_n5242 (.I0(n5228), .I1(n5231), .I2(n5232), .O(n5242));
  LUT3 #(.INIT(8'hE8)) lut_n5243 (.I0(n5238), .I1(n5241), .I2(n5242), .O(n5243));
  LUT3 #(.INIT(8'h96)) lut_n5244 (.I0(x1890), .I1(x1891), .I2(x1892), .O(n5244));
  LUT5 #(.INIT(32'h96696996)) lut_n5245 (.I0(x1881), .I1(x1882), .I2(x1883), .I3(n5239), .I4(n5240), .O(n5245));
  LUT5 #(.INIT(32'hFF969600)) lut_n5246 (.I0(x1887), .I1(x1888), .I2(x1889), .I3(n5244), .I4(n5245), .O(n5246));
  LUT3 #(.INIT(8'h96)) lut_n5247 (.I0(x1896), .I1(x1897), .I2(x1898), .O(n5247));
  LUT5 #(.INIT(32'h96696996)) lut_n5248 (.I0(x1887), .I1(x1888), .I2(x1889), .I3(n5244), .I4(n5245), .O(n5248));
  LUT5 #(.INIT(32'hFF969600)) lut_n5249 (.I0(x1893), .I1(x1894), .I2(x1895), .I3(n5247), .I4(n5248), .O(n5249));
  LUT3 #(.INIT(8'h96)) lut_n5250 (.I0(n5238), .I1(n5241), .I2(n5242), .O(n5250));
  LUT3 #(.INIT(8'hE8)) lut_n5251 (.I0(n5246), .I1(n5249), .I2(n5250), .O(n5251));
  LUT3 #(.INIT(8'h96)) lut_n5252 (.I0(n5225), .I1(n5233), .I2(n5234), .O(n5252));
  LUT3 #(.INIT(8'hE8)) lut_n5253 (.I0(n5243), .I1(n5251), .I2(n5252), .O(n5253));
  LUT3 #(.INIT(8'h96)) lut_n5254 (.I0(n5197), .I1(n5215), .I2(n5216), .O(n5254));
  LUT3 #(.INIT(8'hE8)) lut_n5255 (.I0(n5235), .I1(n5253), .I2(n5254), .O(n5255));
  LUT3 #(.INIT(8'h96)) lut_n5256 (.I0(n5139), .I1(n5177), .I2(n5178), .O(n5256));
  LUT3 #(.INIT(8'hE8)) lut_n5257 (.I0(n5217), .I1(n5255), .I2(n5256), .O(n5257));
  LUT3 #(.INIT(8'h96)) lut_n5258 (.I0(n5020), .I1(n5098), .I2(n5099), .O(n5258));
  LUT3 #(.INIT(8'hE8)) lut_n5259 (.I0(n5179), .I1(n5257), .I2(n5258), .O(n5259));
  LUT3 #(.INIT(8'h96)) lut_n5260 (.I0(x1902), .I1(x1903), .I2(x1904), .O(n5260));
  LUT5 #(.INIT(32'h96696996)) lut_n5261 (.I0(x1893), .I1(x1894), .I2(x1895), .I3(n5247), .I4(n5248), .O(n5261));
  LUT5 #(.INIT(32'hFF969600)) lut_n5262 (.I0(x1899), .I1(x1900), .I2(x1901), .I3(n5260), .I4(n5261), .O(n5262));
  LUT3 #(.INIT(8'h96)) lut_n5263 (.I0(x1908), .I1(x1909), .I2(x1910), .O(n5263));
  LUT5 #(.INIT(32'h96696996)) lut_n5264 (.I0(x1899), .I1(x1900), .I2(x1901), .I3(n5260), .I4(n5261), .O(n5264));
  LUT5 #(.INIT(32'hFF969600)) lut_n5265 (.I0(x1905), .I1(x1906), .I2(x1907), .I3(n5263), .I4(n5264), .O(n5265));
  LUT3 #(.INIT(8'h96)) lut_n5266 (.I0(n5246), .I1(n5249), .I2(n5250), .O(n5266));
  LUT3 #(.INIT(8'hE8)) lut_n5267 (.I0(n5262), .I1(n5265), .I2(n5266), .O(n5267));
  LUT3 #(.INIT(8'h96)) lut_n5268 (.I0(x1914), .I1(x1915), .I2(x1916), .O(n5268));
  LUT5 #(.INIT(32'h96696996)) lut_n5269 (.I0(x1905), .I1(x1906), .I2(x1907), .I3(n5263), .I4(n5264), .O(n5269));
  LUT5 #(.INIT(32'hFF969600)) lut_n5270 (.I0(x1911), .I1(x1912), .I2(x1913), .I3(n5268), .I4(n5269), .O(n5270));
  LUT3 #(.INIT(8'h96)) lut_n5271 (.I0(x1920), .I1(x1921), .I2(x1922), .O(n5271));
  LUT5 #(.INIT(32'h96696996)) lut_n5272 (.I0(x1911), .I1(x1912), .I2(x1913), .I3(n5268), .I4(n5269), .O(n5272));
  LUT5 #(.INIT(32'hFF969600)) lut_n5273 (.I0(x1917), .I1(x1918), .I2(x1919), .I3(n5271), .I4(n5272), .O(n5273));
  LUT3 #(.INIT(8'h96)) lut_n5274 (.I0(n5262), .I1(n5265), .I2(n5266), .O(n5274));
  LUT3 #(.INIT(8'hE8)) lut_n5275 (.I0(n5270), .I1(n5273), .I2(n5274), .O(n5275));
  LUT3 #(.INIT(8'h96)) lut_n5276 (.I0(n5243), .I1(n5251), .I2(n5252), .O(n5276));
  LUT3 #(.INIT(8'hE8)) lut_n5277 (.I0(n5267), .I1(n5275), .I2(n5276), .O(n5277));
  LUT3 #(.INIT(8'h96)) lut_n5278 (.I0(x1926), .I1(x1927), .I2(x1928), .O(n5278));
  LUT5 #(.INIT(32'h96696996)) lut_n5279 (.I0(x1917), .I1(x1918), .I2(x1919), .I3(n5271), .I4(n5272), .O(n5279));
  LUT5 #(.INIT(32'hFF969600)) lut_n5280 (.I0(x1923), .I1(x1924), .I2(x1925), .I3(n5278), .I4(n5279), .O(n5280));
  LUT3 #(.INIT(8'h96)) lut_n5281 (.I0(x1932), .I1(x1933), .I2(x1934), .O(n5281));
  LUT5 #(.INIT(32'h96696996)) lut_n5282 (.I0(x1923), .I1(x1924), .I2(x1925), .I3(n5278), .I4(n5279), .O(n5282));
  LUT5 #(.INIT(32'hFF969600)) lut_n5283 (.I0(x1929), .I1(x1930), .I2(x1931), .I3(n5281), .I4(n5282), .O(n5283));
  LUT3 #(.INIT(8'h96)) lut_n5284 (.I0(n5270), .I1(n5273), .I2(n5274), .O(n5284));
  LUT3 #(.INIT(8'hE8)) lut_n5285 (.I0(n5280), .I1(n5283), .I2(n5284), .O(n5285));
  LUT3 #(.INIT(8'h96)) lut_n5286 (.I0(x1938), .I1(x1939), .I2(x1940), .O(n5286));
  LUT5 #(.INIT(32'h96696996)) lut_n5287 (.I0(x1929), .I1(x1930), .I2(x1931), .I3(n5281), .I4(n5282), .O(n5287));
  LUT5 #(.INIT(32'hFF969600)) lut_n5288 (.I0(x1935), .I1(x1936), .I2(x1937), .I3(n5286), .I4(n5287), .O(n5288));
  LUT3 #(.INIT(8'h96)) lut_n5289 (.I0(x1944), .I1(x1945), .I2(x1946), .O(n5289));
  LUT5 #(.INIT(32'h96696996)) lut_n5290 (.I0(x1935), .I1(x1936), .I2(x1937), .I3(n5286), .I4(n5287), .O(n5290));
  LUT5 #(.INIT(32'hFF969600)) lut_n5291 (.I0(x1941), .I1(x1942), .I2(x1943), .I3(n5289), .I4(n5290), .O(n5291));
  LUT3 #(.INIT(8'h96)) lut_n5292 (.I0(n5280), .I1(n5283), .I2(n5284), .O(n5292));
  LUT3 #(.INIT(8'hE8)) lut_n5293 (.I0(n5288), .I1(n5291), .I2(n5292), .O(n5293));
  LUT3 #(.INIT(8'h96)) lut_n5294 (.I0(n5267), .I1(n5275), .I2(n5276), .O(n5294));
  LUT3 #(.INIT(8'hE8)) lut_n5295 (.I0(n5285), .I1(n5293), .I2(n5294), .O(n5295));
  LUT3 #(.INIT(8'h96)) lut_n5296 (.I0(n5235), .I1(n5253), .I2(n5254), .O(n5296));
  LUT3 #(.INIT(8'hE8)) lut_n5297 (.I0(n5277), .I1(n5295), .I2(n5296), .O(n5297));
  LUT3 #(.INIT(8'h96)) lut_n5298 (.I0(x1950), .I1(x1951), .I2(x1952), .O(n5298));
  LUT5 #(.INIT(32'h96696996)) lut_n5299 (.I0(x1941), .I1(x1942), .I2(x1943), .I3(n5289), .I4(n5290), .O(n5299));
  LUT5 #(.INIT(32'hFF969600)) lut_n5300 (.I0(x1947), .I1(x1948), .I2(x1949), .I3(n5298), .I4(n5299), .O(n5300));
  LUT3 #(.INIT(8'h96)) lut_n5301 (.I0(x1956), .I1(x1957), .I2(x1958), .O(n5301));
  LUT5 #(.INIT(32'h96696996)) lut_n5302 (.I0(x1947), .I1(x1948), .I2(x1949), .I3(n5298), .I4(n5299), .O(n5302));
  LUT5 #(.INIT(32'hFF969600)) lut_n5303 (.I0(x1953), .I1(x1954), .I2(x1955), .I3(n5301), .I4(n5302), .O(n5303));
  LUT3 #(.INIT(8'h96)) lut_n5304 (.I0(n5288), .I1(n5291), .I2(n5292), .O(n5304));
  LUT3 #(.INIT(8'hE8)) lut_n5305 (.I0(n5300), .I1(n5303), .I2(n5304), .O(n5305));
  LUT3 #(.INIT(8'h96)) lut_n5306 (.I0(x1962), .I1(x1963), .I2(x1964), .O(n5306));
  LUT5 #(.INIT(32'h96696996)) lut_n5307 (.I0(x1953), .I1(x1954), .I2(x1955), .I3(n5301), .I4(n5302), .O(n5307));
  LUT5 #(.INIT(32'hFF969600)) lut_n5308 (.I0(x1959), .I1(x1960), .I2(x1961), .I3(n5306), .I4(n5307), .O(n5308));
  LUT3 #(.INIT(8'h96)) lut_n5309 (.I0(x1968), .I1(x1969), .I2(x1970), .O(n5309));
  LUT5 #(.INIT(32'h96696996)) lut_n5310 (.I0(x1959), .I1(x1960), .I2(x1961), .I3(n5306), .I4(n5307), .O(n5310));
  LUT5 #(.INIT(32'hFF969600)) lut_n5311 (.I0(x1965), .I1(x1966), .I2(x1967), .I3(n5309), .I4(n5310), .O(n5311));
  LUT3 #(.INIT(8'h96)) lut_n5312 (.I0(n5300), .I1(n5303), .I2(n5304), .O(n5312));
  LUT3 #(.INIT(8'hE8)) lut_n5313 (.I0(n5308), .I1(n5311), .I2(n5312), .O(n5313));
  LUT3 #(.INIT(8'h96)) lut_n5314 (.I0(n5285), .I1(n5293), .I2(n5294), .O(n5314));
  LUT3 #(.INIT(8'hE8)) lut_n5315 (.I0(n5305), .I1(n5313), .I2(n5314), .O(n5315));
  LUT3 #(.INIT(8'h96)) lut_n5316 (.I0(x1974), .I1(x1975), .I2(x1976), .O(n5316));
  LUT5 #(.INIT(32'h96696996)) lut_n5317 (.I0(x1965), .I1(x1966), .I2(x1967), .I3(n5309), .I4(n5310), .O(n5317));
  LUT5 #(.INIT(32'hFF969600)) lut_n5318 (.I0(x1971), .I1(x1972), .I2(x1973), .I3(n5316), .I4(n5317), .O(n5318));
  LUT3 #(.INIT(8'h96)) lut_n5319 (.I0(x1980), .I1(x1981), .I2(x1982), .O(n5319));
  LUT5 #(.INIT(32'h96696996)) lut_n5320 (.I0(x1971), .I1(x1972), .I2(x1973), .I3(n5316), .I4(n5317), .O(n5320));
  LUT5 #(.INIT(32'hFF969600)) lut_n5321 (.I0(x1977), .I1(x1978), .I2(x1979), .I3(n5319), .I4(n5320), .O(n5321));
  LUT3 #(.INIT(8'h96)) lut_n5322 (.I0(n5308), .I1(n5311), .I2(n5312), .O(n5322));
  LUT3 #(.INIT(8'hE8)) lut_n5323 (.I0(n5318), .I1(n5321), .I2(n5322), .O(n5323));
  LUT3 #(.INIT(8'h96)) lut_n5324 (.I0(x1986), .I1(x1987), .I2(x1988), .O(n5324));
  LUT5 #(.INIT(32'h96696996)) lut_n5325 (.I0(x1977), .I1(x1978), .I2(x1979), .I3(n5319), .I4(n5320), .O(n5325));
  LUT5 #(.INIT(32'hFF969600)) lut_n5326 (.I0(x1983), .I1(x1984), .I2(x1985), .I3(n5324), .I4(n5325), .O(n5326));
  LUT3 #(.INIT(8'h96)) lut_n5327 (.I0(x1992), .I1(x1993), .I2(x1994), .O(n5327));
  LUT5 #(.INIT(32'h96696996)) lut_n5328 (.I0(x1983), .I1(x1984), .I2(x1985), .I3(n5324), .I4(n5325), .O(n5328));
  LUT5 #(.INIT(32'hFF969600)) lut_n5329 (.I0(x1989), .I1(x1990), .I2(x1991), .I3(n5327), .I4(n5328), .O(n5329));
  LUT3 #(.INIT(8'h96)) lut_n5330 (.I0(n5318), .I1(n5321), .I2(n5322), .O(n5330));
  LUT3 #(.INIT(8'hE8)) lut_n5331 (.I0(n5326), .I1(n5329), .I2(n5330), .O(n5331));
  LUT3 #(.INIT(8'h96)) lut_n5332 (.I0(n5305), .I1(n5313), .I2(n5314), .O(n5332));
  LUT3 #(.INIT(8'hE8)) lut_n5333 (.I0(n5323), .I1(n5331), .I2(n5332), .O(n5333));
  LUT3 #(.INIT(8'h96)) lut_n5334 (.I0(n5277), .I1(n5295), .I2(n5296), .O(n5334));
  LUT3 #(.INIT(8'hE8)) lut_n5335 (.I0(n5315), .I1(n5333), .I2(n5334), .O(n5335));
  LUT3 #(.INIT(8'h96)) lut_n5336 (.I0(n5217), .I1(n5255), .I2(n5256), .O(n5336));
  LUT3 #(.INIT(8'hE8)) lut_n5337 (.I0(n5297), .I1(n5335), .I2(n5336), .O(n5337));
  LUT3 #(.INIT(8'h96)) lut_n5338 (.I0(x1998), .I1(x1999), .I2(x2000), .O(n5338));
  LUT5 #(.INIT(32'h96696996)) lut_n5339 (.I0(x1989), .I1(x1990), .I2(x1991), .I3(n5327), .I4(n5328), .O(n5339));
  LUT5 #(.INIT(32'hFF969600)) lut_n5340 (.I0(x1995), .I1(x1996), .I2(x1997), .I3(n5338), .I4(n5339), .O(n5340));
  LUT3 #(.INIT(8'h96)) lut_n5341 (.I0(x2004), .I1(x2005), .I2(x2006), .O(n5341));
  LUT5 #(.INIT(32'h96696996)) lut_n5342 (.I0(x1995), .I1(x1996), .I2(x1997), .I3(n5338), .I4(n5339), .O(n5342));
  LUT5 #(.INIT(32'hFF969600)) lut_n5343 (.I0(x2001), .I1(x2002), .I2(x2003), .I3(n5341), .I4(n5342), .O(n5343));
  LUT3 #(.INIT(8'h96)) lut_n5344 (.I0(n5326), .I1(n5329), .I2(n5330), .O(n5344));
  LUT3 #(.INIT(8'hE8)) lut_n5345 (.I0(n5340), .I1(n5343), .I2(n5344), .O(n5345));
  LUT3 #(.INIT(8'h96)) lut_n5346 (.I0(x2010), .I1(x2011), .I2(x2012), .O(n5346));
  LUT5 #(.INIT(32'h96696996)) lut_n5347 (.I0(x2001), .I1(x2002), .I2(x2003), .I3(n5341), .I4(n5342), .O(n5347));
  LUT5 #(.INIT(32'hFF969600)) lut_n5348 (.I0(x2007), .I1(x2008), .I2(x2009), .I3(n5346), .I4(n5347), .O(n5348));
  LUT3 #(.INIT(8'h96)) lut_n5349 (.I0(x2016), .I1(x2017), .I2(x2018), .O(n5349));
  LUT5 #(.INIT(32'h96696996)) lut_n5350 (.I0(x2007), .I1(x2008), .I2(x2009), .I3(n5346), .I4(n5347), .O(n5350));
  LUT5 #(.INIT(32'hFF969600)) lut_n5351 (.I0(x2013), .I1(x2014), .I2(x2015), .I3(n5349), .I4(n5350), .O(n5351));
  LUT3 #(.INIT(8'h96)) lut_n5352 (.I0(n5340), .I1(n5343), .I2(n5344), .O(n5352));
  LUT3 #(.INIT(8'hE8)) lut_n5353 (.I0(n5348), .I1(n5351), .I2(n5352), .O(n5353));
  LUT3 #(.INIT(8'h96)) lut_n5354 (.I0(n5323), .I1(n5331), .I2(n5332), .O(n5354));
  LUT3 #(.INIT(8'hE8)) lut_n5355 (.I0(n5345), .I1(n5353), .I2(n5354), .O(n5355));
  LUT3 #(.INIT(8'h96)) lut_n5356 (.I0(x2022), .I1(x2023), .I2(x2024), .O(n5356));
  LUT5 #(.INIT(32'h96696996)) lut_n5357 (.I0(x2013), .I1(x2014), .I2(x2015), .I3(n5349), .I4(n5350), .O(n5357));
  LUT5 #(.INIT(32'hFF969600)) lut_n5358 (.I0(x2019), .I1(x2020), .I2(x2021), .I3(n5356), .I4(n5357), .O(n5358));
  LUT5 #(.INIT(32'h96696996)) lut_n5359 (.I0(x2019), .I1(x2020), .I2(x2021), .I3(n5356), .I4(n5357), .O(n5359));
  LUT3 #(.INIT(8'h96)) lut_n5360 (.I0(n5348), .I1(n5351), .I2(n5352), .O(n5360));
  LUT6 #(.INIT(64'hFF96969696969600)) lut_n5361 (.I0(n5345), .I1(n5353), .I2(n5354), .I3(n5358), .I4(n5359), .I5(n5360), .O(n5361));
  LUT3 #(.INIT(8'h96)) lut_n5362 (.I0(n5315), .I1(n5333), .I2(n5334), .O(n5362));
  LUT6 #(.INIT(64'hFF96969696969600)) lut_n5363 (.I0(n5297), .I1(n5335), .I2(n5336), .I3(n5355), .I4(n5361), .I5(n5362), .O(n5363));
  LUT5 #(.INIT(32'hFF969600)) lut_n5364 (.I0(n5179), .I1(n5257), .I2(n5258), .I3(n5337), .I4(n5363), .O(n5364));
  LUT3 #(.INIT(8'h96)) lut_n5365 (.I0(n4464), .I1(n4782), .I2(n4783), .O(n5365));
  LUT6 #(.INIT(64'hFFFEFEE8E8808000)) lut_n5366 (.I0(n4942), .I1(n5100), .I2(n5101), .I3(n5259), .I4(n5364), .I5(n5365), .O(n5366));
  LUT5 #(.INIT(32'hFF969600)) lut_n5367 (.I0(n3596), .I1(n4144), .I2(n4145), .I3(n4784), .I4(n5366), .O(n5367));
  LUT3 #(.INIT(8'hE8)) lut_n5368 (.I0(n3278), .I1(n4146), .I2(n5367), .O(n5368));
  assign y0 = n5368;
endmodule
