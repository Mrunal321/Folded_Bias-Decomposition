module top (x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, y0);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24;
  output y0;
  wire n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56;
  LUT3 #(.INIT(8'hE8)) lut_n27 (.I0(x0), .I1(x1), .I2(x2), .O(n27));
  LUT3 #(.INIT(8'hE8)) lut_n28 (.I0(x6), .I1(x7), .I2(x8), .O(n28));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n29 (.I0(x3), .I1(x4), .I2(x5), .I3(n27), .I4(n28), .O(n29));
  LUT3 #(.INIT(8'hE8)) lut_n30 (.I0(x12), .I1(x13), .I2(x14), .O(n30));
  LUT5 #(.INIT(32'hE81717E8)) lut_n31 (.I0(x3), .I1(x4), .I2(x5), .I3(n27), .I4(n28), .O(n31));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n32 (.I0(x9), .I1(x10), .I2(x11), .I3(n30), .I4(n31), .O(n32));
  LUT3 #(.INIT(8'hE8)) lut_n33 (.I0(x18), .I1(x19), .I2(x20), .O(n33));
  LUT5 #(.INIT(32'hE81717E8)) lut_n34 (.I0(x9), .I1(x10), .I2(x11), .I3(n30), .I4(n31), .O(n34));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n35 (.I0(x15), .I1(x16), .I2(x17), .I3(n33), .I4(n34), .O(n35));
  LUT3 #(.INIT(8'hE8)) lut_n36 (.I0(n29), .I1(n32), .I2(n35), .O(n36));
  LUT5 #(.INIT(32'hE81717E8)) lut_n37 (.I0(x15), .I1(x16), .I2(x17), .I3(n33), .I4(n34), .O(n37));
  LUT4 #(.INIT(16'hFFE8)) lut_n38 (.I0(x21), .I1(x22), .I2(x23), .I3(n37), .O(n38));
  LUT3 #(.INIT(8'h96)) lut_n39 (.I0(x0), .I1(x1), .I2(x2), .O(n39));
  LUT3 #(.INIT(8'h96)) lut_n40 (.I0(x6), .I1(x7), .I2(x8), .O(n40));
  LUT5 #(.INIT(32'hFF969600)) lut_n41 (.I0(x3), .I1(x4), .I2(x5), .I3(n39), .I4(n40), .O(n41));
  LUT4 #(.INIT(16'h17E8)) lut_n42 (.I0(x21), .I1(x22), .I2(x23), .I3(n37), .O(n42));
  LUT2 #(.INIT(4'h2)) lut_n43 (.I0(n41), .I1(n42), .O(n43));
  LUT3 #(.INIT(8'h96)) lut_n44 (.I0(n29), .I1(n32), .I2(n35), .O(n44));
  LUT3 #(.INIT(8'h96)) lut_n45 (.I0(x12), .I1(x13), .I2(x14), .O(n45));
  LUT5 #(.INIT(32'h96696996)) lut_n46 (.I0(x3), .I1(x4), .I2(x5), .I3(n39), .I4(n40), .O(n46));
  LUT5 #(.INIT(32'hFF969600)) lut_n47 (.I0(x9), .I1(x10), .I2(x11), .I3(n45), .I4(n46), .O(n47));
  LUT3 #(.INIT(8'h96)) lut_n48 (.I0(x18), .I1(x19), .I2(x20), .O(n48));
  LUT5 #(.INIT(32'h96696996)) lut_n49 (.I0(x9), .I1(x10), .I2(x11), .I3(n45), .I4(n46), .O(n49));
  LUT5 #(.INIT(32'hFF969600)) lut_n50 (.I0(x15), .I1(x16), .I2(x17), .I3(n48), .I4(n49), .O(n50));
  LUT2 #(.INIT(4'h6)) lut_n51 (.I0(n41), .I1(n42), .O(n51));
  LUT3 #(.INIT(8'h8E)) lut_n52 (.I0(n47), .I1(n50), .I2(n51), .O(n52));
  LUT3 #(.INIT(8'h96)) lut_n53 (.I0(x21), .I1(x22), .I2(x23), .O(n53));
  LUT5 #(.INIT(32'h96696996)) lut_n54 (.I0(x15), .I1(x16), .I2(x17), .I3(n48), .I4(n49), .O(n54));
  LUT6 #(.INIT(64'hBEEB3CC33CC32882)) lut_n55 (.I0(x24), .I1(n47), .I2(n50), .I3(n51), .I4(n53), .I5(n54), .O(n55));
  LUT6 #(.INIT(64'hFEEAEAA8EAA8A880)) lut_n56 (.I0(n36), .I1(n38), .I2(n43), .I3(n44), .I4(n52), .I5(n55), .O(n56));
  assign y0 = n56;
endmodule
