module top (x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, y0);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254;
  output y0;
  wire n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650;
  LUT3 #(.INIT(8'hE8)) lut_n257 (.I0(x0), .I1(x1), .I2(x2), .O(n257));
  LUT3 #(.INIT(8'hE8)) lut_n258 (.I0(x6), .I1(x7), .I2(x8), .O(n258));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n259 (.I0(x3), .I1(x4), .I2(x5), .I3(n257), .I4(n258), .O(n259));
  LUT3 #(.INIT(8'hE8)) lut_n260 (.I0(x12), .I1(x13), .I2(x14), .O(n260));
  LUT5 #(.INIT(32'hE81717E8)) lut_n261 (.I0(x3), .I1(x4), .I2(x5), .I3(n257), .I4(n258), .O(n261));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n262 (.I0(x9), .I1(x10), .I2(x11), .I3(n260), .I4(n261), .O(n262));
  LUT3 #(.INIT(8'hE8)) lut_n263 (.I0(x18), .I1(x19), .I2(x20), .O(n263));
  LUT5 #(.INIT(32'hE81717E8)) lut_n264 (.I0(x9), .I1(x10), .I2(x11), .I3(n260), .I4(n261), .O(n264));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n265 (.I0(x15), .I1(x16), .I2(x17), .I3(n263), .I4(n264), .O(n265));
  LUT3 #(.INIT(8'hE8)) lut_n266 (.I0(n259), .I1(n262), .I2(n265), .O(n266));
  LUT3 #(.INIT(8'hE8)) lut_n267 (.I0(x24), .I1(x25), .I2(x26), .O(n267));
  LUT5 #(.INIT(32'hE81717E8)) lut_n268 (.I0(x15), .I1(x16), .I2(x17), .I3(n263), .I4(n264), .O(n268));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n269 (.I0(x21), .I1(x22), .I2(x23), .I3(n267), .I4(n268), .O(n269));
  LUT3 #(.INIT(8'hE8)) lut_n270 (.I0(x27), .I1(x28), .I2(x29), .O(n270));
  LUT5 #(.INIT(32'hE81717E8)) lut_n271 (.I0(x21), .I1(x22), .I2(x23), .I3(n267), .I4(n268), .O(n271));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n272 (.I0(x30), .I1(x31), .I2(x32), .I3(n270), .I4(n271), .O(n272));
  LUT3 #(.INIT(8'h96)) lut_n273 (.I0(n259), .I1(n262), .I2(n265), .O(n273));
  LUT3 #(.INIT(8'hE8)) lut_n274 (.I0(n269), .I1(n272), .I2(n273), .O(n274));
  LUT3 #(.INIT(8'hE8)) lut_n275 (.I0(x36), .I1(x37), .I2(x38), .O(n275));
  LUT5 #(.INIT(32'hE81717E8)) lut_n276 (.I0(x30), .I1(x31), .I2(x32), .I3(n270), .I4(n271), .O(n276));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n277 (.I0(x33), .I1(x34), .I2(x35), .I3(n275), .I4(n276), .O(n277));
  LUT3 #(.INIT(8'hE8)) lut_n278 (.I0(x42), .I1(x43), .I2(x44), .O(n278));
  LUT5 #(.INIT(32'hE81717E8)) lut_n279 (.I0(x33), .I1(x34), .I2(x35), .I3(n275), .I4(n276), .O(n279));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n280 (.I0(x39), .I1(x40), .I2(x41), .I3(n278), .I4(n279), .O(n280));
  LUT3 #(.INIT(8'h96)) lut_n281 (.I0(n269), .I1(n272), .I2(n273), .O(n281));
  LUT3 #(.INIT(8'hE8)) lut_n282 (.I0(n277), .I1(n280), .I2(n281), .O(n282));
  LUT3 #(.INIT(8'hE8)) lut_n283 (.I0(n266), .I1(n274), .I2(n282), .O(n283));
  LUT3 #(.INIT(8'hE8)) lut_n284 (.I0(x48), .I1(x49), .I2(x50), .O(n284));
  LUT5 #(.INIT(32'hE81717E8)) lut_n285 (.I0(x39), .I1(x40), .I2(x41), .I3(n278), .I4(n279), .O(n285));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n286 (.I0(x45), .I1(x46), .I2(x47), .I3(n284), .I4(n285), .O(n286));
  LUT3 #(.INIT(8'hE8)) lut_n287 (.I0(x54), .I1(x55), .I2(x56), .O(n287));
  LUT5 #(.INIT(32'hE81717E8)) lut_n288 (.I0(x45), .I1(x46), .I2(x47), .I3(n284), .I4(n285), .O(n288));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n289 (.I0(x51), .I1(x52), .I2(x53), .I3(n287), .I4(n288), .O(n289));
  LUT3 #(.INIT(8'h96)) lut_n290 (.I0(n277), .I1(n280), .I2(n281), .O(n290));
  LUT3 #(.INIT(8'hE8)) lut_n291 (.I0(n286), .I1(n289), .I2(n290), .O(n291));
  LUT3 #(.INIT(8'hE8)) lut_n292 (.I0(x60), .I1(x61), .I2(x62), .O(n292));
  LUT5 #(.INIT(32'hE81717E8)) lut_n293 (.I0(x51), .I1(x52), .I2(x53), .I3(n287), .I4(n288), .O(n293));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n294 (.I0(x57), .I1(x58), .I2(x59), .I3(n292), .I4(n293), .O(n294));
  LUT3 #(.INIT(8'hE8)) lut_n295 (.I0(x66), .I1(x67), .I2(x68), .O(n295));
  LUT5 #(.INIT(32'hE81717E8)) lut_n296 (.I0(x57), .I1(x58), .I2(x59), .I3(n292), .I4(n293), .O(n296));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n297 (.I0(x63), .I1(x64), .I2(x65), .I3(n295), .I4(n296), .O(n297));
  LUT3 #(.INIT(8'h96)) lut_n298 (.I0(n286), .I1(n289), .I2(n290), .O(n298));
  LUT3 #(.INIT(8'hE8)) lut_n299 (.I0(n294), .I1(n297), .I2(n298), .O(n299));
  LUT3 #(.INIT(8'h96)) lut_n300 (.I0(n266), .I1(n274), .I2(n282), .O(n300));
  LUT3 #(.INIT(8'hE8)) lut_n301 (.I0(n291), .I1(n299), .I2(n300), .O(n301));
  LUT3 #(.INIT(8'hE8)) lut_n302 (.I0(x72), .I1(x73), .I2(x74), .O(n302));
  LUT5 #(.INIT(32'hE81717E8)) lut_n303 (.I0(x63), .I1(x64), .I2(x65), .I3(n295), .I4(n296), .O(n303));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n304 (.I0(x69), .I1(x70), .I2(x71), .I3(n302), .I4(n303), .O(n304));
  LUT3 #(.INIT(8'hE8)) lut_n305 (.I0(x78), .I1(x79), .I2(x80), .O(n305));
  LUT5 #(.INIT(32'hE81717E8)) lut_n306 (.I0(x69), .I1(x70), .I2(x71), .I3(n302), .I4(n303), .O(n306));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n307 (.I0(x75), .I1(x76), .I2(x77), .I3(n305), .I4(n306), .O(n307));
  LUT3 #(.INIT(8'h96)) lut_n308 (.I0(n294), .I1(n297), .I2(n298), .O(n308));
  LUT3 #(.INIT(8'hE8)) lut_n309 (.I0(n304), .I1(n307), .I2(n308), .O(n309));
  LUT3 #(.INIT(8'hE8)) lut_n310 (.I0(x84), .I1(x85), .I2(x86), .O(n310));
  LUT5 #(.INIT(32'hE81717E8)) lut_n311 (.I0(x75), .I1(x76), .I2(x77), .I3(n305), .I4(n306), .O(n311));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n312 (.I0(x81), .I1(x82), .I2(x83), .I3(n310), .I4(n311), .O(n312));
  LUT3 #(.INIT(8'hE8)) lut_n313 (.I0(x90), .I1(x91), .I2(x92), .O(n313));
  LUT5 #(.INIT(32'hE81717E8)) lut_n314 (.I0(x81), .I1(x82), .I2(x83), .I3(n310), .I4(n311), .O(n314));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n315 (.I0(x87), .I1(x88), .I2(x89), .I3(n313), .I4(n314), .O(n315));
  LUT3 #(.INIT(8'h96)) lut_n316 (.I0(n304), .I1(n307), .I2(n308), .O(n316));
  LUT3 #(.INIT(8'hE8)) lut_n317 (.I0(n312), .I1(n315), .I2(n316), .O(n317));
  LUT3 #(.INIT(8'h96)) lut_n318 (.I0(n291), .I1(n299), .I2(n300), .O(n318));
  LUT3 #(.INIT(8'hE8)) lut_n319 (.I0(n309), .I1(n317), .I2(n318), .O(n319));
  LUT3 #(.INIT(8'hE8)) lut_n320 (.I0(n283), .I1(n301), .I2(n319), .O(n320));
  LUT3 #(.INIT(8'hE8)) lut_n321 (.I0(x96), .I1(x97), .I2(x98), .O(n321));
  LUT5 #(.INIT(32'hE81717E8)) lut_n322 (.I0(x87), .I1(x88), .I2(x89), .I3(n313), .I4(n314), .O(n322));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n323 (.I0(x93), .I1(x94), .I2(x95), .I3(n321), .I4(n322), .O(n323));
  LUT3 #(.INIT(8'hE8)) lut_n324 (.I0(x102), .I1(x103), .I2(x104), .O(n324));
  LUT5 #(.INIT(32'hE81717E8)) lut_n325 (.I0(x93), .I1(x94), .I2(x95), .I3(n321), .I4(n322), .O(n325));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n326 (.I0(x99), .I1(x100), .I2(x101), .I3(n324), .I4(n325), .O(n326));
  LUT3 #(.INIT(8'h96)) lut_n327 (.I0(n312), .I1(n315), .I2(n316), .O(n327));
  LUT3 #(.INIT(8'hE8)) lut_n328 (.I0(n323), .I1(n326), .I2(n327), .O(n328));
  LUT3 #(.INIT(8'hE8)) lut_n329 (.I0(x108), .I1(x109), .I2(x110), .O(n329));
  LUT5 #(.INIT(32'hE81717E8)) lut_n330 (.I0(x99), .I1(x100), .I2(x101), .I3(n324), .I4(n325), .O(n330));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n331 (.I0(x105), .I1(x106), .I2(x107), .I3(n329), .I4(n330), .O(n331));
  LUT3 #(.INIT(8'hE8)) lut_n332 (.I0(x114), .I1(x115), .I2(x116), .O(n332));
  LUT5 #(.INIT(32'hE81717E8)) lut_n333 (.I0(x105), .I1(x106), .I2(x107), .I3(n329), .I4(n330), .O(n333));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n334 (.I0(x111), .I1(x112), .I2(x113), .I3(n332), .I4(n333), .O(n334));
  LUT3 #(.INIT(8'h96)) lut_n335 (.I0(n323), .I1(n326), .I2(n327), .O(n335));
  LUT3 #(.INIT(8'hE8)) lut_n336 (.I0(n331), .I1(n334), .I2(n335), .O(n336));
  LUT3 #(.INIT(8'h96)) lut_n337 (.I0(n309), .I1(n317), .I2(n318), .O(n337));
  LUT3 #(.INIT(8'hE8)) lut_n338 (.I0(n328), .I1(n336), .I2(n337), .O(n338));
  LUT3 #(.INIT(8'hE8)) lut_n339 (.I0(x120), .I1(x121), .I2(x122), .O(n339));
  LUT5 #(.INIT(32'hE81717E8)) lut_n340 (.I0(x111), .I1(x112), .I2(x113), .I3(n332), .I4(n333), .O(n340));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n341 (.I0(x117), .I1(x118), .I2(x119), .I3(n339), .I4(n340), .O(n341));
  LUT3 #(.INIT(8'hE8)) lut_n342 (.I0(x126), .I1(x127), .I2(x128), .O(n342));
  LUT5 #(.INIT(32'hE81717E8)) lut_n343 (.I0(x117), .I1(x118), .I2(x119), .I3(n339), .I4(n340), .O(n343));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n344 (.I0(x123), .I1(x124), .I2(x125), .I3(n342), .I4(n343), .O(n344));
  LUT3 #(.INIT(8'h96)) lut_n345 (.I0(n331), .I1(n334), .I2(n335), .O(n345));
  LUT3 #(.INIT(8'hE8)) lut_n346 (.I0(n341), .I1(n344), .I2(n345), .O(n346));
  LUT3 #(.INIT(8'hE8)) lut_n347 (.I0(x132), .I1(x133), .I2(x134), .O(n347));
  LUT5 #(.INIT(32'hE81717E8)) lut_n348 (.I0(x123), .I1(x124), .I2(x125), .I3(n342), .I4(n343), .O(n348));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n349 (.I0(x129), .I1(x130), .I2(x131), .I3(n347), .I4(n348), .O(n349));
  LUT3 #(.INIT(8'hE8)) lut_n350 (.I0(x138), .I1(x139), .I2(x140), .O(n350));
  LUT5 #(.INIT(32'hE81717E8)) lut_n351 (.I0(x129), .I1(x130), .I2(x131), .I3(n347), .I4(n348), .O(n351));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n352 (.I0(x135), .I1(x136), .I2(x137), .I3(n350), .I4(n351), .O(n352));
  LUT3 #(.INIT(8'h96)) lut_n353 (.I0(n341), .I1(n344), .I2(n345), .O(n353));
  LUT3 #(.INIT(8'hE8)) lut_n354 (.I0(n349), .I1(n352), .I2(n353), .O(n354));
  LUT3 #(.INIT(8'h96)) lut_n355 (.I0(n328), .I1(n336), .I2(n337), .O(n355));
  LUT3 #(.INIT(8'hE8)) lut_n356 (.I0(n346), .I1(n354), .I2(n355), .O(n356));
  LUT3 #(.INIT(8'h96)) lut_n357 (.I0(n283), .I1(n301), .I2(n319), .O(n357));
  LUT3 #(.INIT(8'hE8)) lut_n358 (.I0(n338), .I1(n356), .I2(n357), .O(n358));
  LUT3 #(.INIT(8'hE8)) lut_n359 (.I0(x144), .I1(x145), .I2(x146), .O(n359));
  LUT5 #(.INIT(32'hE81717E8)) lut_n360 (.I0(x135), .I1(x136), .I2(x137), .I3(n350), .I4(n351), .O(n360));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n361 (.I0(x141), .I1(x142), .I2(x143), .I3(n359), .I4(n360), .O(n361));
  LUT3 #(.INIT(8'hE8)) lut_n362 (.I0(x150), .I1(x151), .I2(x152), .O(n362));
  LUT5 #(.INIT(32'hE81717E8)) lut_n363 (.I0(x141), .I1(x142), .I2(x143), .I3(n359), .I4(n360), .O(n363));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n364 (.I0(x147), .I1(x148), .I2(x149), .I3(n362), .I4(n363), .O(n364));
  LUT3 #(.INIT(8'h96)) lut_n365 (.I0(n349), .I1(n352), .I2(n353), .O(n365));
  LUT3 #(.INIT(8'hE8)) lut_n366 (.I0(n361), .I1(n364), .I2(n365), .O(n366));
  LUT3 #(.INIT(8'hE8)) lut_n367 (.I0(x156), .I1(x157), .I2(x158), .O(n367));
  LUT5 #(.INIT(32'hE81717E8)) lut_n368 (.I0(x147), .I1(x148), .I2(x149), .I3(n362), .I4(n363), .O(n368));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n369 (.I0(x153), .I1(x154), .I2(x155), .I3(n367), .I4(n368), .O(n369));
  LUT3 #(.INIT(8'hE8)) lut_n370 (.I0(x162), .I1(x163), .I2(x164), .O(n370));
  LUT5 #(.INIT(32'hE81717E8)) lut_n371 (.I0(x153), .I1(x154), .I2(x155), .I3(n367), .I4(n368), .O(n371));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n372 (.I0(x159), .I1(x160), .I2(x161), .I3(n370), .I4(n371), .O(n372));
  LUT3 #(.INIT(8'h96)) lut_n373 (.I0(n361), .I1(n364), .I2(n365), .O(n373));
  LUT3 #(.INIT(8'hE8)) lut_n374 (.I0(n369), .I1(n372), .I2(n373), .O(n374));
  LUT3 #(.INIT(8'h96)) lut_n375 (.I0(n346), .I1(n354), .I2(n355), .O(n375));
  LUT3 #(.INIT(8'hE8)) lut_n376 (.I0(n366), .I1(n374), .I2(n375), .O(n376));
  LUT3 #(.INIT(8'hE8)) lut_n377 (.I0(x168), .I1(x169), .I2(x170), .O(n377));
  LUT5 #(.INIT(32'hE81717E8)) lut_n378 (.I0(x159), .I1(x160), .I2(x161), .I3(n370), .I4(n371), .O(n378));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n379 (.I0(x165), .I1(x166), .I2(x167), .I3(n377), .I4(n378), .O(n379));
  LUT3 #(.INIT(8'hE8)) lut_n380 (.I0(x174), .I1(x175), .I2(x176), .O(n380));
  LUT5 #(.INIT(32'hE81717E8)) lut_n381 (.I0(x165), .I1(x166), .I2(x167), .I3(n377), .I4(n378), .O(n381));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n382 (.I0(x171), .I1(x172), .I2(x173), .I3(n380), .I4(n381), .O(n382));
  LUT3 #(.INIT(8'h96)) lut_n383 (.I0(n369), .I1(n372), .I2(n373), .O(n383));
  LUT3 #(.INIT(8'hE8)) lut_n384 (.I0(n379), .I1(n382), .I2(n383), .O(n384));
  LUT3 #(.INIT(8'hE8)) lut_n385 (.I0(x180), .I1(x181), .I2(x182), .O(n385));
  LUT5 #(.INIT(32'hE81717E8)) lut_n386 (.I0(x171), .I1(x172), .I2(x173), .I3(n380), .I4(n381), .O(n386));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n387 (.I0(x177), .I1(x178), .I2(x179), .I3(n385), .I4(n386), .O(n387));
  LUT3 #(.INIT(8'hE8)) lut_n388 (.I0(x186), .I1(x187), .I2(x188), .O(n388));
  LUT5 #(.INIT(32'hE81717E8)) lut_n389 (.I0(x177), .I1(x178), .I2(x179), .I3(n385), .I4(n386), .O(n389));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n390 (.I0(x183), .I1(x184), .I2(x185), .I3(n388), .I4(n389), .O(n390));
  LUT3 #(.INIT(8'h96)) lut_n391 (.I0(n379), .I1(n382), .I2(n383), .O(n391));
  LUT3 #(.INIT(8'hE8)) lut_n392 (.I0(n387), .I1(n390), .I2(n391), .O(n392));
  LUT3 #(.INIT(8'h96)) lut_n393 (.I0(n366), .I1(n374), .I2(n375), .O(n393));
  LUT3 #(.INIT(8'hE8)) lut_n394 (.I0(n384), .I1(n392), .I2(n393), .O(n394));
  LUT3 #(.INIT(8'h96)) lut_n395 (.I0(n338), .I1(n356), .I2(n357), .O(n395));
  LUT3 #(.INIT(8'hE8)) lut_n396 (.I0(n376), .I1(n394), .I2(n395), .O(n396));
  LUT3 #(.INIT(8'hE8)) lut_n397 (.I0(n320), .I1(n358), .I2(n396), .O(n397));
  LUT3 #(.INIT(8'hE8)) lut_n398 (.I0(x192), .I1(x193), .I2(x194), .O(n398));
  LUT5 #(.INIT(32'hE81717E8)) lut_n399 (.I0(x183), .I1(x184), .I2(x185), .I3(n388), .I4(n389), .O(n399));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n400 (.I0(x189), .I1(x190), .I2(x191), .I3(n398), .I4(n399), .O(n400));
  LUT3 #(.INIT(8'hE8)) lut_n401 (.I0(x198), .I1(x199), .I2(x200), .O(n401));
  LUT5 #(.INIT(32'hE81717E8)) lut_n402 (.I0(x189), .I1(x190), .I2(x191), .I3(n398), .I4(n399), .O(n402));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n403 (.I0(x195), .I1(x196), .I2(x197), .I3(n401), .I4(n402), .O(n403));
  LUT3 #(.INIT(8'h96)) lut_n404 (.I0(n387), .I1(n390), .I2(n391), .O(n404));
  LUT3 #(.INIT(8'hE8)) lut_n405 (.I0(n400), .I1(n403), .I2(n404), .O(n405));
  LUT3 #(.INIT(8'hE8)) lut_n406 (.I0(x204), .I1(x205), .I2(x206), .O(n406));
  LUT5 #(.INIT(32'hE81717E8)) lut_n407 (.I0(x195), .I1(x196), .I2(x197), .I3(n401), .I4(n402), .O(n407));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n408 (.I0(x201), .I1(x202), .I2(x203), .I3(n406), .I4(n407), .O(n408));
  LUT3 #(.INIT(8'hE8)) lut_n409 (.I0(x210), .I1(x211), .I2(x212), .O(n409));
  LUT5 #(.INIT(32'hE81717E8)) lut_n410 (.I0(x201), .I1(x202), .I2(x203), .I3(n406), .I4(n407), .O(n410));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n411 (.I0(x207), .I1(x208), .I2(x209), .I3(n409), .I4(n410), .O(n411));
  LUT3 #(.INIT(8'h96)) lut_n412 (.I0(n400), .I1(n403), .I2(n404), .O(n412));
  LUT3 #(.INIT(8'hE8)) lut_n413 (.I0(n408), .I1(n411), .I2(n412), .O(n413));
  LUT3 #(.INIT(8'h96)) lut_n414 (.I0(n384), .I1(n392), .I2(n393), .O(n414));
  LUT3 #(.INIT(8'hE8)) lut_n415 (.I0(n405), .I1(n413), .I2(n414), .O(n415));
  LUT3 #(.INIT(8'hE8)) lut_n416 (.I0(x216), .I1(x217), .I2(x218), .O(n416));
  LUT5 #(.INIT(32'hE81717E8)) lut_n417 (.I0(x207), .I1(x208), .I2(x209), .I3(n409), .I4(n410), .O(n417));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n418 (.I0(x213), .I1(x214), .I2(x215), .I3(n416), .I4(n417), .O(n418));
  LUT3 #(.INIT(8'hE8)) lut_n419 (.I0(x222), .I1(x223), .I2(x224), .O(n419));
  LUT5 #(.INIT(32'hE81717E8)) lut_n420 (.I0(x213), .I1(x214), .I2(x215), .I3(n416), .I4(n417), .O(n420));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n421 (.I0(x219), .I1(x220), .I2(x221), .I3(n419), .I4(n420), .O(n421));
  LUT3 #(.INIT(8'h96)) lut_n422 (.I0(n408), .I1(n411), .I2(n412), .O(n422));
  LUT3 #(.INIT(8'hE8)) lut_n423 (.I0(n418), .I1(n421), .I2(n422), .O(n423));
  LUT3 #(.INIT(8'hE8)) lut_n424 (.I0(x228), .I1(x229), .I2(x230), .O(n424));
  LUT5 #(.INIT(32'hE81717E8)) lut_n425 (.I0(x219), .I1(x220), .I2(x221), .I3(n419), .I4(n420), .O(n425));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n426 (.I0(x225), .I1(x226), .I2(x227), .I3(n424), .I4(n425), .O(n426));
  LUT3 #(.INIT(8'hE8)) lut_n427 (.I0(x234), .I1(x235), .I2(x236), .O(n427));
  LUT5 #(.INIT(32'hE81717E8)) lut_n428 (.I0(x225), .I1(x226), .I2(x227), .I3(n424), .I4(n425), .O(n428));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n429 (.I0(x231), .I1(x232), .I2(x233), .I3(n427), .I4(n428), .O(n429));
  LUT3 #(.INIT(8'h96)) lut_n430 (.I0(n418), .I1(n421), .I2(n422), .O(n430));
  LUT3 #(.INIT(8'hE8)) lut_n431 (.I0(n426), .I1(n429), .I2(n430), .O(n431));
  LUT3 #(.INIT(8'h96)) lut_n432 (.I0(n405), .I1(n413), .I2(n414), .O(n432));
  LUT3 #(.INIT(8'hE8)) lut_n433 (.I0(n423), .I1(n431), .I2(n432), .O(n433));
  LUT3 #(.INIT(8'h96)) lut_n434 (.I0(n376), .I1(n394), .I2(n395), .O(n434));
  LUT3 #(.INIT(8'hE8)) lut_n435 (.I0(n415), .I1(n433), .I2(n434), .O(n435));
  LUT3 #(.INIT(8'hE8)) lut_n436 (.I0(x240), .I1(x241), .I2(x242), .O(n436));
  LUT5 #(.INIT(32'hE81717E8)) lut_n437 (.I0(x231), .I1(x232), .I2(x233), .I3(n427), .I4(n428), .O(n437));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n438 (.I0(x237), .I1(x238), .I2(x239), .I3(n436), .I4(n437), .O(n438));
  LUT3 #(.INIT(8'hE8)) lut_n439 (.I0(x246), .I1(x247), .I2(x248), .O(n439));
  LUT5 #(.INIT(32'hE81717E8)) lut_n440 (.I0(x237), .I1(x238), .I2(x239), .I3(n436), .I4(n437), .O(n440));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n441 (.I0(x243), .I1(x244), .I2(x245), .I3(n439), .I4(n440), .O(n441));
  LUT3 #(.INIT(8'h96)) lut_n442 (.I0(n426), .I1(n429), .I2(n430), .O(n442));
  LUT3 #(.INIT(8'hE8)) lut_n443 (.I0(n438), .I1(n441), .I2(n442), .O(n443));
  LUT3 #(.INIT(8'hE8)) lut_n444 (.I0(x252), .I1(x253), .I2(x254), .O(n444));
  LUT5 #(.INIT(32'hE81717E8)) lut_n445 (.I0(x243), .I1(x244), .I2(x245), .I3(n439), .I4(n440), .O(n445));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n446 (.I0(x249), .I1(x250), .I2(x251), .I3(n444), .I4(n445), .O(n446));
  LUT3 #(.INIT(8'h96)) lut_n447 (.I0(x0), .I1(x1), .I2(x2), .O(n447));
  LUT3 #(.INIT(8'h96)) lut_n448 (.I0(x6), .I1(x7), .I2(x8), .O(n448));
  LUT5 #(.INIT(32'hFF969600)) lut_n449 (.I0(x3), .I1(x4), .I2(x5), .I3(n447), .I4(n448), .O(n449));
  LUT3 #(.INIT(8'h96)) lut_n450 (.I0(x12), .I1(x13), .I2(x14), .O(n450));
  LUT5 #(.INIT(32'h96696996)) lut_n451 (.I0(x3), .I1(x4), .I2(x5), .I3(n447), .I4(n448), .O(n451));
  LUT5 #(.INIT(32'hFF969600)) lut_n452 (.I0(x9), .I1(x10), .I2(x11), .I3(n450), .I4(n451), .O(n452));
  LUT5 #(.INIT(32'hE81717E8)) lut_n453 (.I0(x249), .I1(x250), .I2(x251), .I3(n444), .I4(n445), .O(n453));
  LUT3 #(.INIT(8'hE8)) lut_n454 (.I0(n449), .I1(n452), .I2(n453), .O(n454));
  LUT3 #(.INIT(8'h96)) lut_n455 (.I0(n438), .I1(n441), .I2(n442), .O(n455));
  LUT3 #(.INIT(8'hE8)) lut_n456 (.I0(n446), .I1(n454), .I2(n455), .O(n456));
  LUT3 #(.INIT(8'h96)) lut_n457 (.I0(n423), .I1(n431), .I2(n432), .O(n457));
  LUT3 #(.INIT(8'hE8)) lut_n458 (.I0(n443), .I1(n456), .I2(n457), .O(n458));
  LUT3 #(.INIT(8'h96)) lut_n459 (.I0(x18), .I1(x19), .I2(x20), .O(n459));
  LUT5 #(.INIT(32'h96696996)) lut_n460 (.I0(x9), .I1(x10), .I2(x11), .I3(n450), .I4(n451), .O(n460));
  LUT5 #(.INIT(32'hFF969600)) lut_n461 (.I0(x15), .I1(x16), .I2(x17), .I3(n459), .I4(n460), .O(n461));
  LUT3 #(.INIT(8'h96)) lut_n462 (.I0(x24), .I1(x25), .I2(x26), .O(n462));
  LUT5 #(.INIT(32'h96696996)) lut_n463 (.I0(x15), .I1(x16), .I2(x17), .I3(n459), .I4(n460), .O(n463));
  LUT5 #(.INIT(32'hFF969600)) lut_n464 (.I0(x21), .I1(x22), .I2(x23), .I3(n462), .I4(n463), .O(n464));
  LUT3 #(.INIT(8'h96)) lut_n465 (.I0(n449), .I1(n452), .I2(n453), .O(n465));
  LUT3 #(.INIT(8'hE8)) lut_n466 (.I0(n461), .I1(n464), .I2(n465), .O(n466));
  LUT3 #(.INIT(8'h96)) lut_n467 (.I0(x27), .I1(x28), .I2(x29), .O(n467));
  LUT5 #(.INIT(32'h96696996)) lut_n468 (.I0(x21), .I1(x22), .I2(x23), .I3(n462), .I4(n463), .O(n468));
  LUT5 #(.INIT(32'hFF969600)) lut_n469 (.I0(x30), .I1(x31), .I2(x32), .I3(n467), .I4(n468), .O(n469));
  LUT3 #(.INIT(8'h96)) lut_n470 (.I0(x36), .I1(x37), .I2(x38), .O(n470));
  LUT5 #(.INIT(32'h96696996)) lut_n471 (.I0(x30), .I1(x31), .I2(x32), .I3(n467), .I4(n468), .O(n471));
  LUT5 #(.INIT(32'hFF969600)) lut_n472 (.I0(x33), .I1(x34), .I2(x35), .I3(n470), .I4(n471), .O(n472));
  LUT3 #(.INIT(8'h96)) lut_n473 (.I0(n461), .I1(n464), .I2(n465), .O(n473));
  LUT3 #(.INIT(8'hE8)) lut_n474 (.I0(n469), .I1(n472), .I2(n473), .O(n474));
  LUT3 #(.INIT(8'h96)) lut_n475 (.I0(n446), .I1(n454), .I2(n455), .O(n475));
  LUT3 #(.INIT(8'hE8)) lut_n476 (.I0(n466), .I1(n474), .I2(n475), .O(n476));
  LUT3 #(.INIT(8'h96)) lut_n477 (.I0(x42), .I1(x43), .I2(x44), .O(n477));
  LUT5 #(.INIT(32'h96696996)) lut_n478 (.I0(x33), .I1(x34), .I2(x35), .I3(n470), .I4(n471), .O(n478));
  LUT5 #(.INIT(32'hFF969600)) lut_n479 (.I0(x39), .I1(x40), .I2(x41), .I3(n477), .I4(n478), .O(n479));
  LUT3 #(.INIT(8'h96)) lut_n480 (.I0(x48), .I1(x49), .I2(x50), .O(n480));
  LUT5 #(.INIT(32'h96696996)) lut_n481 (.I0(x39), .I1(x40), .I2(x41), .I3(n477), .I4(n478), .O(n481));
  LUT5 #(.INIT(32'hFF969600)) lut_n482 (.I0(x45), .I1(x46), .I2(x47), .I3(n480), .I4(n481), .O(n482));
  LUT3 #(.INIT(8'h96)) lut_n483 (.I0(n469), .I1(n472), .I2(n473), .O(n483));
  LUT3 #(.INIT(8'hE8)) lut_n484 (.I0(n479), .I1(n482), .I2(n483), .O(n484));
  LUT3 #(.INIT(8'h96)) lut_n485 (.I0(x54), .I1(x55), .I2(x56), .O(n485));
  LUT5 #(.INIT(32'h96696996)) lut_n486 (.I0(x45), .I1(x46), .I2(x47), .I3(n480), .I4(n481), .O(n486));
  LUT5 #(.INIT(32'hFF969600)) lut_n487 (.I0(x51), .I1(x52), .I2(x53), .I3(n485), .I4(n486), .O(n487));
  LUT3 #(.INIT(8'h96)) lut_n488 (.I0(x60), .I1(x61), .I2(x62), .O(n488));
  LUT5 #(.INIT(32'h96696996)) lut_n489 (.I0(x51), .I1(x52), .I2(x53), .I3(n485), .I4(n486), .O(n489));
  LUT5 #(.INIT(32'hFF969600)) lut_n490 (.I0(x57), .I1(x58), .I2(x59), .I3(n488), .I4(n489), .O(n490));
  LUT3 #(.INIT(8'h96)) lut_n491 (.I0(n479), .I1(n482), .I2(n483), .O(n491));
  LUT3 #(.INIT(8'hE8)) lut_n492 (.I0(n487), .I1(n490), .I2(n491), .O(n492));
  LUT3 #(.INIT(8'h96)) lut_n493 (.I0(n466), .I1(n474), .I2(n475), .O(n493));
  LUT3 #(.INIT(8'hE8)) lut_n494 (.I0(n484), .I1(n492), .I2(n493), .O(n494));
  LUT3 #(.INIT(8'h96)) lut_n495 (.I0(n443), .I1(n456), .I2(n457), .O(n495));
  LUT3 #(.INIT(8'hE8)) lut_n496 (.I0(n476), .I1(n494), .I2(n495), .O(n496));
  LUT3 #(.INIT(8'h96)) lut_n497 (.I0(n415), .I1(n433), .I2(n434), .O(n497));
  LUT3 #(.INIT(8'hE8)) lut_n498 (.I0(n458), .I1(n496), .I2(n497), .O(n498));
  LUT3 #(.INIT(8'h96)) lut_n499 (.I0(n320), .I1(n358), .I2(n396), .O(n499));
  LUT3 #(.INIT(8'h96)) lut_n500 (.I0(x66), .I1(x67), .I2(x68), .O(n500));
  LUT5 #(.INIT(32'h96696996)) lut_n501 (.I0(x57), .I1(x58), .I2(x59), .I3(n488), .I4(n489), .O(n501));
  LUT5 #(.INIT(32'hFF969600)) lut_n502 (.I0(x63), .I1(x64), .I2(x65), .I3(n500), .I4(n501), .O(n502));
  LUT3 #(.INIT(8'h96)) lut_n503 (.I0(x72), .I1(x73), .I2(x74), .O(n503));
  LUT5 #(.INIT(32'h96696996)) lut_n504 (.I0(x63), .I1(x64), .I2(x65), .I3(n500), .I4(n501), .O(n504));
  LUT5 #(.INIT(32'hFF969600)) lut_n505 (.I0(x69), .I1(x70), .I2(x71), .I3(n503), .I4(n504), .O(n505));
  LUT3 #(.INIT(8'h96)) lut_n506 (.I0(n487), .I1(n490), .I2(n491), .O(n506));
  LUT3 #(.INIT(8'hE8)) lut_n507 (.I0(n502), .I1(n505), .I2(n506), .O(n507));
  LUT3 #(.INIT(8'h96)) lut_n508 (.I0(x78), .I1(x79), .I2(x80), .O(n508));
  LUT5 #(.INIT(32'h96696996)) lut_n509 (.I0(x69), .I1(x70), .I2(x71), .I3(n503), .I4(n504), .O(n509));
  LUT5 #(.INIT(32'hFF969600)) lut_n510 (.I0(x75), .I1(x76), .I2(x77), .I3(n508), .I4(n509), .O(n510));
  LUT3 #(.INIT(8'h96)) lut_n511 (.I0(x84), .I1(x85), .I2(x86), .O(n511));
  LUT5 #(.INIT(32'h96696996)) lut_n512 (.I0(x75), .I1(x76), .I2(x77), .I3(n508), .I4(n509), .O(n512));
  LUT5 #(.INIT(32'hFF969600)) lut_n513 (.I0(x81), .I1(x82), .I2(x83), .I3(n511), .I4(n512), .O(n513));
  LUT3 #(.INIT(8'h96)) lut_n514 (.I0(n502), .I1(n505), .I2(n506), .O(n514));
  LUT3 #(.INIT(8'hE8)) lut_n515 (.I0(n510), .I1(n513), .I2(n514), .O(n515));
  LUT3 #(.INIT(8'h96)) lut_n516 (.I0(n484), .I1(n492), .I2(n493), .O(n516));
  LUT3 #(.INIT(8'hE8)) lut_n517 (.I0(n507), .I1(n515), .I2(n516), .O(n517));
  LUT3 #(.INIT(8'h96)) lut_n518 (.I0(x90), .I1(x91), .I2(x92), .O(n518));
  LUT5 #(.INIT(32'h96696996)) lut_n519 (.I0(x81), .I1(x82), .I2(x83), .I3(n511), .I4(n512), .O(n519));
  LUT5 #(.INIT(32'hFF969600)) lut_n520 (.I0(x87), .I1(x88), .I2(x89), .I3(n518), .I4(n519), .O(n520));
  LUT3 #(.INIT(8'h96)) lut_n521 (.I0(x96), .I1(x97), .I2(x98), .O(n521));
  LUT5 #(.INIT(32'h96696996)) lut_n522 (.I0(x87), .I1(x88), .I2(x89), .I3(n518), .I4(n519), .O(n522));
  LUT5 #(.INIT(32'hFF969600)) lut_n523 (.I0(x93), .I1(x94), .I2(x95), .I3(n521), .I4(n522), .O(n523));
  LUT3 #(.INIT(8'h96)) lut_n524 (.I0(n510), .I1(n513), .I2(n514), .O(n524));
  LUT3 #(.INIT(8'hE8)) lut_n525 (.I0(n520), .I1(n523), .I2(n524), .O(n525));
  LUT3 #(.INIT(8'h96)) lut_n526 (.I0(x102), .I1(x103), .I2(x104), .O(n526));
  LUT5 #(.INIT(32'h96696996)) lut_n527 (.I0(x93), .I1(x94), .I2(x95), .I3(n521), .I4(n522), .O(n527));
  LUT5 #(.INIT(32'hFF969600)) lut_n528 (.I0(x99), .I1(x100), .I2(x101), .I3(n526), .I4(n527), .O(n528));
  LUT3 #(.INIT(8'h96)) lut_n529 (.I0(x108), .I1(x109), .I2(x110), .O(n529));
  LUT5 #(.INIT(32'h96696996)) lut_n530 (.I0(x99), .I1(x100), .I2(x101), .I3(n526), .I4(n527), .O(n530));
  LUT5 #(.INIT(32'hFF969600)) lut_n531 (.I0(x105), .I1(x106), .I2(x107), .I3(n529), .I4(n530), .O(n531));
  LUT3 #(.INIT(8'h96)) lut_n532 (.I0(n520), .I1(n523), .I2(n524), .O(n532));
  LUT3 #(.INIT(8'hE8)) lut_n533 (.I0(n528), .I1(n531), .I2(n532), .O(n533));
  LUT3 #(.INIT(8'h96)) lut_n534 (.I0(n507), .I1(n515), .I2(n516), .O(n534));
  LUT3 #(.INIT(8'hE8)) lut_n535 (.I0(n525), .I1(n533), .I2(n534), .O(n535));
  LUT3 #(.INIT(8'h96)) lut_n536 (.I0(n476), .I1(n494), .I2(n495), .O(n536));
  LUT3 #(.INIT(8'hE8)) lut_n537 (.I0(n517), .I1(n535), .I2(n536), .O(n537));
  LUT3 #(.INIT(8'h96)) lut_n538 (.I0(x114), .I1(x115), .I2(x116), .O(n538));
  LUT5 #(.INIT(32'h96696996)) lut_n539 (.I0(x105), .I1(x106), .I2(x107), .I3(n529), .I4(n530), .O(n539));
  LUT5 #(.INIT(32'hFF969600)) lut_n540 (.I0(x111), .I1(x112), .I2(x113), .I3(n538), .I4(n539), .O(n540));
  LUT3 #(.INIT(8'h96)) lut_n541 (.I0(x120), .I1(x121), .I2(x122), .O(n541));
  LUT5 #(.INIT(32'h96696996)) lut_n542 (.I0(x111), .I1(x112), .I2(x113), .I3(n538), .I4(n539), .O(n542));
  LUT5 #(.INIT(32'hFF969600)) lut_n543 (.I0(x117), .I1(x118), .I2(x119), .I3(n541), .I4(n542), .O(n543));
  LUT3 #(.INIT(8'h96)) lut_n544 (.I0(n528), .I1(n531), .I2(n532), .O(n544));
  LUT3 #(.INIT(8'hE8)) lut_n545 (.I0(n540), .I1(n543), .I2(n544), .O(n545));
  LUT3 #(.INIT(8'h96)) lut_n546 (.I0(x126), .I1(x127), .I2(x128), .O(n546));
  LUT5 #(.INIT(32'h96696996)) lut_n547 (.I0(x117), .I1(x118), .I2(x119), .I3(n541), .I4(n542), .O(n547));
  LUT5 #(.INIT(32'hFF969600)) lut_n548 (.I0(x123), .I1(x124), .I2(x125), .I3(n546), .I4(n547), .O(n548));
  LUT3 #(.INIT(8'h96)) lut_n549 (.I0(x132), .I1(x133), .I2(x134), .O(n549));
  LUT5 #(.INIT(32'h96696996)) lut_n550 (.I0(x123), .I1(x124), .I2(x125), .I3(n546), .I4(n547), .O(n550));
  LUT5 #(.INIT(32'hFF969600)) lut_n551 (.I0(x129), .I1(x130), .I2(x131), .I3(n549), .I4(n550), .O(n551));
  LUT3 #(.INIT(8'h96)) lut_n552 (.I0(n540), .I1(n543), .I2(n544), .O(n552));
  LUT3 #(.INIT(8'hE8)) lut_n553 (.I0(n548), .I1(n551), .I2(n552), .O(n553));
  LUT3 #(.INIT(8'h96)) lut_n554 (.I0(n525), .I1(n533), .I2(n534), .O(n554));
  LUT3 #(.INIT(8'hE8)) lut_n555 (.I0(n545), .I1(n553), .I2(n554), .O(n555));
  LUT3 #(.INIT(8'h96)) lut_n556 (.I0(x138), .I1(x139), .I2(x140), .O(n556));
  LUT5 #(.INIT(32'h96696996)) lut_n557 (.I0(x129), .I1(x130), .I2(x131), .I3(n549), .I4(n550), .O(n557));
  LUT5 #(.INIT(32'hFF969600)) lut_n558 (.I0(x135), .I1(x136), .I2(x137), .I3(n556), .I4(n557), .O(n558));
  LUT3 #(.INIT(8'h96)) lut_n559 (.I0(x144), .I1(x145), .I2(x146), .O(n559));
  LUT5 #(.INIT(32'h96696996)) lut_n560 (.I0(x135), .I1(x136), .I2(x137), .I3(n556), .I4(n557), .O(n560));
  LUT5 #(.INIT(32'hFF969600)) lut_n561 (.I0(x141), .I1(x142), .I2(x143), .I3(n559), .I4(n560), .O(n561));
  LUT3 #(.INIT(8'h96)) lut_n562 (.I0(n548), .I1(n551), .I2(n552), .O(n562));
  LUT3 #(.INIT(8'hE8)) lut_n563 (.I0(n558), .I1(n561), .I2(n562), .O(n563));
  LUT3 #(.INIT(8'h96)) lut_n564 (.I0(x150), .I1(x151), .I2(x152), .O(n564));
  LUT5 #(.INIT(32'h96696996)) lut_n565 (.I0(x141), .I1(x142), .I2(x143), .I3(n559), .I4(n560), .O(n565));
  LUT5 #(.INIT(32'hFF969600)) lut_n566 (.I0(x147), .I1(x148), .I2(x149), .I3(n564), .I4(n565), .O(n566));
  LUT3 #(.INIT(8'h96)) lut_n567 (.I0(x156), .I1(x157), .I2(x158), .O(n567));
  LUT5 #(.INIT(32'h96696996)) lut_n568 (.I0(x147), .I1(x148), .I2(x149), .I3(n564), .I4(n565), .O(n568));
  LUT5 #(.INIT(32'hFF969600)) lut_n569 (.I0(x153), .I1(x154), .I2(x155), .I3(n567), .I4(n568), .O(n569));
  LUT3 #(.INIT(8'h96)) lut_n570 (.I0(n558), .I1(n561), .I2(n562), .O(n570));
  LUT3 #(.INIT(8'hE8)) lut_n571 (.I0(n566), .I1(n569), .I2(n570), .O(n571));
  LUT3 #(.INIT(8'h96)) lut_n572 (.I0(n545), .I1(n553), .I2(n554), .O(n572));
  LUT3 #(.INIT(8'hE8)) lut_n573 (.I0(n563), .I1(n571), .I2(n572), .O(n573));
  LUT3 #(.INIT(8'h96)) lut_n574 (.I0(n517), .I1(n535), .I2(n536), .O(n574));
  LUT3 #(.INIT(8'hE8)) lut_n575 (.I0(n555), .I1(n573), .I2(n574), .O(n575));
  LUT3 #(.INIT(8'h96)) lut_n576 (.I0(n458), .I1(n496), .I2(n497), .O(n576));
  LUT3 #(.INIT(8'hE8)) lut_n577 (.I0(n537), .I1(n575), .I2(n576), .O(n577));
  LUT3 #(.INIT(8'h96)) lut_n578 (.I0(x162), .I1(x163), .I2(x164), .O(n578));
  LUT5 #(.INIT(32'h96696996)) lut_n579 (.I0(x153), .I1(x154), .I2(x155), .I3(n567), .I4(n568), .O(n579));
  LUT5 #(.INIT(32'hFF969600)) lut_n580 (.I0(x159), .I1(x160), .I2(x161), .I3(n578), .I4(n579), .O(n580));
  LUT3 #(.INIT(8'h96)) lut_n581 (.I0(x168), .I1(x169), .I2(x170), .O(n581));
  LUT5 #(.INIT(32'h96696996)) lut_n582 (.I0(x159), .I1(x160), .I2(x161), .I3(n578), .I4(n579), .O(n582));
  LUT5 #(.INIT(32'hFF969600)) lut_n583 (.I0(x165), .I1(x166), .I2(x167), .I3(n581), .I4(n582), .O(n583));
  LUT3 #(.INIT(8'h96)) lut_n584 (.I0(n566), .I1(n569), .I2(n570), .O(n584));
  LUT3 #(.INIT(8'hE8)) lut_n585 (.I0(n580), .I1(n583), .I2(n584), .O(n585));
  LUT3 #(.INIT(8'h96)) lut_n586 (.I0(x174), .I1(x175), .I2(x176), .O(n586));
  LUT5 #(.INIT(32'h96696996)) lut_n587 (.I0(x165), .I1(x166), .I2(x167), .I3(n581), .I4(n582), .O(n587));
  LUT5 #(.INIT(32'hFF969600)) lut_n588 (.I0(x171), .I1(x172), .I2(x173), .I3(n586), .I4(n587), .O(n588));
  LUT3 #(.INIT(8'h96)) lut_n589 (.I0(x180), .I1(x181), .I2(x182), .O(n589));
  LUT5 #(.INIT(32'h96696996)) lut_n590 (.I0(x171), .I1(x172), .I2(x173), .I3(n586), .I4(n587), .O(n590));
  LUT5 #(.INIT(32'hFF969600)) lut_n591 (.I0(x177), .I1(x178), .I2(x179), .I3(n589), .I4(n590), .O(n591));
  LUT3 #(.INIT(8'h96)) lut_n592 (.I0(n580), .I1(n583), .I2(n584), .O(n592));
  LUT3 #(.INIT(8'hE8)) lut_n593 (.I0(n588), .I1(n591), .I2(n592), .O(n593));
  LUT3 #(.INIT(8'h96)) lut_n594 (.I0(n563), .I1(n571), .I2(n572), .O(n594));
  LUT3 #(.INIT(8'hE8)) lut_n595 (.I0(n585), .I1(n593), .I2(n594), .O(n595));
  LUT3 #(.INIT(8'h96)) lut_n596 (.I0(x186), .I1(x187), .I2(x188), .O(n596));
  LUT5 #(.INIT(32'h96696996)) lut_n597 (.I0(x177), .I1(x178), .I2(x179), .I3(n589), .I4(n590), .O(n597));
  LUT5 #(.INIT(32'hFF969600)) lut_n598 (.I0(x183), .I1(x184), .I2(x185), .I3(n596), .I4(n597), .O(n598));
  LUT3 #(.INIT(8'h96)) lut_n599 (.I0(x192), .I1(x193), .I2(x194), .O(n599));
  LUT5 #(.INIT(32'h96696996)) lut_n600 (.I0(x183), .I1(x184), .I2(x185), .I3(n596), .I4(n597), .O(n600));
  LUT5 #(.INIT(32'hFF969600)) lut_n601 (.I0(x189), .I1(x190), .I2(x191), .I3(n599), .I4(n600), .O(n601));
  LUT3 #(.INIT(8'h96)) lut_n602 (.I0(n588), .I1(n591), .I2(n592), .O(n602));
  LUT3 #(.INIT(8'hE8)) lut_n603 (.I0(n598), .I1(n601), .I2(n602), .O(n603));
  LUT3 #(.INIT(8'h96)) lut_n604 (.I0(x198), .I1(x199), .I2(x200), .O(n604));
  LUT5 #(.INIT(32'h96696996)) lut_n605 (.I0(x189), .I1(x190), .I2(x191), .I3(n599), .I4(n600), .O(n605));
  LUT5 #(.INIT(32'hFF969600)) lut_n606 (.I0(x195), .I1(x196), .I2(x197), .I3(n604), .I4(n605), .O(n606));
  LUT3 #(.INIT(8'h96)) lut_n607 (.I0(x204), .I1(x205), .I2(x206), .O(n607));
  LUT5 #(.INIT(32'h96696996)) lut_n608 (.I0(x195), .I1(x196), .I2(x197), .I3(n604), .I4(n605), .O(n608));
  LUT5 #(.INIT(32'hFF969600)) lut_n609 (.I0(x201), .I1(x202), .I2(x203), .I3(n607), .I4(n608), .O(n609));
  LUT3 #(.INIT(8'h96)) lut_n610 (.I0(n598), .I1(n601), .I2(n602), .O(n610));
  LUT3 #(.INIT(8'hE8)) lut_n611 (.I0(n606), .I1(n609), .I2(n610), .O(n611));
  LUT3 #(.INIT(8'h96)) lut_n612 (.I0(n585), .I1(n593), .I2(n594), .O(n612));
  LUT3 #(.INIT(8'hE8)) lut_n613 (.I0(n603), .I1(n611), .I2(n612), .O(n613));
  LUT3 #(.INIT(8'h96)) lut_n614 (.I0(n555), .I1(n573), .I2(n574), .O(n614));
  LUT3 #(.INIT(8'h96)) lut_n615 (.I0(x210), .I1(x211), .I2(x212), .O(n615));
  LUT5 #(.INIT(32'h96696996)) lut_n616 (.I0(x201), .I1(x202), .I2(x203), .I3(n607), .I4(n608), .O(n616));
  LUT5 #(.INIT(32'hFF969600)) lut_n617 (.I0(x207), .I1(x208), .I2(x209), .I3(n615), .I4(n616), .O(n617));
  LUT3 #(.INIT(8'h96)) lut_n618 (.I0(x216), .I1(x217), .I2(x218), .O(n618));
  LUT5 #(.INIT(32'h96696996)) lut_n619 (.I0(x207), .I1(x208), .I2(x209), .I3(n615), .I4(n616), .O(n619));
  LUT5 #(.INIT(32'hFF969600)) lut_n620 (.I0(x213), .I1(x214), .I2(x215), .I3(n618), .I4(n619), .O(n620));
  LUT3 #(.INIT(8'h96)) lut_n621 (.I0(n606), .I1(n609), .I2(n610), .O(n621));
  LUT3 #(.INIT(8'hE8)) lut_n622 (.I0(n617), .I1(n620), .I2(n621), .O(n622));
  LUT3 #(.INIT(8'h96)) lut_n623 (.I0(x222), .I1(x223), .I2(x224), .O(n623));
  LUT5 #(.INIT(32'h96696996)) lut_n624 (.I0(x213), .I1(x214), .I2(x215), .I3(n618), .I4(n619), .O(n624));
  LUT5 #(.INIT(32'hFF969600)) lut_n625 (.I0(x219), .I1(x220), .I2(x221), .I3(n623), .I4(n624), .O(n625));
  LUT3 #(.INIT(8'h96)) lut_n626 (.I0(x228), .I1(x229), .I2(x230), .O(n626));
  LUT5 #(.INIT(32'h96696996)) lut_n627 (.I0(x219), .I1(x220), .I2(x221), .I3(n623), .I4(n624), .O(n627));
  LUT5 #(.INIT(32'hFF969600)) lut_n628 (.I0(x225), .I1(x226), .I2(x227), .I3(n626), .I4(n627), .O(n628));
  LUT3 #(.INIT(8'h96)) lut_n629 (.I0(n617), .I1(n620), .I2(n621), .O(n629));
  LUT3 #(.INIT(8'hE8)) lut_n630 (.I0(n625), .I1(n628), .I2(n629), .O(n630));
  LUT3 #(.INIT(8'h96)) lut_n631 (.I0(n603), .I1(n611), .I2(n612), .O(n631));
  LUT3 #(.INIT(8'hE8)) lut_n632 (.I0(n622), .I1(n630), .I2(n631), .O(n632));
  LUT3 #(.INIT(8'h96)) lut_n633 (.I0(x234), .I1(x235), .I2(x236), .O(n633));
  LUT5 #(.INIT(32'h96696996)) lut_n634 (.I0(x225), .I1(x226), .I2(x227), .I3(n626), .I4(n627), .O(n634));
  LUT5 #(.INIT(32'hFF969600)) lut_n635 (.I0(x231), .I1(x232), .I2(x233), .I3(n633), .I4(n634), .O(n635));
  LUT3 #(.INIT(8'h96)) lut_n636 (.I0(x240), .I1(x241), .I2(x242), .O(n636));
  LUT5 #(.INIT(32'h96696996)) lut_n637 (.I0(x231), .I1(x232), .I2(x233), .I3(n633), .I4(n634), .O(n637));
  LUT5 #(.INIT(32'hFF969600)) lut_n638 (.I0(x237), .I1(x238), .I2(x239), .I3(n636), .I4(n637), .O(n638));
  LUT3 #(.INIT(8'h96)) lut_n639 (.I0(n625), .I1(n628), .I2(n629), .O(n639));
  LUT3 #(.INIT(8'h96)) lut_n640 (.I0(x246), .I1(x247), .I2(x248), .O(n640));
  LUT5 #(.INIT(32'h96696996)) lut_n641 (.I0(x237), .I1(x238), .I2(x239), .I3(n636), .I4(n637), .O(n641));
  LUT5 #(.INIT(32'hFF969600)) lut_n642 (.I0(x243), .I1(x244), .I2(x245), .I3(n640), .I4(n641), .O(n642));
  LUT3 #(.INIT(8'h96)) lut_n643 (.I0(x249), .I1(x250), .I2(x251), .O(n643));
  LUT5 #(.INIT(32'h96696996)) lut_n644 (.I0(x243), .I1(x244), .I2(x245), .I3(n640), .I4(n641), .O(n644));
  LUT5 #(.INIT(32'hFF969600)) lut_n645 (.I0(x252), .I1(x253), .I2(x254), .I3(n643), .I4(n644), .O(n645));
  LUT3 #(.INIT(8'h96)) lut_n646 (.I0(n622), .I1(n630), .I2(n631), .O(n646));
  LUT6 #(.INIT(64'hFFFEFEE8E8808000)) lut_n647 (.I0(n635), .I1(n638), .I2(n639), .I3(n642), .I4(n645), .I5(n646), .O(n647));
  LUT3 #(.INIT(8'h96)) lut_n648 (.I0(n537), .I1(n575), .I2(n576), .O(n648));
  LUT6 #(.INIT(64'hFFFEFEE8E8808000)) lut_n649 (.I0(n595), .I1(n613), .I2(n614), .I3(n632), .I4(n647), .I5(n648), .O(n649));
  LUT6 #(.INIT(64'hFEEAEAA8EAA8A880)) lut_n650 (.I0(n397), .I1(n435), .I2(n498), .I3(n499), .I4(n577), .I5(n649), .O(n650));
  assign y0 = n650;
endmodule
