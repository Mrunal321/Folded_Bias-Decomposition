module top (x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, y0);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28;
  output y0;
  wire n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63;
  LUT3 #(.INIT(8'hE8)) lut_n31 (.I0(x0), .I1(x1), .I2(x2), .O(n31));
  LUT3 #(.INIT(8'hE8)) lut_n32 (.I0(x6), .I1(x7), .I2(x8), .O(n32));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n33 (.I0(x3), .I1(x4), .I2(x5), .I3(n31), .I4(n32), .O(n33));
  LUT3 #(.INIT(8'hE8)) lut_n34 (.I0(x12), .I1(x13), .I2(x14), .O(n34));
  LUT5 #(.INIT(32'hE81717E8)) lut_n35 (.I0(x3), .I1(x4), .I2(x5), .I3(n31), .I4(n32), .O(n35));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n36 (.I0(x9), .I1(x10), .I2(x11), .I3(n34), .I4(n35), .O(n36));
  LUT3 #(.INIT(8'hE8)) lut_n37 (.I0(x18), .I1(x19), .I2(x20), .O(n37));
  LUT5 #(.INIT(32'hE81717E8)) lut_n38 (.I0(x9), .I1(x10), .I2(x11), .I3(n34), .I4(n35), .O(n38));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n39 (.I0(x15), .I1(x16), .I2(x17), .I3(n37), .I4(n38), .O(n39));
  LUT3 #(.INIT(8'hE8)) lut_n40 (.I0(n33), .I1(n36), .I2(n39), .O(n40));
  LUT3 #(.INIT(8'hE8)) lut_n41 (.I0(x24), .I1(x25), .I2(x26), .O(n41));
  LUT5 #(.INIT(32'hE81717E8)) lut_n42 (.I0(x15), .I1(x16), .I2(x17), .I3(n37), .I4(n38), .O(n42));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n43 (.I0(x21), .I1(x22), .I2(x23), .I3(n41), .I4(n42), .O(n43));
  LUT3 #(.INIT(8'h96)) lut_n44 (.I0(x0), .I1(x1), .I2(x2), .O(n44));
  LUT3 #(.INIT(8'h96)) lut_n45 (.I0(x6), .I1(x7), .I2(x8), .O(n45));
  LUT5 #(.INIT(32'hFF969600)) lut_n46 (.I0(x3), .I1(x4), .I2(x5), .I3(n44), .I4(n45), .O(n46));
  LUT5 #(.INIT(32'hE81717E8)) lut_n47 (.I0(x21), .I1(x22), .I2(x23), .I3(n41), .I4(n42), .O(n47));
  LUT4 #(.INIT(16'hFEE0)) lut_n48 (.I0(x27), .I1(x28), .I2(n46), .I3(n47), .O(n48));
  LUT3 #(.INIT(8'h96)) lut_n49 (.I0(n33), .I1(n36), .I2(n39), .O(n49));
  LUT3 #(.INIT(8'h96)) lut_n50 (.I0(x12), .I1(x13), .I2(x14), .O(n50));
  LUT5 #(.INIT(32'h96696996)) lut_n51 (.I0(x3), .I1(x4), .I2(x5), .I3(n44), .I4(n45), .O(n51));
  LUT5 #(.INIT(32'hFF969600)) lut_n52 (.I0(x9), .I1(x10), .I2(x11), .I3(n50), .I4(n51), .O(n52));
  LUT3 #(.INIT(8'h96)) lut_n53 (.I0(x18), .I1(x19), .I2(x20), .O(n53));
  LUT5 #(.INIT(32'h96696996)) lut_n54 (.I0(x9), .I1(x10), .I2(x11), .I3(n50), .I4(n51), .O(n54));
  LUT5 #(.INIT(32'hFF969600)) lut_n55 (.I0(x15), .I1(x16), .I2(x17), .I3(n53), .I4(n54), .O(n55));
  LUT4 #(.INIT(16'hE11E)) lut_n56 (.I0(x27), .I1(x28), .I2(n46), .I3(n47), .O(n56));
  LUT3 #(.INIT(8'hE8)) lut_n57 (.I0(n52), .I1(n55), .I2(n56), .O(n57));
  LUT3 #(.INIT(8'h96)) lut_n58 (.I0(x21), .I1(x22), .I2(x23), .O(n58));
  LUT3 #(.INIT(8'h96)) lut_n59 (.I0(x24), .I1(x25), .I2(x26), .O(n59));
  LUT5 #(.INIT(32'h96696996)) lut_n60 (.I0(x15), .I1(x16), .I2(x17), .I3(n53), .I4(n54), .O(n60));
  LUT3 #(.INIT(8'h96)) lut_n61 (.I0(n52), .I1(n55), .I2(n56), .O(n61));
  LUT6 #(.INIT(64'hFFF9F99090000000)) lut_n62 (.I0(x27), .I1(x28), .I2(n58), .I3(n59), .I4(n60), .I5(n61), .O(n62));
  LUT6 #(.INIT(64'hFEEAEAA8EAA8A880)) lut_n63 (.I0(n40), .I1(n43), .I2(n48), .I3(n49), .I4(n57), .I5(n62), .O(n63));
  assign y0 = n63;
endmodule
