module top (x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, y0);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54;
  output y0;
  wire n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131;
  LUT3 #(.INIT(8'hE8)) lut_n57 (.I0(x0), .I1(x1), .I2(x2), .O(n57));
  LUT3 #(.INIT(8'hE8)) lut_n58 (.I0(x6), .I1(x7), .I2(x8), .O(n58));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n59 (.I0(x3), .I1(x4), .I2(x5), .I3(n57), .I4(n58), .O(n59));
  LUT3 #(.INIT(8'hE8)) lut_n60 (.I0(x12), .I1(x13), .I2(x14), .O(n60));
  LUT5 #(.INIT(32'hE81717E8)) lut_n61 (.I0(x3), .I1(x4), .I2(x5), .I3(n57), .I4(n58), .O(n61));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n62 (.I0(x9), .I1(x10), .I2(x11), .I3(n60), .I4(n61), .O(n62));
  LUT3 #(.INIT(8'hE8)) lut_n63 (.I0(x18), .I1(x19), .I2(x20), .O(n63));
  LUT5 #(.INIT(32'hE81717E8)) lut_n64 (.I0(x9), .I1(x10), .I2(x11), .I3(n60), .I4(n61), .O(n64));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n65 (.I0(x15), .I1(x16), .I2(x17), .I3(n63), .I4(n64), .O(n65));
  LUT3 #(.INIT(8'hE8)) lut_n66 (.I0(n59), .I1(n62), .I2(n65), .O(n66));
  LUT3 #(.INIT(8'hE8)) lut_n67 (.I0(x24), .I1(x25), .I2(x26), .O(n67));
  LUT5 #(.INIT(32'hE81717E8)) lut_n68 (.I0(x15), .I1(x16), .I2(x17), .I3(n63), .I4(n64), .O(n68));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n69 (.I0(x21), .I1(x22), .I2(x23), .I3(n67), .I4(n68), .O(n69));
  LUT3 #(.INIT(8'hE8)) lut_n70 (.I0(x27), .I1(x28), .I2(x29), .O(n70));
  LUT5 #(.INIT(32'hE81717E8)) lut_n71 (.I0(x21), .I1(x22), .I2(x23), .I3(n67), .I4(n68), .O(n71));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n72 (.I0(x30), .I1(x31), .I2(x32), .I3(n70), .I4(n71), .O(n72));
  LUT3 #(.INIT(8'h96)) lut_n73 (.I0(n59), .I1(n62), .I2(n65), .O(n73));
  LUT3 #(.INIT(8'hE8)) lut_n74 (.I0(n69), .I1(n72), .I2(n73), .O(n74));
  LUT3 #(.INIT(8'hE8)) lut_n75 (.I0(x36), .I1(x37), .I2(x38), .O(n75));
  LUT5 #(.INIT(32'hE81717E8)) lut_n76 (.I0(x30), .I1(x31), .I2(x32), .I3(n70), .I4(n71), .O(n76));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n77 (.I0(x33), .I1(x34), .I2(x35), .I3(n75), .I4(n76), .O(n77));
  LUT3 #(.INIT(8'hE8)) lut_n78 (.I0(x42), .I1(x43), .I2(x44), .O(n78));
  LUT5 #(.INIT(32'hE81717E8)) lut_n79 (.I0(x33), .I1(x34), .I2(x35), .I3(n75), .I4(n76), .O(n79));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n80 (.I0(x39), .I1(x40), .I2(x41), .I3(n78), .I4(n79), .O(n80));
  LUT3 #(.INIT(8'h96)) lut_n81 (.I0(n69), .I1(n72), .I2(n73), .O(n81));
  LUT3 #(.INIT(8'hE8)) lut_n82 (.I0(n77), .I1(n80), .I2(n81), .O(n82));
  LUT3 #(.INIT(8'hE8)) lut_n83 (.I0(n66), .I1(n74), .I2(n82), .O(n83));
  LUT3 #(.INIT(8'hE8)) lut_n84 (.I0(x48), .I1(x49), .I2(x50), .O(n84));
  LUT5 #(.INIT(32'hE81717E8)) lut_n85 (.I0(x39), .I1(x40), .I2(x41), .I3(n78), .I4(n79), .O(n85));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n86 (.I0(x45), .I1(x46), .I2(x47), .I3(n84), .I4(n85), .O(n86));
  LUT5 #(.INIT(32'hE81717E8)) lut_n87 (.I0(x45), .I1(x46), .I2(x47), .I3(n84), .I4(n85), .O(n87));
  LUT4 #(.INIT(16'hFFE8)) lut_n88 (.I0(x51), .I1(x52), .I2(x53), .I3(n87), .O(n88));
  LUT3 #(.INIT(8'h96)) lut_n89 (.I0(n77), .I1(n80), .I2(n81), .O(n89));
  LUT3 #(.INIT(8'hE8)) lut_n90 (.I0(n86), .I1(n88), .I2(n89), .O(n90));
  LUT4 #(.INIT(16'h17E8)) lut_n91 (.I0(x51), .I1(x52), .I2(x53), .I3(n87), .O(n91));
  LUT3 #(.INIT(8'h96)) lut_n92 (.I0(x0), .I1(x1), .I2(x2), .O(n92));
  LUT3 #(.INIT(8'h96)) lut_n93 (.I0(x6), .I1(x7), .I2(x8), .O(n93));
  LUT5 #(.INIT(32'hFF969600)) lut_n94 (.I0(x3), .I1(x4), .I2(x5), .I3(n92), .I4(n93), .O(n94));
  LUT3 #(.INIT(8'h96)) lut_n95 (.I0(x12), .I1(x13), .I2(x14), .O(n95));
  LUT5 #(.INIT(32'h96696996)) lut_n96 (.I0(x3), .I1(x4), .I2(x5), .I3(n92), .I4(n93), .O(n96));
  LUT5 #(.INIT(32'hFF969600)) lut_n97 (.I0(x9), .I1(x10), .I2(x11), .I3(n95), .I4(n96), .O(n97));
  LUT3 #(.INIT(8'hE8)) lut_n98 (.I0(n91), .I1(n94), .I2(n97), .O(n98));
  LUT3 #(.INIT(8'h96)) lut_n99 (.I0(n86), .I1(n88), .I2(n89), .O(n99));
  LUT3 #(.INIT(8'hD4)) lut_n100 (.I0(n91), .I1(n98), .I2(n99), .O(n100));
  LUT3 #(.INIT(8'h96)) lut_n101 (.I0(n66), .I1(n74), .I2(n82), .O(n101));
  LUT3 #(.INIT(8'h96)) lut_n102 (.I0(x18), .I1(x19), .I2(x20), .O(n102));
  LUT5 #(.INIT(32'h96696996)) lut_n103 (.I0(x9), .I1(x10), .I2(x11), .I3(n95), .I4(n96), .O(n103));
  LUT5 #(.INIT(32'hFF969600)) lut_n104 (.I0(x15), .I1(x16), .I2(x17), .I3(n102), .I4(n103), .O(n104));
  LUT3 #(.INIT(8'h96)) lut_n105 (.I0(x24), .I1(x25), .I2(x26), .O(n105));
  LUT5 #(.INIT(32'h96696996)) lut_n106 (.I0(x15), .I1(x16), .I2(x17), .I3(n102), .I4(n103), .O(n106));
  LUT5 #(.INIT(32'hFF969600)) lut_n107 (.I0(x21), .I1(x22), .I2(x23), .I3(n105), .I4(n106), .O(n107));
  LUT3 #(.INIT(8'h96)) lut_n108 (.I0(n91), .I1(n94), .I2(n97), .O(n108));
  LUT3 #(.INIT(8'hE8)) lut_n109 (.I0(n104), .I1(n107), .I2(n108), .O(n109));
  LUT3 #(.INIT(8'h96)) lut_n110 (.I0(x27), .I1(x28), .I2(x29), .O(n110));
  LUT5 #(.INIT(32'h96696996)) lut_n111 (.I0(x21), .I1(x22), .I2(x23), .I3(n105), .I4(n106), .O(n111));
  LUT5 #(.INIT(32'hFF969600)) lut_n112 (.I0(x30), .I1(x31), .I2(x32), .I3(n110), .I4(n111), .O(n112));
  LUT3 #(.INIT(8'h96)) lut_n113 (.I0(x36), .I1(x37), .I2(x38), .O(n113));
  LUT5 #(.INIT(32'h96696996)) lut_n114 (.I0(x30), .I1(x31), .I2(x32), .I3(n110), .I4(n111), .O(n114));
  LUT5 #(.INIT(32'hFF969600)) lut_n115 (.I0(x33), .I1(x34), .I2(x35), .I3(n113), .I4(n114), .O(n115));
  LUT3 #(.INIT(8'h96)) lut_n116 (.I0(n104), .I1(n107), .I2(n108), .O(n116));
  LUT3 #(.INIT(8'hE8)) lut_n117 (.I0(n112), .I1(n115), .I2(n116), .O(n117));
  LUT3 #(.INIT(8'h96)) lut_n118 (.I0(n91), .I1(n98), .I2(n99), .O(n118));
  LUT3 #(.INIT(8'h8E)) lut_n119 (.I0(n109), .I1(n117), .I2(n118), .O(n119));
  LUT3 #(.INIT(8'h96)) lut_n120 (.I0(x42), .I1(x43), .I2(x44), .O(n120));
  LUT5 #(.INIT(32'h96696996)) lut_n121 (.I0(x33), .I1(x34), .I2(x35), .I3(n113), .I4(n114), .O(n121));
  LUT5 #(.INIT(32'hFF969600)) lut_n122 (.I0(x39), .I1(x40), .I2(x41), .I3(n120), .I4(n121), .O(n122));
  LUT3 #(.INIT(8'h96)) lut_n123 (.I0(x48), .I1(x49), .I2(x50), .O(n123));
  LUT5 #(.INIT(32'h96696996)) lut_n124 (.I0(x39), .I1(x40), .I2(x41), .I3(n120), .I4(n121), .O(n124));
  LUT5 #(.INIT(32'hFF969600)) lut_n125 (.I0(x45), .I1(x46), .I2(x47), .I3(n123), .I4(n124), .O(n125));
  LUT3 #(.INIT(8'h96)) lut_n126 (.I0(n112), .I1(n115), .I2(n116), .O(n126));
  LUT5 #(.INIT(32'h96696996)) lut_n127 (.I0(x45), .I1(x46), .I2(x47), .I3(n123), .I4(n124), .O(n127));
  LUT5 #(.INIT(32'hFF969600)) lut_n128 (.I0(x51), .I1(x52), .I2(x53), .I3(x54), .I4(n127), .O(n128));
  LUT3 #(.INIT(8'h96)) lut_n129 (.I0(n109), .I1(n117), .I2(n118), .O(n129));
  LUT5 #(.INIT(32'h8000FEE8)) lut_n130 (.I0(n122), .I1(n125), .I2(n126), .I3(n128), .I4(n129), .O(n130));
  LUT6 #(.INIT(64'hFEEAEAA8EAA8A880)) lut_n131 (.I0(n83), .I1(n90), .I2(n100), .I3(n101), .I4(n119), .I5(n130), .O(n131));
  assign y0 = n131;
endmodule
