module top (x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, y0);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126;
  output y0;
  wire n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313;
  LUT3 #(.INIT(8'hE8)) lut_n129 (.I0(x0), .I1(x1), .I2(x2), .O(n129));
  LUT3 #(.INIT(8'hE8)) lut_n130 (.I0(x6), .I1(x7), .I2(x8), .O(n130));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n131 (.I0(x3), .I1(x4), .I2(x5), .I3(n129), .I4(n130), .O(n131));
  LUT3 #(.INIT(8'hE8)) lut_n132 (.I0(x12), .I1(x13), .I2(x14), .O(n132));
  LUT5 #(.INIT(32'hE81717E8)) lut_n133 (.I0(x3), .I1(x4), .I2(x5), .I3(n129), .I4(n130), .O(n133));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n134 (.I0(x9), .I1(x10), .I2(x11), .I3(n132), .I4(n133), .O(n134));
  LUT3 #(.INIT(8'hE8)) lut_n135 (.I0(x18), .I1(x19), .I2(x20), .O(n135));
  LUT5 #(.INIT(32'hE81717E8)) lut_n136 (.I0(x9), .I1(x10), .I2(x11), .I3(n132), .I4(n133), .O(n136));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n137 (.I0(x15), .I1(x16), .I2(x17), .I3(n135), .I4(n136), .O(n137));
  LUT3 #(.INIT(8'hE8)) lut_n138 (.I0(n131), .I1(n134), .I2(n137), .O(n138));
  LUT3 #(.INIT(8'hE8)) lut_n139 (.I0(x24), .I1(x25), .I2(x26), .O(n139));
  LUT5 #(.INIT(32'hE81717E8)) lut_n140 (.I0(x15), .I1(x16), .I2(x17), .I3(n135), .I4(n136), .O(n140));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n141 (.I0(x21), .I1(x22), .I2(x23), .I3(n139), .I4(n140), .O(n141));
  LUT3 #(.INIT(8'hE8)) lut_n142 (.I0(x27), .I1(x28), .I2(x29), .O(n142));
  LUT5 #(.INIT(32'hE81717E8)) lut_n143 (.I0(x21), .I1(x22), .I2(x23), .I3(n139), .I4(n140), .O(n143));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n144 (.I0(x30), .I1(x31), .I2(x32), .I3(n142), .I4(n143), .O(n144));
  LUT3 #(.INIT(8'h96)) lut_n145 (.I0(n131), .I1(n134), .I2(n137), .O(n145));
  LUT3 #(.INIT(8'hE8)) lut_n146 (.I0(n141), .I1(n144), .I2(n145), .O(n146));
  LUT3 #(.INIT(8'hE8)) lut_n147 (.I0(x36), .I1(x37), .I2(x38), .O(n147));
  LUT5 #(.INIT(32'hE81717E8)) lut_n148 (.I0(x30), .I1(x31), .I2(x32), .I3(n142), .I4(n143), .O(n148));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n149 (.I0(x33), .I1(x34), .I2(x35), .I3(n147), .I4(n148), .O(n149));
  LUT3 #(.INIT(8'hE8)) lut_n150 (.I0(x42), .I1(x43), .I2(x44), .O(n150));
  LUT5 #(.INIT(32'hE81717E8)) lut_n151 (.I0(x33), .I1(x34), .I2(x35), .I3(n147), .I4(n148), .O(n151));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n152 (.I0(x39), .I1(x40), .I2(x41), .I3(n150), .I4(n151), .O(n152));
  LUT3 #(.INIT(8'h96)) lut_n153 (.I0(n141), .I1(n144), .I2(n145), .O(n153));
  LUT3 #(.INIT(8'hE8)) lut_n154 (.I0(n149), .I1(n152), .I2(n153), .O(n154));
  LUT3 #(.INIT(8'hE8)) lut_n155 (.I0(n138), .I1(n146), .I2(n154), .O(n155));
  LUT3 #(.INIT(8'hE8)) lut_n156 (.I0(x48), .I1(x49), .I2(x50), .O(n156));
  LUT5 #(.INIT(32'hE81717E8)) lut_n157 (.I0(x39), .I1(x40), .I2(x41), .I3(n150), .I4(n151), .O(n157));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n158 (.I0(x45), .I1(x46), .I2(x47), .I3(n156), .I4(n157), .O(n158));
  LUT3 #(.INIT(8'hE8)) lut_n159 (.I0(x54), .I1(x55), .I2(x56), .O(n159));
  LUT5 #(.INIT(32'hE81717E8)) lut_n160 (.I0(x45), .I1(x46), .I2(x47), .I3(n156), .I4(n157), .O(n160));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n161 (.I0(x51), .I1(x52), .I2(x53), .I3(n159), .I4(n160), .O(n161));
  LUT3 #(.INIT(8'h96)) lut_n162 (.I0(n149), .I1(n152), .I2(n153), .O(n162));
  LUT3 #(.INIT(8'hE8)) lut_n163 (.I0(n158), .I1(n161), .I2(n162), .O(n163));
  LUT3 #(.INIT(8'hE8)) lut_n164 (.I0(x60), .I1(x61), .I2(x62), .O(n164));
  LUT5 #(.INIT(32'hE81717E8)) lut_n165 (.I0(x51), .I1(x52), .I2(x53), .I3(n159), .I4(n160), .O(n165));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n166 (.I0(x57), .I1(x58), .I2(x59), .I3(n164), .I4(n165), .O(n166));
  LUT3 #(.INIT(8'hE8)) lut_n167 (.I0(x66), .I1(x67), .I2(x68), .O(n167));
  LUT5 #(.INIT(32'hE81717E8)) lut_n168 (.I0(x57), .I1(x58), .I2(x59), .I3(n164), .I4(n165), .O(n168));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n169 (.I0(x63), .I1(x64), .I2(x65), .I3(n167), .I4(n168), .O(n169));
  LUT3 #(.INIT(8'h96)) lut_n170 (.I0(n158), .I1(n161), .I2(n162), .O(n170));
  LUT3 #(.INIT(8'hE8)) lut_n171 (.I0(n166), .I1(n169), .I2(n170), .O(n171));
  LUT3 #(.INIT(8'h96)) lut_n172 (.I0(n138), .I1(n146), .I2(n154), .O(n172));
  LUT3 #(.INIT(8'hE8)) lut_n173 (.I0(n163), .I1(n171), .I2(n172), .O(n173));
  LUT3 #(.INIT(8'hE8)) lut_n174 (.I0(x72), .I1(x73), .I2(x74), .O(n174));
  LUT5 #(.INIT(32'hE81717E8)) lut_n175 (.I0(x63), .I1(x64), .I2(x65), .I3(n167), .I4(n168), .O(n175));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n176 (.I0(x69), .I1(x70), .I2(x71), .I3(n174), .I4(n175), .O(n176));
  LUT3 #(.INIT(8'hE8)) lut_n177 (.I0(x78), .I1(x79), .I2(x80), .O(n177));
  LUT5 #(.INIT(32'hE81717E8)) lut_n178 (.I0(x69), .I1(x70), .I2(x71), .I3(n174), .I4(n175), .O(n178));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n179 (.I0(x75), .I1(x76), .I2(x77), .I3(n177), .I4(n178), .O(n179));
  LUT3 #(.INIT(8'h96)) lut_n180 (.I0(n166), .I1(n169), .I2(n170), .O(n180));
  LUT3 #(.INIT(8'hE8)) lut_n181 (.I0(n176), .I1(n179), .I2(n180), .O(n181));
  LUT3 #(.INIT(8'hE8)) lut_n182 (.I0(x84), .I1(x85), .I2(x86), .O(n182));
  LUT5 #(.INIT(32'hE81717E8)) lut_n183 (.I0(x75), .I1(x76), .I2(x77), .I3(n177), .I4(n178), .O(n183));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n184 (.I0(x81), .I1(x82), .I2(x83), .I3(n182), .I4(n183), .O(n184));
  LUT3 #(.INIT(8'hE8)) lut_n185 (.I0(x90), .I1(x91), .I2(x92), .O(n185));
  LUT5 #(.INIT(32'hE81717E8)) lut_n186 (.I0(x81), .I1(x82), .I2(x83), .I3(n182), .I4(n183), .O(n186));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n187 (.I0(x87), .I1(x88), .I2(x89), .I3(n185), .I4(n186), .O(n187));
  LUT3 #(.INIT(8'h96)) lut_n188 (.I0(n176), .I1(n179), .I2(n180), .O(n188));
  LUT3 #(.INIT(8'hE8)) lut_n189 (.I0(n184), .I1(n187), .I2(n188), .O(n189));
  LUT3 #(.INIT(8'h96)) lut_n190 (.I0(n163), .I1(n171), .I2(n172), .O(n190));
  LUT3 #(.INIT(8'hE8)) lut_n191 (.I0(n181), .I1(n189), .I2(n190), .O(n191));
  LUT3 #(.INIT(8'hE8)) lut_n192 (.I0(n155), .I1(n173), .I2(n191), .O(n192));
  LUT3 #(.INIT(8'hE8)) lut_n193 (.I0(x96), .I1(x97), .I2(x98), .O(n193));
  LUT5 #(.INIT(32'hE81717E8)) lut_n194 (.I0(x87), .I1(x88), .I2(x89), .I3(n185), .I4(n186), .O(n194));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n195 (.I0(x93), .I1(x94), .I2(x95), .I3(n193), .I4(n194), .O(n195));
  LUT3 #(.INIT(8'hE8)) lut_n196 (.I0(x102), .I1(x103), .I2(x104), .O(n196));
  LUT5 #(.INIT(32'hE81717E8)) lut_n197 (.I0(x93), .I1(x94), .I2(x95), .I3(n193), .I4(n194), .O(n197));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n198 (.I0(x99), .I1(x100), .I2(x101), .I3(n196), .I4(n197), .O(n198));
  LUT3 #(.INIT(8'h96)) lut_n199 (.I0(n184), .I1(n187), .I2(n188), .O(n199));
  LUT3 #(.INIT(8'hE8)) lut_n200 (.I0(n195), .I1(n198), .I2(n199), .O(n200));
  LUT3 #(.INIT(8'hE8)) lut_n201 (.I0(x108), .I1(x109), .I2(x110), .O(n201));
  LUT5 #(.INIT(32'hE81717E8)) lut_n202 (.I0(x99), .I1(x100), .I2(x101), .I3(n196), .I4(n197), .O(n202));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n203 (.I0(x105), .I1(x106), .I2(x107), .I3(n201), .I4(n202), .O(n203));
  LUT3 #(.INIT(8'hE8)) lut_n204 (.I0(x114), .I1(x115), .I2(x116), .O(n204));
  LUT5 #(.INIT(32'hE81717E8)) lut_n205 (.I0(x105), .I1(x106), .I2(x107), .I3(n201), .I4(n202), .O(n205));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n206 (.I0(x111), .I1(x112), .I2(x113), .I3(n204), .I4(n205), .O(n206));
  LUT3 #(.INIT(8'h96)) lut_n207 (.I0(n195), .I1(n198), .I2(n199), .O(n207));
  LUT3 #(.INIT(8'hE8)) lut_n208 (.I0(n203), .I1(n206), .I2(n207), .O(n208));
  LUT3 #(.INIT(8'h96)) lut_n209 (.I0(n181), .I1(n189), .I2(n190), .O(n209));
  LUT3 #(.INIT(8'hE8)) lut_n210 (.I0(n200), .I1(n208), .I2(n209), .O(n210));
  LUT3 #(.INIT(8'hE8)) lut_n211 (.I0(x120), .I1(x121), .I2(x122), .O(n211));
  LUT5 #(.INIT(32'hE81717E8)) lut_n212 (.I0(x111), .I1(x112), .I2(x113), .I3(n204), .I4(n205), .O(n212));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n213 (.I0(x117), .I1(x118), .I2(x119), .I3(n211), .I4(n212), .O(n213));
  LUT3 #(.INIT(8'h96)) lut_n214 (.I0(x0), .I1(x1), .I2(x2), .O(n214));
  LUT3 #(.INIT(8'h96)) lut_n215 (.I0(x6), .I1(x7), .I2(x8), .O(n215));
  LUT5 #(.INIT(32'hFF969600)) lut_n216 (.I0(x3), .I1(x4), .I2(x5), .I3(n214), .I4(n215), .O(n216));
  LUT5 #(.INIT(32'hE81717E8)) lut_n217 (.I0(x117), .I1(x118), .I2(x119), .I3(n211), .I4(n212), .O(n217));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n218 (.I0(x123), .I1(x124), .I2(x125), .I3(n216), .I4(n217), .O(n218));
  LUT3 #(.INIT(8'h96)) lut_n219 (.I0(n203), .I1(n206), .I2(n207), .O(n219));
  LUT3 #(.INIT(8'hE8)) lut_n220 (.I0(n213), .I1(n218), .I2(n219), .O(n220));
  LUT3 #(.INIT(8'h96)) lut_n221 (.I0(x12), .I1(x13), .I2(x14), .O(n221));
  LUT5 #(.INIT(32'h96696996)) lut_n222 (.I0(x3), .I1(x4), .I2(x5), .I3(n214), .I4(n215), .O(n222));
  LUT5 #(.INIT(32'hFF969600)) lut_n223 (.I0(x9), .I1(x10), .I2(x11), .I3(n221), .I4(n222), .O(n223));
  LUT3 #(.INIT(8'h96)) lut_n224 (.I0(x18), .I1(x19), .I2(x20), .O(n224));
  LUT5 #(.INIT(32'h96696996)) lut_n225 (.I0(x9), .I1(x10), .I2(x11), .I3(n221), .I4(n222), .O(n225));
  LUT5 #(.INIT(32'hFF969600)) lut_n226 (.I0(x15), .I1(x16), .I2(x17), .I3(n224), .I4(n225), .O(n226));
  LUT5 #(.INIT(32'hE81717E8)) lut_n227 (.I0(x123), .I1(x124), .I2(x125), .I3(n216), .I4(n217), .O(n227));
  LUT3 #(.INIT(8'hE8)) lut_n228 (.I0(n223), .I1(n226), .I2(n227), .O(n228));
  LUT3 #(.INIT(8'h96)) lut_n229 (.I0(x24), .I1(x25), .I2(x26), .O(n229));
  LUT5 #(.INIT(32'h96696996)) lut_n230 (.I0(x15), .I1(x16), .I2(x17), .I3(n224), .I4(n225), .O(n230));
  LUT5 #(.INIT(32'hFF969600)) lut_n231 (.I0(x21), .I1(x22), .I2(x23), .I3(n229), .I4(n230), .O(n231));
  LUT3 #(.INIT(8'h96)) lut_n232 (.I0(x27), .I1(x28), .I2(x29), .O(n232));
  LUT5 #(.INIT(32'h96696996)) lut_n233 (.I0(x21), .I1(x22), .I2(x23), .I3(n229), .I4(n230), .O(n233));
  LUT5 #(.INIT(32'hFF969600)) lut_n234 (.I0(x30), .I1(x31), .I2(x32), .I3(n232), .I4(n233), .O(n234));
  LUT3 #(.INIT(8'h96)) lut_n235 (.I0(n223), .I1(n226), .I2(n227), .O(n235));
  LUT3 #(.INIT(8'hE8)) lut_n236 (.I0(n231), .I1(n234), .I2(n235), .O(n236));
  LUT3 #(.INIT(8'h96)) lut_n237 (.I0(n213), .I1(n218), .I2(n219), .O(n237));
  LUT3 #(.INIT(8'hE8)) lut_n238 (.I0(n228), .I1(n236), .I2(n237), .O(n238));
  LUT3 #(.INIT(8'h96)) lut_n239 (.I0(n200), .I1(n208), .I2(n209), .O(n239));
  LUT3 #(.INIT(8'hE8)) lut_n240 (.I0(n220), .I1(n238), .I2(n239), .O(n240));
  LUT3 #(.INIT(8'h96)) lut_n241 (.I0(n155), .I1(n173), .I2(n191), .O(n241));
  LUT3 #(.INIT(8'h96)) lut_n242 (.I0(x36), .I1(x37), .I2(x38), .O(n242));
  LUT5 #(.INIT(32'h96696996)) lut_n243 (.I0(x30), .I1(x31), .I2(x32), .I3(n232), .I4(n233), .O(n243));
  LUT5 #(.INIT(32'hFF969600)) lut_n244 (.I0(x33), .I1(x34), .I2(x35), .I3(n242), .I4(n243), .O(n244));
  LUT3 #(.INIT(8'h96)) lut_n245 (.I0(x42), .I1(x43), .I2(x44), .O(n245));
  LUT5 #(.INIT(32'h96696996)) lut_n246 (.I0(x33), .I1(x34), .I2(x35), .I3(n242), .I4(n243), .O(n246));
  LUT5 #(.INIT(32'hFF969600)) lut_n247 (.I0(x39), .I1(x40), .I2(x41), .I3(n245), .I4(n246), .O(n247));
  LUT3 #(.INIT(8'h96)) lut_n248 (.I0(n231), .I1(n234), .I2(n235), .O(n248));
  LUT3 #(.INIT(8'hE8)) lut_n249 (.I0(n244), .I1(n247), .I2(n248), .O(n249));
  LUT3 #(.INIT(8'h96)) lut_n250 (.I0(x48), .I1(x49), .I2(x50), .O(n250));
  LUT5 #(.INIT(32'h96696996)) lut_n251 (.I0(x39), .I1(x40), .I2(x41), .I3(n245), .I4(n246), .O(n251));
  LUT5 #(.INIT(32'hFF969600)) lut_n252 (.I0(x45), .I1(x46), .I2(x47), .I3(n250), .I4(n251), .O(n252));
  LUT3 #(.INIT(8'h96)) lut_n253 (.I0(x54), .I1(x55), .I2(x56), .O(n253));
  LUT5 #(.INIT(32'h96696996)) lut_n254 (.I0(x45), .I1(x46), .I2(x47), .I3(n250), .I4(n251), .O(n254));
  LUT5 #(.INIT(32'hFF969600)) lut_n255 (.I0(x51), .I1(x52), .I2(x53), .I3(n253), .I4(n254), .O(n255));
  LUT3 #(.INIT(8'h96)) lut_n256 (.I0(n244), .I1(n247), .I2(n248), .O(n256));
  LUT3 #(.INIT(8'hE8)) lut_n257 (.I0(n252), .I1(n255), .I2(n256), .O(n257));
  LUT3 #(.INIT(8'h96)) lut_n258 (.I0(n228), .I1(n236), .I2(n237), .O(n258));
  LUT3 #(.INIT(8'hE8)) lut_n259 (.I0(n249), .I1(n257), .I2(n258), .O(n259));
  LUT3 #(.INIT(8'h96)) lut_n260 (.I0(x60), .I1(x61), .I2(x62), .O(n260));
  LUT5 #(.INIT(32'h96696996)) lut_n261 (.I0(x51), .I1(x52), .I2(x53), .I3(n253), .I4(n254), .O(n261));
  LUT5 #(.INIT(32'hFF969600)) lut_n262 (.I0(x57), .I1(x58), .I2(x59), .I3(n260), .I4(n261), .O(n262));
  LUT3 #(.INIT(8'h96)) lut_n263 (.I0(x66), .I1(x67), .I2(x68), .O(n263));
  LUT5 #(.INIT(32'h96696996)) lut_n264 (.I0(x57), .I1(x58), .I2(x59), .I3(n260), .I4(n261), .O(n264));
  LUT5 #(.INIT(32'hFF969600)) lut_n265 (.I0(x63), .I1(x64), .I2(x65), .I3(n263), .I4(n264), .O(n265));
  LUT3 #(.INIT(8'h96)) lut_n266 (.I0(n252), .I1(n255), .I2(n256), .O(n266));
  LUT3 #(.INIT(8'hE8)) lut_n267 (.I0(n262), .I1(n265), .I2(n266), .O(n267));
  LUT3 #(.INIT(8'h96)) lut_n268 (.I0(x72), .I1(x73), .I2(x74), .O(n268));
  LUT5 #(.INIT(32'h96696996)) lut_n269 (.I0(x63), .I1(x64), .I2(x65), .I3(n263), .I4(n264), .O(n269));
  LUT5 #(.INIT(32'hFF969600)) lut_n270 (.I0(x69), .I1(x70), .I2(x71), .I3(n268), .I4(n269), .O(n270));
  LUT3 #(.INIT(8'h96)) lut_n271 (.I0(x78), .I1(x79), .I2(x80), .O(n271));
  LUT5 #(.INIT(32'h96696996)) lut_n272 (.I0(x69), .I1(x70), .I2(x71), .I3(n268), .I4(n269), .O(n272));
  LUT5 #(.INIT(32'hFF969600)) lut_n273 (.I0(x75), .I1(x76), .I2(x77), .I3(n271), .I4(n272), .O(n273));
  LUT3 #(.INIT(8'h96)) lut_n274 (.I0(n262), .I1(n265), .I2(n266), .O(n274));
  LUT3 #(.INIT(8'hE8)) lut_n275 (.I0(n270), .I1(n273), .I2(n274), .O(n275));
  LUT3 #(.INIT(8'h96)) lut_n276 (.I0(n249), .I1(n257), .I2(n258), .O(n276));
  LUT3 #(.INIT(8'hE8)) lut_n277 (.I0(n267), .I1(n275), .I2(n276), .O(n277));
  LUT3 #(.INIT(8'h96)) lut_n278 (.I0(n220), .I1(n238), .I2(n239), .O(n278));
  LUT3 #(.INIT(8'hE8)) lut_n279 (.I0(n259), .I1(n277), .I2(n278), .O(n279));
  LUT3 #(.INIT(8'h96)) lut_n280 (.I0(x84), .I1(x85), .I2(x86), .O(n280));
  LUT5 #(.INIT(32'h96696996)) lut_n281 (.I0(x75), .I1(x76), .I2(x77), .I3(n271), .I4(n272), .O(n281));
  LUT5 #(.INIT(32'hFF969600)) lut_n282 (.I0(x81), .I1(x82), .I2(x83), .I3(n280), .I4(n281), .O(n282));
  LUT3 #(.INIT(8'h96)) lut_n283 (.I0(x90), .I1(x91), .I2(x92), .O(n283));
  LUT5 #(.INIT(32'h96696996)) lut_n284 (.I0(x81), .I1(x82), .I2(x83), .I3(n280), .I4(n281), .O(n284));
  LUT5 #(.INIT(32'hFF969600)) lut_n285 (.I0(x87), .I1(x88), .I2(x89), .I3(n283), .I4(n284), .O(n285));
  LUT3 #(.INIT(8'h96)) lut_n286 (.I0(n270), .I1(n273), .I2(n274), .O(n286));
  LUT3 #(.INIT(8'hE8)) lut_n287 (.I0(n282), .I1(n285), .I2(n286), .O(n287));
  LUT3 #(.INIT(8'h96)) lut_n288 (.I0(x96), .I1(x97), .I2(x98), .O(n288));
  LUT5 #(.INIT(32'h96696996)) lut_n289 (.I0(x87), .I1(x88), .I2(x89), .I3(n283), .I4(n284), .O(n289));
  LUT5 #(.INIT(32'hFF969600)) lut_n290 (.I0(x93), .I1(x94), .I2(x95), .I3(n288), .I4(n289), .O(n290));
  LUT3 #(.INIT(8'h96)) lut_n291 (.I0(x102), .I1(x103), .I2(x104), .O(n291));
  LUT5 #(.INIT(32'h96696996)) lut_n292 (.I0(x93), .I1(x94), .I2(x95), .I3(n288), .I4(n289), .O(n292));
  LUT5 #(.INIT(32'hFF969600)) lut_n293 (.I0(x99), .I1(x100), .I2(x101), .I3(n291), .I4(n292), .O(n293));
  LUT3 #(.INIT(8'h96)) lut_n294 (.I0(n282), .I1(n285), .I2(n286), .O(n294));
  LUT3 #(.INIT(8'hE8)) lut_n295 (.I0(n290), .I1(n293), .I2(n294), .O(n295));
  LUT3 #(.INIT(8'h96)) lut_n296 (.I0(n267), .I1(n275), .I2(n276), .O(n296));
  LUT3 #(.INIT(8'h96)) lut_n297 (.I0(x108), .I1(x109), .I2(x110), .O(n297));
  LUT5 #(.INIT(32'h96696996)) lut_n298 (.I0(x99), .I1(x100), .I2(x101), .I3(n291), .I4(n292), .O(n298));
  LUT5 #(.INIT(32'hFF969600)) lut_n299 (.I0(x105), .I1(x106), .I2(x107), .I3(n297), .I4(n298), .O(n299));
  LUT3 #(.INIT(8'h96)) lut_n300 (.I0(x114), .I1(x115), .I2(x116), .O(n300));
  LUT5 #(.INIT(32'h96696996)) lut_n301 (.I0(x105), .I1(x106), .I2(x107), .I3(n297), .I4(n298), .O(n301));
  LUT5 #(.INIT(32'hFF969600)) lut_n302 (.I0(x111), .I1(x112), .I2(x113), .I3(n300), .I4(n301), .O(n302));
  LUT3 #(.INIT(8'h96)) lut_n303 (.I0(n290), .I1(n293), .I2(n294), .O(n303));
  LUT3 #(.INIT(8'hE8)) lut_n304 (.I0(n299), .I1(n302), .I2(n303), .O(n304));
  LUT3 #(.INIT(8'h96)) lut_n305 (.I0(x117), .I1(x118), .I2(x119), .O(n305));
  LUT3 #(.INIT(8'h96)) lut_n306 (.I0(x120), .I1(x121), .I2(x122), .O(n306));
  LUT5 #(.INIT(32'h96696996)) lut_n307 (.I0(x111), .I1(x112), .I2(x113), .I3(n300), .I4(n301), .O(n307));
  LUT3 #(.INIT(8'h96)) lut_n308 (.I0(x123), .I1(x124), .I2(x125), .O(n308));
  LUT3 #(.INIT(8'h96)) lut_n309 (.I0(n299), .I1(n302), .I2(n303), .O(n309));
  LUT6 #(.INIT(64'hFFFEFEE8E8808000)) lut_n310 (.I0(x126), .I1(n305), .I2(n306), .I3(n307), .I4(n308), .I5(n309), .O(n310));
  LUT3 #(.INIT(8'h96)) lut_n311 (.I0(n259), .I1(n277), .I2(n278), .O(n311));
  LUT6 #(.INIT(64'hFFFEFEE8E8808000)) lut_n312 (.I0(n287), .I1(n295), .I2(n296), .I3(n304), .I4(n310), .I5(n311), .O(n312));
  LUT6 #(.INIT(64'hFEEAEAA8EAA8A880)) lut_n313 (.I0(n192), .I1(n210), .I2(n240), .I3(n241), .I4(n279), .I5(n312), .O(n313));
  assign y0 = n313;
endmodule
