module top (x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, y0);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62;
  output y0;
  wire n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147;
  LUT3 #(.INIT(8'hE8)) lut_n65 (.I0(x0), .I1(x1), .I2(x2), .O(n65));
  LUT3 #(.INIT(8'hE8)) lut_n66 (.I0(x6), .I1(x7), .I2(x8), .O(n66));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n67 (.I0(x3), .I1(x4), .I2(x5), .I3(n65), .I4(n66), .O(n67));
  LUT3 #(.INIT(8'hE8)) lut_n68 (.I0(x12), .I1(x13), .I2(x14), .O(n68));
  LUT5 #(.INIT(32'hE81717E8)) lut_n69 (.I0(x3), .I1(x4), .I2(x5), .I3(n65), .I4(n66), .O(n69));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n70 (.I0(x9), .I1(x10), .I2(x11), .I3(n68), .I4(n69), .O(n70));
  LUT3 #(.INIT(8'hE8)) lut_n71 (.I0(x18), .I1(x19), .I2(x20), .O(n71));
  LUT5 #(.INIT(32'hE81717E8)) lut_n72 (.I0(x9), .I1(x10), .I2(x11), .I3(n68), .I4(n69), .O(n72));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n73 (.I0(x15), .I1(x16), .I2(x17), .I3(n71), .I4(n72), .O(n73));
  LUT3 #(.INIT(8'hE8)) lut_n74 (.I0(n67), .I1(n70), .I2(n73), .O(n74));
  LUT3 #(.INIT(8'hE8)) lut_n75 (.I0(x24), .I1(x25), .I2(x26), .O(n75));
  LUT5 #(.INIT(32'hE81717E8)) lut_n76 (.I0(x15), .I1(x16), .I2(x17), .I3(n71), .I4(n72), .O(n76));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n77 (.I0(x21), .I1(x22), .I2(x23), .I3(n75), .I4(n76), .O(n77));
  LUT3 #(.INIT(8'hE8)) lut_n78 (.I0(x27), .I1(x28), .I2(x29), .O(n78));
  LUT5 #(.INIT(32'hE81717E8)) lut_n79 (.I0(x21), .I1(x22), .I2(x23), .I3(n75), .I4(n76), .O(n79));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n80 (.I0(x30), .I1(x31), .I2(x32), .I3(n78), .I4(n79), .O(n80));
  LUT3 #(.INIT(8'h96)) lut_n81 (.I0(n67), .I1(n70), .I2(n73), .O(n81));
  LUT3 #(.INIT(8'hE8)) lut_n82 (.I0(n77), .I1(n80), .I2(n81), .O(n82));
  LUT3 #(.INIT(8'hE8)) lut_n83 (.I0(x36), .I1(x37), .I2(x38), .O(n83));
  LUT5 #(.INIT(32'hE81717E8)) lut_n84 (.I0(x30), .I1(x31), .I2(x32), .I3(n78), .I4(n79), .O(n84));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n85 (.I0(x33), .I1(x34), .I2(x35), .I3(n83), .I4(n84), .O(n85));
  LUT3 #(.INIT(8'hE8)) lut_n86 (.I0(x42), .I1(x43), .I2(x44), .O(n86));
  LUT5 #(.INIT(32'hE81717E8)) lut_n87 (.I0(x33), .I1(x34), .I2(x35), .I3(n83), .I4(n84), .O(n87));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n88 (.I0(x39), .I1(x40), .I2(x41), .I3(n86), .I4(n87), .O(n88));
  LUT3 #(.INIT(8'h96)) lut_n89 (.I0(n77), .I1(n80), .I2(n81), .O(n89));
  LUT3 #(.INIT(8'hE8)) lut_n90 (.I0(n85), .I1(n88), .I2(n89), .O(n90));
  LUT3 #(.INIT(8'hE8)) lut_n91 (.I0(n74), .I1(n82), .I2(n90), .O(n91));
  LUT3 #(.INIT(8'hE8)) lut_n92 (.I0(x48), .I1(x49), .I2(x50), .O(n92));
  LUT5 #(.INIT(32'hE81717E8)) lut_n93 (.I0(x39), .I1(x40), .I2(x41), .I3(n86), .I4(n87), .O(n93));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n94 (.I0(x45), .I1(x46), .I2(x47), .I3(n92), .I4(n93), .O(n94));
  LUT3 #(.INIT(8'hE8)) lut_n95 (.I0(x54), .I1(x55), .I2(x56), .O(n95));
  LUT5 #(.INIT(32'hE81717E8)) lut_n96 (.I0(x45), .I1(x46), .I2(x47), .I3(n92), .I4(n93), .O(n96));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n97 (.I0(x51), .I1(x52), .I2(x53), .I3(n95), .I4(n96), .O(n97));
  LUT3 #(.INIT(8'h96)) lut_n98 (.I0(n85), .I1(n88), .I2(n89), .O(n98));
  LUT3 #(.INIT(8'hE8)) lut_n99 (.I0(n94), .I1(n97), .I2(n98), .O(n99));
  LUT3 #(.INIT(8'hE8)) lut_n100 (.I0(x60), .I1(x61), .I2(x62), .O(n100));
  LUT5 #(.INIT(32'hE81717E8)) lut_n101 (.I0(x51), .I1(x52), .I2(x53), .I3(n95), .I4(n96), .O(n101));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n102 (.I0(x57), .I1(x58), .I2(x59), .I3(n100), .I4(n101), .O(n102));
  LUT3 #(.INIT(8'h96)) lut_n103 (.I0(x0), .I1(x1), .I2(x2), .O(n103));
  LUT3 #(.INIT(8'h96)) lut_n104 (.I0(x6), .I1(x7), .I2(x8), .O(n104));
  LUT5 #(.INIT(32'hFF969600)) lut_n105 (.I0(x3), .I1(x4), .I2(x5), .I3(n103), .I4(n104), .O(n105));
  LUT3 #(.INIT(8'h96)) lut_n106 (.I0(x12), .I1(x13), .I2(x14), .O(n106));
  LUT5 #(.INIT(32'h96696996)) lut_n107 (.I0(x3), .I1(x4), .I2(x5), .I3(n103), .I4(n104), .O(n107));
  LUT5 #(.INIT(32'hFF969600)) lut_n108 (.I0(x9), .I1(x10), .I2(x11), .I3(n106), .I4(n107), .O(n108));
  LUT5 #(.INIT(32'hE81717E8)) lut_n109 (.I0(x57), .I1(x58), .I2(x59), .I3(n100), .I4(n101), .O(n109));
  LUT3 #(.INIT(8'hE8)) lut_n110 (.I0(n105), .I1(n108), .I2(n109), .O(n110));
  LUT3 #(.INIT(8'h96)) lut_n111 (.I0(n94), .I1(n97), .I2(n98), .O(n111));
  LUT3 #(.INIT(8'hE8)) lut_n112 (.I0(n102), .I1(n110), .I2(n111), .O(n112));
  LUT3 #(.INIT(8'h96)) lut_n113 (.I0(n74), .I1(n82), .I2(n90), .O(n113));
  LUT3 #(.INIT(8'h96)) lut_n114 (.I0(x18), .I1(x19), .I2(x20), .O(n114));
  LUT5 #(.INIT(32'h96696996)) lut_n115 (.I0(x9), .I1(x10), .I2(x11), .I3(n106), .I4(n107), .O(n115));
  LUT5 #(.INIT(32'hFF969600)) lut_n116 (.I0(x15), .I1(x16), .I2(x17), .I3(n114), .I4(n115), .O(n116));
  LUT3 #(.INIT(8'h96)) lut_n117 (.I0(x24), .I1(x25), .I2(x26), .O(n117));
  LUT5 #(.INIT(32'h96696996)) lut_n118 (.I0(x15), .I1(x16), .I2(x17), .I3(n114), .I4(n115), .O(n118));
  LUT5 #(.INIT(32'hFF969600)) lut_n119 (.I0(x21), .I1(x22), .I2(x23), .I3(n117), .I4(n118), .O(n119));
  LUT3 #(.INIT(8'h96)) lut_n120 (.I0(n105), .I1(n108), .I2(n109), .O(n120));
  LUT3 #(.INIT(8'hE8)) lut_n121 (.I0(n116), .I1(n119), .I2(n120), .O(n121));
  LUT3 #(.INIT(8'h96)) lut_n122 (.I0(x27), .I1(x28), .I2(x29), .O(n122));
  LUT5 #(.INIT(32'h96696996)) lut_n123 (.I0(x21), .I1(x22), .I2(x23), .I3(n117), .I4(n118), .O(n123));
  LUT5 #(.INIT(32'hFF969600)) lut_n124 (.I0(x30), .I1(x31), .I2(x32), .I3(n122), .I4(n123), .O(n124));
  LUT3 #(.INIT(8'h96)) lut_n125 (.I0(x36), .I1(x37), .I2(x38), .O(n125));
  LUT5 #(.INIT(32'h96696996)) lut_n126 (.I0(x30), .I1(x31), .I2(x32), .I3(n122), .I4(n123), .O(n126));
  LUT5 #(.INIT(32'hFF969600)) lut_n127 (.I0(x33), .I1(x34), .I2(x35), .I3(n125), .I4(n126), .O(n127));
  LUT3 #(.INIT(8'h96)) lut_n128 (.I0(n116), .I1(n119), .I2(n120), .O(n128));
  LUT3 #(.INIT(8'hE8)) lut_n129 (.I0(n124), .I1(n127), .I2(n128), .O(n129));
  LUT3 #(.INIT(8'h96)) lut_n130 (.I0(n102), .I1(n110), .I2(n111), .O(n130));
  LUT3 #(.INIT(8'hE8)) lut_n131 (.I0(n121), .I1(n129), .I2(n130), .O(n131));
  LUT3 #(.INIT(8'h96)) lut_n132 (.I0(x42), .I1(x43), .I2(x44), .O(n132));
  LUT5 #(.INIT(32'h96696996)) lut_n133 (.I0(x33), .I1(x34), .I2(x35), .I3(n125), .I4(n126), .O(n133));
  LUT5 #(.INIT(32'hFF969600)) lut_n134 (.I0(x39), .I1(x40), .I2(x41), .I3(n132), .I4(n133), .O(n134));
  LUT3 #(.INIT(8'h96)) lut_n135 (.I0(x48), .I1(x49), .I2(x50), .O(n135));
  LUT5 #(.INIT(32'h96696996)) lut_n136 (.I0(x39), .I1(x40), .I2(x41), .I3(n132), .I4(n133), .O(n136));
  LUT5 #(.INIT(32'hFF969600)) lut_n137 (.I0(x45), .I1(x46), .I2(x47), .I3(n135), .I4(n136), .O(n137));
  LUT3 #(.INIT(8'h96)) lut_n138 (.I0(n124), .I1(n127), .I2(n128), .O(n138));
  LUT3 #(.INIT(8'h96)) lut_n139 (.I0(x54), .I1(x55), .I2(x56), .O(n139));
  LUT5 #(.INIT(32'h96696996)) lut_n140 (.I0(x45), .I1(x46), .I2(x47), .I3(n135), .I4(n136), .O(n140));
  LUT5 #(.INIT(32'hFF969600)) lut_n141 (.I0(x51), .I1(x52), .I2(x53), .I3(n139), .I4(n140), .O(n141));
  LUT3 #(.INIT(8'h96)) lut_n142 (.I0(x57), .I1(x58), .I2(x59), .O(n142));
  LUT5 #(.INIT(32'h96696996)) lut_n143 (.I0(x51), .I1(x52), .I2(x53), .I3(n139), .I4(n140), .O(n143));
  LUT5 #(.INIT(32'hFF969600)) lut_n144 (.I0(x60), .I1(x61), .I2(x62), .I3(n142), .I4(n143), .O(n144));
  LUT3 #(.INIT(8'h96)) lut_n145 (.I0(n121), .I1(n129), .I2(n130), .O(n145));
  LUT6 #(.INIT(64'hFFFEFEE8E8808000)) lut_n146 (.I0(n134), .I1(n137), .I2(n138), .I3(n141), .I4(n144), .I5(n145), .O(n146));
  LUT6 #(.INIT(64'hFEEAEAA8EAA8A880)) lut_n147 (.I0(n91), .I1(n99), .I2(n112), .I3(n113), .I4(n131), .I5(n146), .O(n147));
  assign y0 = n147;
endmodule
