module top (x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255, x256, x257, x258, x259, x260, x261, x262, x263, x264, x265, x266, x267, x268, x269, x270, x271, x272, x273, x274, x275, x276, x277, x278, x279, x280, x281, x282, x283, x284, x285, x286, x287, x288, x289, x290, x291, x292, x293, x294, x295, x296, x297, x298, x299, x300, x301, x302, x303, x304, x305, x306, x307, x308, x309, x310, x311, x312, x313, x314, x315, x316, x317, x318, x319, x320, x321, x322, x323, x324, x325, x326, x327, x328, x329, x330, x331, x332, x333, x334, x335, x336, x337, x338, x339, x340, x341, x342, x343, x344, x345, x346, x347, x348, x349, x350, x351, x352, x353, x354, x355, x356, x357, x358, x359, x360, x361, x362, x363, x364, x365, x366, x367, x368, x369, x370, x371, x372, x373, x374, x375, x376, x377, x378, x379, x380, x381, x382, x383, x384, x385, x386, x387, x388, x389, x390, x391, x392, x393, x394, x395, x396, x397, x398, x399, x400, x401, x402, x403, x404, x405, x406, x407, x408, x409, x410, x411, x412, x413, x414, x415, x416, x417, x418, x419, x420, x421, x422, x423, x424, x425, x426, x427, x428, x429, x430, x431, x432, x433, x434, x435, x436, x437, x438, x439, x440, x441, x442, x443, x444, x445, x446, x447, x448, x449, x450, x451, x452, x453, x454, x455, x456, x457, x458, x459, x460, x461, x462, x463, x464, x465, x466, x467, x468, x469, x470, x471, x472, x473, x474, x475, x476, x477, x478, x479, x480, x481, x482, x483, x484, x485, x486, x487, x488, x489, x490, x491, x492, x493, x494, x495, x496, x497, x498, x499, x500, x501, x502, x503, x504, x505, x506, x507, x508, x509, x510, x511, x512, x513, x514, x515, x516, x517, x518, x519, x520, x521, x522, x523, x524, x525, x526, x527, x528, x529, x530, x531, x532, x533, x534, x535, x536, x537, x538, x539, x540, x541, x542, x543, x544, x545, x546, x547, x548, x549, x550, x551, x552, x553, x554, x555, x556, x557, x558, x559, x560, x561, x562, x563, x564, x565, x566, x567, x568, x569, x570, x571, x572, x573, x574, x575, x576, x577, x578, x579, x580, x581, x582, x583, x584, x585, x586, x587, x588, x589, x590, x591, x592, x593, x594, x595, x596, x597, x598, x599, x600, x601, x602, x603, x604, x605, x606, x607, x608, x609, x610, x611, x612, x613, x614, x615, x616, x617, x618, x619, x620, x621, x622, x623, x624, x625, x626, x627, x628, x629, x630, x631, x632, x633, x634, x635, x636, x637, x638, x639, x640, x641, x642, x643, x644, x645, x646, x647, x648, x649, x650, x651, x652, x653, x654, x655, x656, x657, x658, x659, x660, x661, x662, x663, x664, x665, x666, x667, x668, x669, x670, x671, x672, x673, x674, x675, x676, x677, x678, x679, x680, x681, x682, x683, x684, x685, x686, x687, x688, x689, x690, x691, x692, x693, x694, x695, x696, x697, x698, x699, x700, y0);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255, x256, x257, x258, x259, x260, x261, x262, x263, x264, x265, x266, x267, x268, x269, x270, x271, x272, x273, x274, x275, x276, x277, x278, x279, x280, x281, x282, x283, x284, x285, x286, x287, x288, x289, x290, x291, x292, x293, x294, x295, x296, x297, x298, x299, x300, x301, x302, x303, x304, x305, x306, x307, x308, x309, x310, x311, x312, x313, x314, x315, x316, x317, x318, x319, x320, x321, x322, x323, x324, x325, x326, x327, x328, x329, x330, x331, x332, x333, x334, x335, x336, x337, x338, x339, x340, x341, x342, x343, x344, x345, x346, x347, x348, x349, x350, x351, x352, x353, x354, x355, x356, x357, x358, x359, x360, x361, x362, x363, x364, x365, x366, x367, x368, x369, x370, x371, x372, x373, x374, x375, x376, x377, x378, x379, x380, x381, x382, x383, x384, x385, x386, x387, x388, x389, x390, x391, x392, x393, x394, x395, x396, x397, x398, x399, x400, x401, x402, x403, x404, x405, x406, x407, x408, x409, x410, x411, x412, x413, x414, x415, x416, x417, x418, x419, x420, x421, x422, x423, x424, x425, x426, x427, x428, x429, x430, x431, x432, x433, x434, x435, x436, x437, x438, x439, x440, x441, x442, x443, x444, x445, x446, x447, x448, x449, x450, x451, x452, x453, x454, x455, x456, x457, x458, x459, x460, x461, x462, x463, x464, x465, x466, x467, x468, x469, x470, x471, x472, x473, x474, x475, x476, x477, x478, x479, x480, x481, x482, x483, x484, x485, x486, x487, x488, x489, x490, x491, x492, x493, x494, x495, x496, x497, x498, x499, x500, x501, x502, x503, x504, x505, x506, x507, x508, x509, x510, x511, x512, x513, x514, x515, x516, x517, x518, x519, x520, x521, x522, x523, x524, x525, x526, x527, x528, x529, x530, x531, x532, x533, x534, x535, x536, x537, x538, x539, x540, x541, x542, x543, x544, x545, x546, x547, x548, x549, x550, x551, x552, x553, x554, x555, x556, x557, x558, x559, x560, x561, x562, x563, x564, x565, x566, x567, x568, x569, x570, x571, x572, x573, x574, x575, x576, x577, x578, x579, x580, x581, x582, x583, x584, x585, x586, x587, x588, x589, x590, x591, x592, x593, x594, x595, x596, x597, x598, x599, x600, x601, x602, x603, x604, x605, x606, x607, x608, x609, x610, x611, x612, x613, x614, x615, x616, x617, x618, x619, x620, x621, x622, x623, x624, x625, x626, x627, x628, x629, x630, x631, x632, x633, x634, x635, x636, x637, x638, x639, x640, x641, x642, x643, x644, x645, x646, x647, x648, x649, x650, x651, x652, x653, x654, x655, x656, x657, x658, x659, x660, x661, x662, x663, x664, x665, x666, x667, x668, x669, x670, x671, x672, x673, x674, x675, x676, x677, x678, x679, x680, x681, x682, x683, x684, x685, x686, x687, x688, x689, x690, x691, x692, x693, x694, x695, x696, x697, x698, x699, x700;
  output y0;
  wire n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862;
  LUT3 #(.INIT(8'hE8)) lut_n703 (.I0(x0), .I1(x1), .I2(x2), .O(n703));
  LUT3 #(.INIT(8'hE8)) lut_n704 (.I0(x6), .I1(x7), .I2(x8), .O(n704));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n705 (.I0(x3), .I1(x4), .I2(x5), .I3(n703), .I4(n704), .O(n705));
  LUT3 #(.INIT(8'hE8)) lut_n706 (.I0(x12), .I1(x13), .I2(x14), .O(n706));
  LUT5 #(.INIT(32'hE81717E8)) lut_n707 (.I0(x3), .I1(x4), .I2(x5), .I3(n703), .I4(n704), .O(n707));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n708 (.I0(x9), .I1(x10), .I2(x11), .I3(n706), .I4(n707), .O(n708));
  LUT3 #(.INIT(8'hE8)) lut_n709 (.I0(x18), .I1(x19), .I2(x20), .O(n709));
  LUT5 #(.INIT(32'hE81717E8)) lut_n710 (.I0(x9), .I1(x10), .I2(x11), .I3(n706), .I4(n707), .O(n710));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n711 (.I0(x15), .I1(x16), .I2(x17), .I3(n709), .I4(n710), .O(n711));
  LUT3 #(.INIT(8'hE8)) lut_n712 (.I0(n705), .I1(n708), .I2(n711), .O(n712));
  LUT3 #(.INIT(8'hE8)) lut_n713 (.I0(x24), .I1(x25), .I2(x26), .O(n713));
  LUT5 #(.INIT(32'hE81717E8)) lut_n714 (.I0(x15), .I1(x16), .I2(x17), .I3(n709), .I4(n710), .O(n714));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n715 (.I0(x21), .I1(x22), .I2(x23), .I3(n713), .I4(n714), .O(n715));
  LUT3 #(.INIT(8'hE8)) lut_n716 (.I0(x27), .I1(x28), .I2(x29), .O(n716));
  LUT5 #(.INIT(32'hE81717E8)) lut_n717 (.I0(x21), .I1(x22), .I2(x23), .I3(n713), .I4(n714), .O(n717));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n718 (.I0(x30), .I1(x31), .I2(x32), .I3(n716), .I4(n717), .O(n718));
  LUT3 #(.INIT(8'h96)) lut_n719 (.I0(n705), .I1(n708), .I2(n711), .O(n719));
  LUT3 #(.INIT(8'hE8)) lut_n720 (.I0(n715), .I1(n718), .I2(n719), .O(n720));
  LUT3 #(.INIT(8'hE8)) lut_n721 (.I0(x36), .I1(x37), .I2(x38), .O(n721));
  LUT5 #(.INIT(32'hE81717E8)) lut_n722 (.I0(x30), .I1(x31), .I2(x32), .I3(n716), .I4(n717), .O(n722));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n723 (.I0(x33), .I1(x34), .I2(x35), .I3(n721), .I4(n722), .O(n723));
  LUT3 #(.INIT(8'hE8)) lut_n724 (.I0(x42), .I1(x43), .I2(x44), .O(n724));
  LUT5 #(.INIT(32'hE81717E8)) lut_n725 (.I0(x33), .I1(x34), .I2(x35), .I3(n721), .I4(n722), .O(n725));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n726 (.I0(x39), .I1(x40), .I2(x41), .I3(n724), .I4(n725), .O(n726));
  LUT3 #(.INIT(8'h96)) lut_n727 (.I0(n715), .I1(n718), .I2(n719), .O(n727));
  LUT3 #(.INIT(8'hE8)) lut_n728 (.I0(n723), .I1(n726), .I2(n727), .O(n728));
  LUT3 #(.INIT(8'hE8)) lut_n729 (.I0(n712), .I1(n720), .I2(n728), .O(n729));
  LUT3 #(.INIT(8'hE8)) lut_n730 (.I0(x48), .I1(x49), .I2(x50), .O(n730));
  LUT5 #(.INIT(32'hE81717E8)) lut_n731 (.I0(x39), .I1(x40), .I2(x41), .I3(n724), .I4(n725), .O(n731));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n732 (.I0(x45), .I1(x46), .I2(x47), .I3(n730), .I4(n731), .O(n732));
  LUT3 #(.INIT(8'hE8)) lut_n733 (.I0(x54), .I1(x55), .I2(x56), .O(n733));
  LUT5 #(.INIT(32'hE81717E8)) lut_n734 (.I0(x45), .I1(x46), .I2(x47), .I3(n730), .I4(n731), .O(n734));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n735 (.I0(x51), .I1(x52), .I2(x53), .I3(n733), .I4(n734), .O(n735));
  LUT3 #(.INIT(8'h96)) lut_n736 (.I0(n723), .I1(n726), .I2(n727), .O(n736));
  LUT3 #(.INIT(8'hE8)) lut_n737 (.I0(n732), .I1(n735), .I2(n736), .O(n737));
  LUT3 #(.INIT(8'hE8)) lut_n738 (.I0(x60), .I1(x61), .I2(x62), .O(n738));
  LUT5 #(.INIT(32'hE81717E8)) lut_n739 (.I0(x51), .I1(x52), .I2(x53), .I3(n733), .I4(n734), .O(n739));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n740 (.I0(x57), .I1(x58), .I2(x59), .I3(n738), .I4(n739), .O(n740));
  LUT3 #(.INIT(8'hE8)) lut_n741 (.I0(x66), .I1(x67), .I2(x68), .O(n741));
  LUT5 #(.INIT(32'hE81717E8)) lut_n742 (.I0(x57), .I1(x58), .I2(x59), .I3(n738), .I4(n739), .O(n742));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n743 (.I0(x63), .I1(x64), .I2(x65), .I3(n741), .I4(n742), .O(n743));
  LUT3 #(.INIT(8'h96)) lut_n744 (.I0(n732), .I1(n735), .I2(n736), .O(n744));
  LUT3 #(.INIT(8'hE8)) lut_n745 (.I0(n740), .I1(n743), .I2(n744), .O(n745));
  LUT3 #(.INIT(8'h96)) lut_n746 (.I0(n712), .I1(n720), .I2(n728), .O(n746));
  LUT3 #(.INIT(8'hE8)) lut_n747 (.I0(n737), .I1(n745), .I2(n746), .O(n747));
  LUT3 #(.INIT(8'hE8)) lut_n748 (.I0(x72), .I1(x73), .I2(x74), .O(n748));
  LUT5 #(.INIT(32'hE81717E8)) lut_n749 (.I0(x63), .I1(x64), .I2(x65), .I3(n741), .I4(n742), .O(n749));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n750 (.I0(x69), .I1(x70), .I2(x71), .I3(n748), .I4(n749), .O(n750));
  LUT3 #(.INIT(8'hE8)) lut_n751 (.I0(x78), .I1(x79), .I2(x80), .O(n751));
  LUT5 #(.INIT(32'hE81717E8)) lut_n752 (.I0(x69), .I1(x70), .I2(x71), .I3(n748), .I4(n749), .O(n752));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n753 (.I0(x75), .I1(x76), .I2(x77), .I3(n751), .I4(n752), .O(n753));
  LUT3 #(.INIT(8'h96)) lut_n754 (.I0(n740), .I1(n743), .I2(n744), .O(n754));
  LUT3 #(.INIT(8'hE8)) lut_n755 (.I0(n750), .I1(n753), .I2(n754), .O(n755));
  LUT3 #(.INIT(8'hE8)) lut_n756 (.I0(x84), .I1(x85), .I2(x86), .O(n756));
  LUT5 #(.INIT(32'hE81717E8)) lut_n757 (.I0(x75), .I1(x76), .I2(x77), .I3(n751), .I4(n752), .O(n757));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n758 (.I0(x81), .I1(x82), .I2(x83), .I3(n756), .I4(n757), .O(n758));
  LUT3 #(.INIT(8'hE8)) lut_n759 (.I0(x90), .I1(x91), .I2(x92), .O(n759));
  LUT5 #(.INIT(32'hE81717E8)) lut_n760 (.I0(x81), .I1(x82), .I2(x83), .I3(n756), .I4(n757), .O(n760));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n761 (.I0(x87), .I1(x88), .I2(x89), .I3(n759), .I4(n760), .O(n761));
  LUT3 #(.INIT(8'h96)) lut_n762 (.I0(n750), .I1(n753), .I2(n754), .O(n762));
  LUT3 #(.INIT(8'hE8)) lut_n763 (.I0(n758), .I1(n761), .I2(n762), .O(n763));
  LUT3 #(.INIT(8'h96)) lut_n764 (.I0(n737), .I1(n745), .I2(n746), .O(n764));
  LUT3 #(.INIT(8'hE8)) lut_n765 (.I0(n755), .I1(n763), .I2(n764), .O(n765));
  LUT3 #(.INIT(8'hE8)) lut_n766 (.I0(n729), .I1(n747), .I2(n765), .O(n766));
  LUT3 #(.INIT(8'hE8)) lut_n767 (.I0(x96), .I1(x97), .I2(x98), .O(n767));
  LUT5 #(.INIT(32'hE81717E8)) lut_n768 (.I0(x87), .I1(x88), .I2(x89), .I3(n759), .I4(n760), .O(n768));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n769 (.I0(x93), .I1(x94), .I2(x95), .I3(n767), .I4(n768), .O(n769));
  LUT3 #(.INIT(8'hE8)) lut_n770 (.I0(x102), .I1(x103), .I2(x104), .O(n770));
  LUT5 #(.INIT(32'hE81717E8)) lut_n771 (.I0(x93), .I1(x94), .I2(x95), .I3(n767), .I4(n768), .O(n771));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n772 (.I0(x99), .I1(x100), .I2(x101), .I3(n770), .I4(n771), .O(n772));
  LUT3 #(.INIT(8'h96)) lut_n773 (.I0(n758), .I1(n761), .I2(n762), .O(n773));
  LUT3 #(.INIT(8'hE8)) lut_n774 (.I0(n769), .I1(n772), .I2(n773), .O(n774));
  LUT3 #(.INIT(8'hE8)) lut_n775 (.I0(x108), .I1(x109), .I2(x110), .O(n775));
  LUT5 #(.INIT(32'hE81717E8)) lut_n776 (.I0(x99), .I1(x100), .I2(x101), .I3(n770), .I4(n771), .O(n776));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n777 (.I0(x105), .I1(x106), .I2(x107), .I3(n775), .I4(n776), .O(n777));
  LUT3 #(.INIT(8'hE8)) lut_n778 (.I0(x114), .I1(x115), .I2(x116), .O(n778));
  LUT5 #(.INIT(32'hE81717E8)) lut_n779 (.I0(x105), .I1(x106), .I2(x107), .I3(n775), .I4(n776), .O(n779));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n780 (.I0(x111), .I1(x112), .I2(x113), .I3(n778), .I4(n779), .O(n780));
  LUT3 #(.INIT(8'h96)) lut_n781 (.I0(n769), .I1(n772), .I2(n773), .O(n781));
  LUT3 #(.INIT(8'hE8)) lut_n782 (.I0(n777), .I1(n780), .I2(n781), .O(n782));
  LUT3 #(.INIT(8'h96)) lut_n783 (.I0(n755), .I1(n763), .I2(n764), .O(n783));
  LUT3 #(.INIT(8'hE8)) lut_n784 (.I0(n774), .I1(n782), .I2(n783), .O(n784));
  LUT3 #(.INIT(8'hE8)) lut_n785 (.I0(x120), .I1(x121), .I2(x122), .O(n785));
  LUT5 #(.INIT(32'hE81717E8)) lut_n786 (.I0(x111), .I1(x112), .I2(x113), .I3(n778), .I4(n779), .O(n786));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n787 (.I0(x117), .I1(x118), .I2(x119), .I3(n785), .I4(n786), .O(n787));
  LUT3 #(.INIT(8'hE8)) lut_n788 (.I0(x126), .I1(x127), .I2(x128), .O(n788));
  LUT5 #(.INIT(32'hE81717E8)) lut_n789 (.I0(x117), .I1(x118), .I2(x119), .I3(n785), .I4(n786), .O(n789));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n790 (.I0(x123), .I1(x124), .I2(x125), .I3(n788), .I4(n789), .O(n790));
  LUT3 #(.INIT(8'h96)) lut_n791 (.I0(n777), .I1(n780), .I2(n781), .O(n791));
  LUT3 #(.INIT(8'hE8)) lut_n792 (.I0(n787), .I1(n790), .I2(n791), .O(n792));
  LUT3 #(.INIT(8'hE8)) lut_n793 (.I0(x132), .I1(x133), .I2(x134), .O(n793));
  LUT5 #(.INIT(32'hE81717E8)) lut_n794 (.I0(x123), .I1(x124), .I2(x125), .I3(n788), .I4(n789), .O(n794));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n795 (.I0(x129), .I1(x130), .I2(x131), .I3(n793), .I4(n794), .O(n795));
  LUT3 #(.INIT(8'hE8)) lut_n796 (.I0(x138), .I1(x139), .I2(x140), .O(n796));
  LUT5 #(.INIT(32'hE81717E8)) lut_n797 (.I0(x129), .I1(x130), .I2(x131), .I3(n793), .I4(n794), .O(n797));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n798 (.I0(x135), .I1(x136), .I2(x137), .I3(n796), .I4(n797), .O(n798));
  LUT3 #(.INIT(8'h96)) lut_n799 (.I0(n787), .I1(n790), .I2(n791), .O(n799));
  LUT3 #(.INIT(8'hE8)) lut_n800 (.I0(n795), .I1(n798), .I2(n799), .O(n800));
  LUT3 #(.INIT(8'h96)) lut_n801 (.I0(n774), .I1(n782), .I2(n783), .O(n801));
  LUT3 #(.INIT(8'hE8)) lut_n802 (.I0(n792), .I1(n800), .I2(n801), .O(n802));
  LUT3 #(.INIT(8'h96)) lut_n803 (.I0(n729), .I1(n747), .I2(n765), .O(n803));
  LUT3 #(.INIT(8'hE8)) lut_n804 (.I0(n784), .I1(n802), .I2(n803), .O(n804));
  LUT3 #(.INIT(8'hE8)) lut_n805 (.I0(x144), .I1(x145), .I2(x146), .O(n805));
  LUT5 #(.INIT(32'hE81717E8)) lut_n806 (.I0(x135), .I1(x136), .I2(x137), .I3(n796), .I4(n797), .O(n806));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n807 (.I0(x141), .I1(x142), .I2(x143), .I3(n805), .I4(n806), .O(n807));
  LUT3 #(.INIT(8'hE8)) lut_n808 (.I0(x150), .I1(x151), .I2(x152), .O(n808));
  LUT5 #(.INIT(32'hE81717E8)) lut_n809 (.I0(x141), .I1(x142), .I2(x143), .I3(n805), .I4(n806), .O(n809));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n810 (.I0(x147), .I1(x148), .I2(x149), .I3(n808), .I4(n809), .O(n810));
  LUT3 #(.INIT(8'h96)) lut_n811 (.I0(n795), .I1(n798), .I2(n799), .O(n811));
  LUT3 #(.INIT(8'hE8)) lut_n812 (.I0(n807), .I1(n810), .I2(n811), .O(n812));
  LUT3 #(.INIT(8'hE8)) lut_n813 (.I0(x156), .I1(x157), .I2(x158), .O(n813));
  LUT5 #(.INIT(32'hE81717E8)) lut_n814 (.I0(x147), .I1(x148), .I2(x149), .I3(n808), .I4(n809), .O(n814));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n815 (.I0(x153), .I1(x154), .I2(x155), .I3(n813), .I4(n814), .O(n815));
  LUT3 #(.INIT(8'hE8)) lut_n816 (.I0(x162), .I1(x163), .I2(x164), .O(n816));
  LUT5 #(.INIT(32'hE81717E8)) lut_n817 (.I0(x153), .I1(x154), .I2(x155), .I3(n813), .I4(n814), .O(n817));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n818 (.I0(x159), .I1(x160), .I2(x161), .I3(n816), .I4(n817), .O(n818));
  LUT3 #(.INIT(8'h96)) lut_n819 (.I0(n807), .I1(n810), .I2(n811), .O(n819));
  LUT3 #(.INIT(8'hE8)) lut_n820 (.I0(n815), .I1(n818), .I2(n819), .O(n820));
  LUT3 #(.INIT(8'h96)) lut_n821 (.I0(n792), .I1(n800), .I2(n801), .O(n821));
  LUT3 #(.INIT(8'hE8)) lut_n822 (.I0(n812), .I1(n820), .I2(n821), .O(n822));
  LUT3 #(.INIT(8'hE8)) lut_n823 (.I0(x168), .I1(x169), .I2(x170), .O(n823));
  LUT5 #(.INIT(32'hE81717E8)) lut_n824 (.I0(x159), .I1(x160), .I2(x161), .I3(n816), .I4(n817), .O(n824));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n825 (.I0(x165), .I1(x166), .I2(x167), .I3(n823), .I4(n824), .O(n825));
  LUT3 #(.INIT(8'hE8)) lut_n826 (.I0(x174), .I1(x175), .I2(x176), .O(n826));
  LUT5 #(.INIT(32'hE81717E8)) lut_n827 (.I0(x165), .I1(x166), .I2(x167), .I3(n823), .I4(n824), .O(n827));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n828 (.I0(x171), .I1(x172), .I2(x173), .I3(n826), .I4(n827), .O(n828));
  LUT3 #(.INIT(8'h96)) lut_n829 (.I0(n815), .I1(n818), .I2(n819), .O(n829));
  LUT3 #(.INIT(8'hE8)) lut_n830 (.I0(n825), .I1(n828), .I2(n829), .O(n830));
  LUT3 #(.INIT(8'hE8)) lut_n831 (.I0(x180), .I1(x181), .I2(x182), .O(n831));
  LUT5 #(.INIT(32'hE81717E8)) lut_n832 (.I0(x171), .I1(x172), .I2(x173), .I3(n826), .I4(n827), .O(n832));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n833 (.I0(x177), .I1(x178), .I2(x179), .I3(n831), .I4(n832), .O(n833));
  LUT3 #(.INIT(8'hE8)) lut_n834 (.I0(x186), .I1(x187), .I2(x188), .O(n834));
  LUT5 #(.INIT(32'hE81717E8)) lut_n835 (.I0(x177), .I1(x178), .I2(x179), .I3(n831), .I4(n832), .O(n835));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n836 (.I0(x183), .I1(x184), .I2(x185), .I3(n834), .I4(n835), .O(n836));
  LUT3 #(.INIT(8'h96)) lut_n837 (.I0(n825), .I1(n828), .I2(n829), .O(n837));
  LUT3 #(.INIT(8'hE8)) lut_n838 (.I0(n833), .I1(n836), .I2(n837), .O(n838));
  LUT3 #(.INIT(8'h96)) lut_n839 (.I0(n812), .I1(n820), .I2(n821), .O(n839));
  LUT3 #(.INIT(8'hE8)) lut_n840 (.I0(n830), .I1(n838), .I2(n839), .O(n840));
  LUT3 #(.INIT(8'h96)) lut_n841 (.I0(n784), .I1(n802), .I2(n803), .O(n841));
  LUT3 #(.INIT(8'hE8)) lut_n842 (.I0(n822), .I1(n840), .I2(n841), .O(n842));
  LUT3 #(.INIT(8'hE8)) lut_n843 (.I0(n766), .I1(n804), .I2(n842), .O(n843));
  LUT3 #(.INIT(8'hE8)) lut_n844 (.I0(x192), .I1(x193), .I2(x194), .O(n844));
  LUT5 #(.INIT(32'hE81717E8)) lut_n845 (.I0(x183), .I1(x184), .I2(x185), .I3(n834), .I4(n835), .O(n845));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n846 (.I0(x189), .I1(x190), .I2(x191), .I3(n844), .I4(n845), .O(n846));
  LUT3 #(.INIT(8'hE8)) lut_n847 (.I0(x198), .I1(x199), .I2(x200), .O(n847));
  LUT5 #(.INIT(32'hE81717E8)) lut_n848 (.I0(x189), .I1(x190), .I2(x191), .I3(n844), .I4(n845), .O(n848));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n849 (.I0(x195), .I1(x196), .I2(x197), .I3(n847), .I4(n848), .O(n849));
  LUT3 #(.INIT(8'h96)) lut_n850 (.I0(n833), .I1(n836), .I2(n837), .O(n850));
  LUT3 #(.INIT(8'hE8)) lut_n851 (.I0(n846), .I1(n849), .I2(n850), .O(n851));
  LUT3 #(.INIT(8'hE8)) lut_n852 (.I0(x204), .I1(x205), .I2(x206), .O(n852));
  LUT5 #(.INIT(32'hE81717E8)) lut_n853 (.I0(x195), .I1(x196), .I2(x197), .I3(n847), .I4(n848), .O(n853));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n854 (.I0(x201), .I1(x202), .I2(x203), .I3(n852), .I4(n853), .O(n854));
  LUT3 #(.INIT(8'hE8)) lut_n855 (.I0(x210), .I1(x211), .I2(x212), .O(n855));
  LUT5 #(.INIT(32'hE81717E8)) lut_n856 (.I0(x201), .I1(x202), .I2(x203), .I3(n852), .I4(n853), .O(n856));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n857 (.I0(x207), .I1(x208), .I2(x209), .I3(n855), .I4(n856), .O(n857));
  LUT3 #(.INIT(8'h96)) lut_n858 (.I0(n846), .I1(n849), .I2(n850), .O(n858));
  LUT3 #(.INIT(8'hE8)) lut_n859 (.I0(n854), .I1(n857), .I2(n858), .O(n859));
  LUT3 #(.INIT(8'h96)) lut_n860 (.I0(n830), .I1(n838), .I2(n839), .O(n860));
  LUT3 #(.INIT(8'hE8)) lut_n861 (.I0(n851), .I1(n859), .I2(n860), .O(n861));
  LUT3 #(.INIT(8'hE8)) lut_n862 (.I0(x216), .I1(x217), .I2(x218), .O(n862));
  LUT5 #(.INIT(32'hE81717E8)) lut_n863 (.I0(x207), .I1(x208), .I2(x209), .I3(n855), .I4(n856), .O(n863));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n864 (.I0(x213), .I1(x214), .I2(x215), .I3(n862), .I4(n863), .O(n864));
  LUT3 #(.INIT(8'hE8)) lut_n865 (.I0(x222), .I1(x223), .I2(x224), .O(n865));
  LUT5 #(.INIT(32'hE81717E8)) lut_n866 (.I0(x213), .I1(x214), .I2(x215), .I3(n862), .I4(n863), .O(n866));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n867 (.I0(x219), .I1(x220), .I2(x221), .I3(n865), .I4(n866), .O(n867));
  LUT3 #(.INIT(8'h96)) lut_n868 (.I0(n854), .I1(n857), .I2(n858), .O(n868));
  LUT3 #(.INIT(8'hE8)) lut_n869 (.I0(n864), .I1(n867), .I2(n868), .O(n869));
  LUT3 #(.INIT(8'hE8)) lut_n870 (.I0(x228), .I1(x229), .I2(x230), .O(n870));
  LUT5 #(.INIT(32'hE81717E8)) lut_n871 (.I0(x219), .I1(x220), .I2(x221), .I3(n865), .I4(n866), .O(n871));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n872 (.I0(x225), .I1(x226), .I2(x227), .I3(n870), .I4(n871), .O(n872));
  LUT3 #(.INIT(8'hE8)) lut_n873 (.I0(x234), .I1(x235), .I2(x236), .O(n873));
  LUT5 #(.INIT(32'hE81717E8)) lut_n874 (.I0(x225), .I1(x226), .I2(x227), .I3(n870), .I4(n871), .O(n874));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n875 (.I0(x231), .I1(x232), .I2(x233), .I3(n873), .I4(n874), .O(n875));
  LUT3 #(.INIT(8'h96)) lut_n876 (.I0(n864), .I1(n867), .I2(n868), .O(n876));
  LUT3 #(.INIT(8'hE8)) lut_n877 (.I0(n872), .I1(n875), .I2(n876), .O(n877));
  LUT3 #(.INIT(8'h96)) lut_n878 (.I0(n851), .I1(n859), .I2(n860), .O(n878));
  LUT3 #(.INIT(8'hE8)) lut_n879 (.I0(n869), .I1(n877), .I2(n878), .O(n879));
  LUT3 #(.INIT(8'h96)) lut_n880 (.I0(n822), .I1(n840), .I2(n841), .O(n880));
  LUT3 #(.INIT(8'hE8)) lut_n881 (.I0(n861), .I1(n879), .I2(n880), .O(n881));
  LUT3 #(.INIT(8'hE8)) lut_n882 (.I0(x240), .I1(x241), .I2(x242), .O(n882));
  LUT5 #(.INIT(32'hE81717E8)) lut_n883 (.I0(x231), .I1(x232), .I2(x233), .I3(n873), .I4(n874), .O(n883));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n884 (.I0(x237), .I1(x238), .I2(x239), .I3(n882), .I4(n883), .O(n884));
  LUT3 #(.INIT(8'hE8)) lut_n885 (.I0(x246), .I1(x247), .I2(x248), .O(n885));
  LUT5 #(.INIT(32'hE81717E8)) lut_n886 (.I0(x237), .I1(x238), .I2(x239), .I3(n882), .I4(n883), .O(n886));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n887 (.I0(x243), .I1(x244), .I2(x245), .I3(n885), .I4(n886), .O(n887));
  LUT3 #(.INIT(8'h96)) lut_n888 (.I0(n872), .I1(n875), .I2(n876), .O(n888));
  LUT3 #(.INIT(8'hE8)) lut_n889 (.I0(n884), .I1(n887), .I2(n888), .O(n889));
  LUT3 #(.INIT(8'hE8)) lut_n890 (.I0(x252), .I1(x253), .I2(x254), .O(n890));
  LUT5 #(.INIT(32'hE81717E8)) lut_n891 (.I0(x243), .I1(x244), .I2(x245), .I3(n885), .I4(n886), .O(n891));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n892 (.I0(x249), .I1(x250), .I2(x251), .I3(n890), .I4(n891), .O(n892));
  LUT3 #(.INIT(8'hE8)) lut_n893 (.I0(x258), .I1(x259), .I2(x260), .O(n893));
  LUT5 #(.INIT(32'hE81717E8)) lut_n894 (.I0(x249), .I1(x250), .I2(x251), .I3(n890), .I4(n891), .O(n894));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n895 (.I0(x255), .I1(x256), .I2(x257), .I3(n893), .I4(n894), .O(n895));
  LUT3 #(.INIT(8'h96)) lut_n896 (.I0(n884), .I1(n887), .I2(n888), .O(n896));
  LUT3 #(.INIT(8'hE8)) lut_n897 (.I0(n892), .I1(n895), .I2(n896), .O(n897));
  LUT3 #(.INIT(8'h96)) lut_n898 (.I0(n869), .I1(n877), .I2(n878), .O(n898));
  LUT3 #(.INIT(8'hE8)) lut_n899 (.I0(n889), .I1(n897), .I2(n898), .O(n899));
  LUT3 #(.INIT(8'hE8)) lut_n900 (.I0(x264), .I1(x265), .I2(x266), .O(n900));
  LUT5 #(.INIT(32'hE81717E8)) lut_n901 (.I0(x255), .I1(x256), .I2(x257), .I3(n893), .I4(n894), .O(n901));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n902 (.I0(x261), .I1(x262), .I2(x263), .I3(n900), .I4(n901), .O(n902));
  LUT3 #(.INIT(8'hE8)) lut_n903 (.I0(x270), .I1(x271), .I2(x272), .O(n903));
  LUT5 #(.INIT(32'hE81717E8)) lut_n904 (.I0(x261), .I1(x262), .I2(x263), .I3(n900), .I4(n901), .O(n904));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n905 (.I0(x267), .I1(x268), .I2(x269), .I3(n903), .I4(n904), .O(n905));
  LUT3 #(.INIT(8'h96)) lut_n906 (.I0(n892), .I1(n895), .I2(n896), .O(n906));
  LUT3 #(.INIT(8'hE8)) lut_n907 (.I0(n902), .I1(n905), .I2(n906), .O(n907));
  LUT3 #(.INIT(8'hE8)) lut_n908 (.I0(x276), .I1(x277), .I2(x278), .O(n908));
  LUT5 #(.INIT(32'hE81717E8)) lut_n909 (.I0(x267), .I1(x268), .I2(x269), .I3(n903), .I4(n904), .O(n909));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n910 (.I0(x273), .I1(x274), .I2(x275), .I3(n908), .I4(n909), .O(n910));
  LUT3 #(.INIT(8'hE8)) lut_n911 (.I0(x282), .I1(x283), .I2(x284), .O(n911));
  LUT5 #(.INIT(32'hE81717E8)) lut_n912 (.I0(x273), .I1(x274), .I2(x275), .I3(n908), .I4(n909), .O(n912));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n913 (.I0(x279), .I1(x280), .I2(x281), .I3(n911), .I4(n912), .O(n913));
  LUT3 #(.INIT(8'h96)) lut_n914 (.I0(n902), .I1(n905), .I2(n906), .O(n914));
  LUT3 #(.INIT(8'hE8)) lut_n915 (.I0(n910), .I1(n913), .I2(n914), .O(n915));
  LUT3 #(.INIT(8'h96)) lut_n916 (.I0(n889), .I1(n897), .I2(n898), .O(n916));
  LUT3 #(.INIT(8'hE8)) lut_n917 (.I0(n907), .I1(n915), .I2(n916), .O(n917));
  LUT3 #(.INIT(8'h96)) lut_n918 (.I0(n861), .I1(n879), .I2(n880), .O(n918));
  LUT3 #(.INIT(8'hE8)) lut_n919 (.I0(n899), .I1(n917), .I2(n918), .O(n919));
  LUT3 #(.INIT(8'h96)) lut_n920 (.I0(n766), .I1(n804), .I2(n842), .O(n920));
  LUT3 #(.INIT(8'hE8)) lut_n921 (.I0(n881), .I1(n919), .I2(n920), .O(n921));
  LUT3 #(.INIT(8'hE8)) lut_n922 (.I0(x288), .I1(x289), .I2(x290), .O(n922));
  LUT5 #(.INIT(32'hE81717E8)) lut_n923 (.I0(x279), .I1(x280), .I2(x281), .I3(n911), .I4(n912), .O(n923));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n924 (.I0(x285), .I1(x286), .I2(x287), .I3(n922), .I4(n923), .O(n924));
  LUT3 #(.INIT(8'hE8)) lut_n925 (.I0(x294), .I1(x295), .I2(x296), .O(n925));
  LUT5 #(.INIT(32'hE81717E8)) lut_n926 (.I0(x285), .I1(x286), .I2(x287), .I3(n922), .I4(n923), .O(n926));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n927 (.I0(x291), .I1(x292), .I2(x293), .I3(n925), .I4(n926), .O(n927));
  LUT3 #(.INIT(8'h96)) lut_n928 (.I0(n910), .I1(n913), .I2(n914), .O(n928));
  LUT3 #(.INIT(8'hE8)) lut_n929 (.I0(n924), .I1(n927), .I2(n928), .O(n929));
  LUT3 #(.INIT(8'hE8)) lut_n930 (.I0(x297), .I1(x298), .I2(x299), .O(n930));
  LUT5 #(.INIT(32'hE81717E8)) lut_n931 (.I0(x291), .I1(x292), .I2(x293), .I3(n925), .I4(n926), .O(n931));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n932 (.I0(x300), .I1(x301), .I2(x302), .I3(n930), .I4(n931), .O(n932));
  LUT3 #(.INIT(8'hE8)) lut_n933 (.I0(x306), .I1(x307), .I2(x308), .O(n933));
  LUT5 #(.INIT(32'hE81717E8)) lut_n934 (.I0(x300), .I1(x301), .I2(x302), .I3(n930), .I4(n931), .O(n934));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n935 (.I0(x303), .I1(x304), .I2(x305), .I3(n933), .I4(n934), .O(n935));
  LUT3 #(.INIT(8'h96)) lut_n936 (.I0(n924), .I1(n927), .I2(n928), .O(n936));
  LUT3 #(.INIT(8'hE8)) lut_n937 (.I0(n932), .I1(n935), .I2(n936), .O(n937));
  LUT3 #(.INIT(8'h96)) lut_n938 (.I0(n907), .I1(n915), .I2(n916), .O(n938));
  LUT3 #(.INIT(8'hE8)) lut_n939 (.I0(n929), .I1(n937), .I2(n938), .O(n939));
  LUT3 #(.INIT(8'hE8)) lut_n940 (.I0(x312), .I1(x313), .I2(x314), .O(n940));
  LUT5 #(.INIT(32'hE81717E8)) lut_n941 (.I0(x303), .I1(x304), .I2(x305), .I3(n933), .I4(n934), .O(n941));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n942 (.I0(x309), .I1(x310), .I2(x311), .I3(n940), .I4(n941), .O(n942));
  LUT3 #(.INIT(8'hE8)) lut_n943 (.I0(x318), .I1(x319), .I2(x320), .O(n943));
  LUT5 #(.INIT(32'hE81717E8)) lut_n944 (.I0(x309), .I1(x310), .I2(x311), .I3(n940), .I4(n941), .O(n944));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n945 (.I0(x315), .I1(x316), .I2(x317), .I3(n943), .I4(n944), .O(n945));
  LUT3 #(.INIT(8'h96)) lut_n946 (.I0(n932), .I1(n935), .I2(n936), .O(n946));
  LUT3 #(.INIT(8'hE8)) lut_n947 (.I0(n942), .I1(n945), .I2(n946), .O(n947));
  LUT3 #(.INIT(8'hE8)) lut_n948 (.I0(x324), .I1(x325), .I2(x326), .O(n948));
  LUT5 #(.INIT(32'hE81717E8)) lut_n949 (.I0(x315), .I1(x316), .I2(x317), .I3(n943), .I4(n944), .O(n949));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n950 (.I0(x321), .I1(x322), .I2(x323), .I3(n948), .I4(n949), .O(n950));
  LUT3 #(.INIT(8'hE8)) lut_n951 (.I0(x330), .I1(x331), .I2(x332), .O(n951));
  LUT5 #(.INIT(32'hE81717E8)) lut_n952 (.I0(x321), .I1(x322), .I2(x323), .I3(n948), .I4(n949), .O(n952));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n953 (.I0(x327), .I1(x328), .I2(x329), .I3(n951), .I4(n952), .O(n953));
  LUT3 #(.INIT(8'h96)) lut_n954 (.I0(n942), .I1(n945), .I2(n946), .O(n954));
  LUT3 #(.INIT(8'hE8)) lut_n955 (.I0(n950), .I1(n953), .I2(n954), .O(n955));
  LUT3 #(.INIT(8'h96)) lut_n956 (.I0(n929), .I1(n937), .I2(n938), .O(n956));
  LUT3 #(.INIT(8'hE8)) lut_n957 (.I0(n947), .I1(n955), .I2(n956), .O(n957));
  LUT3 #(.INIT(8'h96)) lut_n958 (.I0(n899), .I1(n917), .I2(n918), .O(n958));
  LUT3 #(.INIT(8'hE8)) lut_n959 (.I0(n939), .I1(n957), .I2(n958), .O(n959));
  LUT3 #(.INIT(8'hE8)) lut_n960 (.I0(x336), .I1(x337), .I2(x338), .O(n960));
  LUT5 #(.INIT(32'hE81717E8)) lut_n961 (.I0(x327), .I1(x328), .I2(x329), .I3(n951), .I4(n952), .O(n961));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n962 (.I0(x333), .I1(x334), .I2(x335), .I3(n960), .I4(n961), .O(n962));
  LUT3 #(.INIT(8'hE8)) lut_n963 (.I0(x342), .I1(x343), .I2(x344), .O(n963));
  LUT5 #(.INIT(32'hE81717E8)) lut_n964 (.I0(x333), .I1(x334), .I2(x335), .I3(n960), .I4(n961), .O(n964));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n965 (.I0(x339), .I1(x340), .I2(x341), .I3(n963), .I4(n964), .O(n965));
  LUT3 #(.INIT(8'h96)) lut_n966 (.I0(n950), .I1(n953), .I2(n954), .O(n966));
  LUT3 #(.INIT(8'hE8)) lut_n967 (.I0(n962), .I1(n965), .I2(n966), .O(n967));
  LUT3 #(.INIT(8'hE8)) lut_n968 (.I0(x348), .I1(x349), .I2(x350), .O(n968));
  LUT5 #(.INIT(32'hE81717E8)) lut_n969 (.I0(x339), .I1(x340), .I2(x341), .I3(n963), .I4(n964), .O(n969));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n970 (.I0(x345), .I1(x346), .I2(x347), .I3(n968), .I4(n969), .O(n970));
  LUT3 #(.INIT(8'hE8)) lut_n971 (.I0(x354), .I1(x355), .I2(x356), .O(n971));
  LUT5 #(.INIT(32'hE81717E8)) lut_n972 (.I0(x345), .I1(x346), .I2(x347), .I3(n968), .I4(n969), .O(n972));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n973 (.I0(x351), .I1(x352), .I2(x353), .I3(n971), .I4(n972), .O(n973));
  LUT3 #(.INIT(8'h96)) lut_n974 (.I0(n962), .I1(n965), .I2(n966), .O(n974));
  LUT3 #(.INIT(8'hE8)) lut_n975 (.I0(n970), .I1(n973), .I2(n974), .O(n975));
  LUT3 #(.INIT(8'h96)) lut_n976 (.I0(n947), .I1(n955), .I2(n956), .O(n976));
  LUT3 #(.INIT(8'hE8)) lut_n977 (.I0(n967), .I1(n975), .I2(n976), .O(n977));
  LUT3 #(.INIT(8'hE8)) lut_n978 (.I0(x360), .I1(x361), .I2(x362), .O(n978));
  LUT5 #(.INIT(32'hE81717E8)) lut_n979 (.I0(x351), .I1(x352), .I2(x353), .I3(n971), .I4(n972), .O(n979));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n980 (.I0(x357), .I1(x358), .I2(x359), .I3(n978), .I4(n979), .O(n980));
  LUT3 #(.INIT(8'hE8)) lut_n981 (.I0(x366), .I1(x367), .I2(x368), .O(n981));
  LUT5 #(.INIT(32'hE81717E8)) lut_n982 (.I0(x357), .I1(x358), .I2(x359), .I3(n978), .I4(n979), .O(n982));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n983 (.I0(x363), .I1(x364), .I2(x365), .I3(n981), .I4(n982), .O(n983));
  LUT3 #(.INIT(8'h96)) lut_n984 (.I0(n970), .I1(n973), .I2(n974), .O(n984));
  LUT3 #(.INIT(8'hE8)) lut_n985 (.I0(n980), .I1(n983), .I2(n984), .O(n985));
  LUT3 #(.INIT(8'hE8)) lut_n986 (.I0(x372), .I1(x373), .I2(x374), .O(n986));
  LUT5 #(.INIT(32'hE81717E8)) lut_n987 (.I0(x363), .I1(x364), .I2(x365), .I3(n981), .I4(n982), .O(n987));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n988 (.I0(x369), .I1(x370), .I2(x371), .I3(n986), .I4(n987), .O(n988));
  LUT3 #(.INIT(8'hE8)) lut_n989 (.I0(x378), .I1(x379), .I2(x380), .O(n989));
  LUT5 #(.INIT(32'hE81717E8)) lut_n990 (.I0(x369), .I1(x370), .I2(x371), .I3(n986), .I4(n987), .O(n990));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n991 (.I0(x375), .I1(x376), .I2(x377), .I3(n989), .I4(n990), .O(n991));
  LUT3 #(.INIT(8'h96)) lut_n992 (.I0(n980), .I1(n983), .I2(n984), .O(n992));
  LUT3 #(.INIT(8'hE8)) lut_n993 (.I0(n988), .I1(n991), .I2(n992), .O(n993));
  LUT3 #(.INIT(8'h96)) lut_n994 (.I0(n967), .I1(n975), .I2(n976), .O(n994));
  LUT3 #(.INIT(8'hE8)) lut_n995 (.I0(n985), .I1(n993), .I2(n994), .O(n995));
  LUT3 #(.INIT(8'h96)) lut_n996 (.I0(n939), .I1(n957), .I2(n958), .O(n996));
  LUT3 #(.INIT(8'hE8)) lut_n997 (.I0(n977), .I1(n995), .I2(n996), .O(n997));
  LUT3 #(.INIT(8'h96)) lut_n998 (.I0(n881), .I1(n919), .I2(n920), .O(n998));
  LUT3 #(.INIT(8'hE8)) lut_n999 (.I0(n959), .I1(n997), .I2(n998), .O(n999));
  LUT3 #(.INIT(8'hE8)) lut_n1000 (.I0(n843), .I1(n921), .I2(n999), .O(n1000));
  LUT3 #(.INIT(8'hE8)) lut_n1001 (.I0(x384), .I1(x385), .I2(x386), .O(n1001));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1002 (.I0(x375), .I1(x376), .I2(x377), .I3(n989), .I4(n990), .O(n1002));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1003 (.I0(x381), .I1(x382), .I2(x383), .I3(n1001), .I4(n1002), .O(n1003));
  LUT3 #(.INIT(8'hE8)) lut_n1004 (.I0(x390), .I1(x391), .I2(x392), .O(n1004));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1005 (.I0(x381), .I1(x382), .I2(x383), .I3(n1001), .I4(n1002), .O(n1005));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1006 (.I0(x387), .I1(x388), .I2(x389), .I3(n1004), .I4(n1005), .O(n1006));
  LUT3 #(.INIT(8'h96)) lut_n1007 (.I0(n988), .I1(n991), .I2(n992), .O(n1007));
  LUT3 #(.INIT(8'hE8)) lut_n1008 (.I0(n1003), .I1(n1006), .I2(n1007), .O(n1008));
  LUT3 #(.INIT(8'hE8)) lut_n1009 (.I0(x396), .I1(x397), .I2(x398), .O(n1009));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1010 (.I0(x387), .I1(x388), .I2(x389), .I3(n1004), .I4(n1005), .O(n1010));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1011 (.I0(x393), .I1(x394), .I2(x395), .I3(n1009), .I4(n1010), .O(n1011));
  LUT3 #(.INIT(8'hE8)) lut_n1012 (.I0(x402), .I1(x403), .I2(x404), .O(n1012));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1013 (.I0(x393), .I1(x394), .I2(x395), .I3(n1009), .I4(n1010), .O(n1013));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1014 (.I0(x399), .I1(x400), .I2(x401), .I3(n1012), .I4(n1013), .O(n1014));
  LUT3 #(.INIT(8'h96)) lut_n1015 (.I0(n1003), .I1(n1006), .I2(n1007), .O(n1015));
  LUT3 #(.INIT(8'hE8)) lut_n1016 (.I0(n1011), .I1(n1014), .I2(n1015), .O(n1016));
  LUT3 #(.INIT(8'h96)) lut_n1017 (.I0(n985), .I1(n993), .I2(n994), .O(n1017));
  LUT3 #(.INIT(8'hE8)) lut_n1018 (.I0(n1008), .I1(n1016), .I2(n1017), .O(n1018));
  LUT3 #(.INIT(8'hE8)) lut_n1019 (.I0(x408), .I1(x409), .I2(x410), .O(n1019));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1020 (.I0(x399), .I1(x400), .I2(x401), .I3(n1012), .I4(n1013), .O(n1020));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1021 (.I0(x405), .I1(x406), .I2(x407), .I3(n1019), .I4(n1020), .O(n1021));
  LUT3 #(.INIT(8'hE8)) lut_n1022 (.I0(x414), .I1(x415), .I2(x416), .O(n1022));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1023 (.I0(x405), .I1(x406), .I2(x407), .I3(n1019), .I4(n1020), .O(n1023));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1024 (.I0(x411), .I1(x412), .I2(x413), .I3(n1022), .I4(n1023), .O(n1024));
  LUT3 #(.INIT(8'h96)) lut_n1025 (.I0(n1011), .I1(n1014), .I2(n1015), .O(n1025));
  LUT3 #(.INIT(8'hE8)) lut_n1026 (.I0(n1021), .I1(n1024), .I2(n1025), .O(n1026));
  LUT3 #(.INIT(8'hE8)) lut_n1027 (.I0(x420), .I1(x421), .I2(x422), .O(n1027));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1028 (.I0(x411), .I1(x412), .I2(x413), .I3(n1022), .I4(n1023), .O(n1028));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1029 (.I0(x417), .I1(x418), .I2(x419), .I3(n1027), .I4(n1028), .O(n1029));
  LUT3 #(.INIT(8'hE8)) lut_n1030 (.I0(x426), .I1(x427), .I2(x428), .O(n1030));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1031 (.I0(x417), .I1(x418), .I2(x419), .I3(n1027), .I4(n1028), .O(n1031));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1032 (.I0(x423), .I1(x424), .I2(x425), .I3(n1030), .I4(n1031), .O(n1032));
  LUT3 #(.INIT(8'h96)) lut_n1033 (.I0(n1021), .I1(n1024), .I2(n1025), .O(n1033));
  LUT3 #(.INIT(8'hE8)) lut_n1034 (.I0(n1029), .I1(n1032), .I2(n1033), .O(n1034));
  LUT3 #(.INIT(8'h96)) lut_n1035 (.I0(n1008), .I1(n1016), .I2(n1017), .O(n1035));
  LUT3 #(.INIT(8'hE8)) lut_n1036 (.I0(n1026), .I1(n1034), .I2(n1035), .O(n1036));
  LUT3 #(.INIT(8'h96)) lut_n1037 (.I0(n977), .I1(n995), .I2(n996), .O(n1037));
  LUT3 #(.INIT(8'hE8)) lut_n1038 (.I0(n1018), .I1(n1036), .I2(n1037), .O(n1038));
  LUT3 #(.INIT(8'hE8)) lut_n1039 (.I0(x432), .I1(x433), .I2(x434), .O(n1039));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1040 (.I0(x423), .I1(x424), .I2(x425), .I3(n1030), .I4(n1031), .O(n1040));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1041 (.I0(x429), .I1(x430), .I2(x431), .I3(n1039), .I4(n1040), .O(n1041));
  LUT3 #(.INIT(8'hE8)) lut_n1042 (.I0(x438), .I1(x439), .I2(x440), .O(n1042));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1043 (.I0(x429), .I1(x430), .I2(x431), .I3(n1039), .I4(n1040), .O(n1043));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1044 (.I0(x435), .I1(x436), .I2(x437), .I3(n1042), .I4(n1043), .O(n1044));
  LUT3 #(.INIT(8'h96)) lut_n1045 (.I0(n1029), .I1(n1032), .I2(n1033), .O(n1045));
  LUT3 #(.INIT(8'hE8)) lut_n1046 (.I0(n1041), .I1(n1044), .I2(n1045), .O(n1046));
  LUT3 #(.INIT(8'hE8)) lut_n1047 (.I0(x444), .I1(x445), .I2(x446), .O(n1047));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1048 (.I0(x435), .I1(x436), .I2(x437), .I3(n1042), .I4(n1043), .O(n1048));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1049 (.I0(x441), .I1(x442), .I2(x443), .I3(n1047), .I4(n1048), .O(n1049));
  LUT3 #(.INIT(8'hE8)) lut_n1050 (.I0(x450), .I1(x451), .I2(x452), .O(n1050));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1051 (.I0(x441), .I1(x442), .I2(x443), .I3(n1047), .I4(n1048), .O(n1051));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1052 (.I0(x447), .I1(x448), .I2(x449), .I3(n1050), .I4(n1051), .O(n1052));
  LUT3 #(.INIT(8'h96)) lut_n1053 (.I0(n1041), .I1(n1044), .I2(n1045), .O(n1053));
  LUT3 #(.INIT(8'hE8)) lut_n1054 (.I0(n1049), .I1(n1052), .I2(n1053), .O(n1054));
  LUT3 #(.INIT(8'h96)) lut_n1055 (.I0(n1026), .I1(n1034), .I2(n1035), .O(n1055));
  LUT3 #(.INIT(8'hE8)) lut_n1056 (.I0(n1046), .I1(n1054), .I2(n1055), .O(n1056));
  LUT3 #(.INIT(8'hE8)) lut_n1057 (.I0(x456), .I1(x457), .I2(x458), .O(n1057));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1058 (.I0(x447), .I1(x448), .I2(x449), .I3(n1050), .I4(n1051), .O(n1058));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1059 (.I0(x453), .I1(x454), .I2(x455), .I3(n1057), .I4(n1058), .O(n1059));
  LUT3 #(.INIT(8'hE8)) lut_n1060 (.I0(x462), .I1(x463), .I2(x464), .O(n1060));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1061 (.I0(x453), .I1(x454), .I2(x455), .I3(n1057), .I4(n1058), .O(n1061));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1062 (.I0(x459), .I1(x460), .I2(x461), .I3(n1060), .I4(n1061), .O(n1062));
  LUT3 #(.INIT(8'h96)) lut_n1063 (.I0(n1049), .I1(n1052), .I2(n1053), .O(n1063));
  LUT3 #(.INIT(8'hE8)) lut_n1064 (.I0(n1059), .I1(n1062), .I2(n1063), .O(n1064));
  LUT3 #(.INIT(8'hE8)) lut_n1065 (.I0(x468), .I1(x469), .I2(x470), .O(n1065));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1066 (.I0(x459), .I1(x460), .I2(x461), .I3(n1060), .I4(n1061), .O(n1066));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1067 (.I0(x465), .I1(x466), .I2(x467), .I3(n1065), .I4(n1066), .O(n1067));
  LUT3 #(.INIT(8'hE8)) lut_n1068 (.I0(x474), .I1(x475), .I2(x476), .O(n1068));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1069 (.I0(x465), .I1(x466), .I2(x467), .I3(n1065), .I4(n1066), .O(n1069));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1070 (.I0(x471), .I1(x472), .I2(x473), .I3(n1068), .I4(n1069), .O(n1070));
  LUT3 #(.INIT(8'h96)) lut_n1071 (.I0(n1059), .I1(n1062), .I2(n1063), .O(n1071));
  LUT3 #(.INIT(8'hE8)) lut_n1072 (.I0(n1067), .I1(n1070), .I2(n1071), .O(n1072));
  LUT3 #(.INIT(8'h96)) lut_n1073 (.I0(n1046), .I1(n1054), .I2(n1055), .O(n1073));
  LUT3 #(.INIT(8'hE8)) lut_n1074 (.I0(n1064), .I1(n1072), .I2(n1073), .O(n1074));
  LUT3 #(.INIT(8'h96)) lut_n1075 (.I0(n1018), .I1(n1036), .I2(n1037), .O(n1075));
  LUT3 #(.INIT(8'hE8)) lut_n1076 (.I0(n1056), .I1(n1074), .I2(n1075), .O(n1076));
  LUT3 #(.INIT(8'h96)) lut_n1077 (.I0(n959), .I1(n997), .I2(n998), .O(n1077));
  LUT3 #(.INIT(8'hE8)) lut_n1078 (.I0(n1038), .I1(n1076), .I2(n1077), .O(n1078));
  LUT3 #(.INIT(8'hE8)) lut_n1079 (.I0(x480), .I1(x481), .I2(x482), .O(n1079));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1080 (.I0(x471), .I1(x472), .I2(x473), .I3(n1068), .I4(n1069), .O(n1080));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1081 (.I0(x477), .I1(x478), .I2(x479), .I3(n1079), .I4(n1080), .O(n1081));
  LUT3 #(.INIT(8'hE8)) lut_n1082 (.I0(x486), .I1(x487), .I2(x488), .O(n1082));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1083 (.I0(x477), .I1(x478), .I2(x479), .I3(n1079), .I4(n1080), .O(n1083));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1084 (.I0(x483), .I1(x484), .I2(x485), .I3(n1082), .I4(n1083), .O(n1084));
  LUT3 #(.INIT(8'h96)) lut_n1085 (.I0(n1067), .I1(n1070), .I2(n1071), .O(n1085));
  LUT3 #(.INIT(8'hE8)) lut_n1086 (.I0(n1081), .I1(n1084), .I2(n1085), .O(n1086));
  LUT3 #(.INIT(8'hE8)) lut_n1087 (.I0(x492), .I1(x493), .I2(x494), .O(n1087));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1088 (.I0(x483), .I1(x484), .I2(x485), .I3(n1082), .I4(n1083), .O(n1088));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1089 (.I0(x489), .I1(x490), .I2(x491), .I3(n1087), .I4(n1088), .O(n1089));
  LUT3 #(.INIT(8'hE8)) lut_n1090 (.I0(x498), .I1(x499), .I2(x500), .O(n1090));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1091 (.I0(x489), .I1(x490), .I2(x491), .I3(n1087), .I4(n1088), .O(n1091));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1092 (.I0(x495), .I1(x496), .I2(x497), .I3(n1090), .I4(n1091), .O(n1092));
  LUT3 #(.INIT(8'h96)) lut_n1093 (.I0(n1081), .I1(n1084), .I2(n1085), .O(n1093));
  LUT3 #(.INIT(8'hE8)) lut_n1094 (.I0(n1089), .I1(n1092), .I2(n1093), .O(n1094));
  LUT3 #(.INIT(8'h96)) lut_n1095 (.I0(n1064), .I1(n1072), .I2(n1073), .O(n1095));
  LUT3 #(.INIT(8'hE8)) lut_n1096 (.I0(n1086), .I1(n1094), .I2(n1095), .O(n1096));
  LUT3 #(.INIT(8'hE8)) lut_n1097 (.I0(x504), .I1(x505), .I2(x506), .O(n1097));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1098 (.I0(x495), .I1(x496), .I2(x497), .I3(n1090), .I4(n1091), .O(n1098));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1099 (.I0(x501), .I1(x502), .I2(x503), .I3(n1097), .I4(n1098), .O(n1099));
  LUT3 #(.INIT(8'hE8)) lut_n1100 (.I0(x510), .I1(x511), .I2(x512), .O(n1100));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1101 (.I0(x501), .I1(x502), .I2(x503), .I3(n1097), .I4(n1098), .O(n1101));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1102 (.I0(x507), .I1(x508), .I2(x509), .I3(n1100), .I4(n1101), .O(n1102));
  LUT3 #(.INIT(8'h96)) lut_n1103 (.I0(n1089), .I1(n1092), .I2(n1093), .O(n1103));
  LUT3 #(.INIT(8'hE8)) lut_n1104 (.I0(n1099), .I1(n1102), .I2(n1103), .O(n1104));
  LUT3 #(.INIT(8'hE8)) lut_n1105 (.I0(x516), .I1(x517), .I2(x518), .O(n1105));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1106 (.I0(x507), .I1(x508), .I2(x509), .I3(n1100), .I4(n1101), .O(n1106));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1107 (.I0(x513), .I1(x514), .I2(x515), .I3(n1105), .I4(n1106), .O(n1107));
  LUT3 #(.INIT(8'hE8)) lut_n1108 (.I0(x522), .I1(x523), .I2(x524), .O(n1108));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1109 (.I0(x513), .I1(x514), .I2(x515), .I3(n1105), .I4(n1106), .O(n1109));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1110 (.I0(x519), .I1(x520), .I2(x521), .I3(n1108), .I4(n1109), .O(n1110));
  LUT3 #(.INIT(8'h96)) lut_n1111 (.I0(n1099), .I1(n1102), .I2(n1103), .O(n1111));
  LUT3 #(.INIT(8'hE8)) lut_n1112 (.I0(n1107), .I1(n1110), .I2(n1111), .O(n1112));
  LUT3 #(.INIT(8'h96)) lut_n1113 (.I0(n1086), .I1(n1094), .I2(n1095), .O(n1113));
  LUT3 #(.INIT(8'hE8)) lut_n1114 (.I0(n1104), .I1(n1112), .I2(n1113), .O(n1114));
  LUT3 #(.INIT(8'h96)) lut_n1115 (.I0(n1056), .I1(n1074), .I2(n1075), .O(n1115));
  LUT3 #(.INIT(8'hE8)) lut_n1116 (.I0(n1096), .I1(n1114), .I2(n1115), .O(n1116));
  LUT3 #(.INIT(8'hE8)) lut_n1117 (.I0(x528), .I1(x529), .I2(x530), .O(n1117));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1118 (.I0(x519), .I1(x520), .I2(x521), .I3(n1108), .I4(n1109), .O(n1118));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1119 (.I0(x525), .I1(x526), .I2(x527), .I3(n1117), .I4(n1118), .O(n1119));
  LUT3 #(.INIT(8'hE8)) lut_n1120 (.I0(x534), .I1(x535), .I2(x536), .O(n1120));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1121 (.I0(x525), .I1(x526), .I2(x527), .I3(n1117), .I4(n1118), .O(n1121));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1122 (.I0(x531), .I1(x532), .I2(x533), .I3(n1120), .I4(n1121), .O(n1122));
  LUT3 #(.INIT(8'h96)) lut_n1123 (.I0(n1107), .I1(n1110), .I2(n1111), .O(n1123));
  LUT3 #(.INIT(8'hE8)) lut_n1124 (.I0(n1119), .I1(n1122), .I2(n1123), .O(n1124));
  LUT3 #(.INIT(8'hE8)) lut_n1125 (.I0(x540), .I1(x541), .I2(x542), .O(n1125));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1126 (.I0(x531), .I1(x532), .I2(x533), .I3(n1120), .I4(n1121), .O(n1126));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1127 (.I0(x537), .I1(x538), .I2(x539), .I3(n1125), .I4(n1126), .O(n1127));
  LUT3 #(.INIT(8'hE8)) lut_n1128 (.I0(x546), .I1(x547), .I2(x548), .O(n1128));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1129 (.I0(x537), .I1(x538), .I2(x539), .I3(n1125), .I4(n1126), .O(n1129));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1130 (.I0(x543), .I1(x544), .I2(x545), .I3(n1128), .I4(n1129), .O(n1130));
  LUT3 #(.INIT(8'h96)) lut_n1131 (.I0(n1119), .I1(n1122), .I2(n1123), .O(n1131));
  LUT3 #(.INIT(8'hE8)) lut_n1132 (.I0(n1127), .I1(n1130), .I2(n1131), .O(n1132));
  LUT3 #(.INIT(8'h96)) lut_n1133 (.I0(n1104), .I1(n1112), .I2(n1113), .O(n1133));
  LUT3 #(.INIT(8'hE8)) lut_n1134 (.I0(n1124), .I1(n1132), .I2(n1133), .O(n1134));
  LUT3 #(.INIT(8'hE8)) lut_n1135 (.I0(x552), .I1(x553), .I2(x554), .O(n1135));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1136 (.I0(x543), .I1(x544), .I2(x545), .I3(n1128), .I4(n1129), .O(n1136));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1137 (.I0(x549), .I1(x550), .I2(x551), .I3(n1135), .I4(n1136), .O(n1137));
  LUT3 #(.INIT(8'hE8)) lut_n1138 (.I0(x558), .I1(x559), .I2(x560), .O(n1138));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1139 (.I0(x549), .I1(x550), .I2(x551), .I3(n1135), .I4(n1136), .O(n1139));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1140 (.I0(x555), .I1(x556), .I2(x557), .I3(n1138), .I4(n1139), .O(n1140));
  LUT3 #(.INIT(8'h96)) lut_n1141 (.I0(n1127), .I1(n1130), .I2(n1131), .O(n1141));
  LUT3 #(.INIT(8'hE8)) lut_n1142 (.I0(n1137), .I1(n1140), .I2(n1141), .O(n1142));
  LUT3 #(.INIT(8'hE8)) lut_n1143 (.I0(x564), .I1(x565), .I2(x566), .O(n1143));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1144 (.I0(x555), .I1(x556), .I2(x557), .I3(n1138), .I4(n1139), .O(n1144));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1145 (.I0(x561), .I1(x562), .I2(x563), .I3(n1143), .I4(n1144), .O(n1145));
  LUT3 #(.INIT(8'hE8)) lut_n1146 (.I0(x570), .I1(x571), .I2(x572), .O(n1146));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1147 (.I0(x561), .I1(x562), .I2(x563), .I3(n1143), .I4(n1144), .O(n1147));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1148 (.I0(x567), .I1(x568), .I2(x569), .I3(n1146), .I4(n1147), .O(n1148));
  LUT3 #(.INIT(8'h96)) lut_n1149 (.I0(n1137), .I1(n1140), .I2(n1141), .O(n1149));
  LUT3 #(.INIT(8'hE8)) lut_n1150 (.I0(n1145), .I1(n1148), .I2(n1149), .O(n1150));
  LUT3 #(.INIT(8'h96)) lut_n1151 (.I0(n1124), .I1(n1132), .I2(n1133), .O(n1151));
  LUT3 #(.INIT(8'hE8)) lut_n1152 (.I0(n1142), .I1(n1150), .I2(n1151), .O(n1152));
  LUT3 #(.INIT(8'h96)) lut_n1153 (.I0(n1096), .I1(n1114), .I2(n1115), .O(n1153));
  LUT3 #(.INIT(8'hE8)) lut_n1154 (.I0(n1134), .I1(n1152), .I2(n1153), .O(n1154));
  LUT3 #(.INIT(8'h96)) lut_n1155 (.I0(n1038), .I1(n1076), .I2(n1077), .O(n1155));
  LUT3 #(.INIT(8'hE8)) lut_n1156 (.I0(n1116), .I1(n1154), .I2(n1155), .O(n1156));
  LUT3 #(.INIT(8'h96)) lut_n1157 (.I0(n843), .I1(n921), .I2(n999), .O(n1157));
  LUT3 #(.INIT(8'hE8)) lut_n1158 (.I0(n1078), .I1(n1156), .I2(n1157), .O(n1158));
  LUT3 #(.INIT(8'hE8)) lut_n1159 (.I0(x576), .I1(x577), .I2(x578), .O(n1159));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1160 (.I0(x567), .I1(x568), .I2(x569), .I3(n1146), .I4(n1147), .O(n1160));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1161 (.I0(x573), .I1(x574), .I2(x575), .I3(n1159), .I4(n1160), .O(n1161));
  LUT3 #(.INIT(8'hE8)) lut_n1162 (.I0(x582), .I1(x583), .I2(x584), .O(n1162));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1163 (.I0(x573), .I1(x574), .I2(x575), .I3(n1159), .I4(n1160), .O(n1163));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1164 (.I0(x579), .I1(x580), .I2(x581), .I3(n1162), .I4(n1163), .O(n1164));
  LUT3 #(.INIT(8'h96)) lut_n1165 (.I0(n1145), .I1(n1148), .I2(n1149), .O(n1165));
  LUT3 #(.INIT(8'hE8)) lut_n1166 (.I0(n1161), .I1(n1164), .I2(n1165), .O(n1166));
  LUT3 #(.INIT(8'hE8)) lut_n1167 (.I0(x588), .I1(x589), .I2(x590), .O(n1167));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1168 (.I0(x579), .I1(x580), .I2(x581), .I3(n1162), .I4(n1163), .O(n1168));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1169 (.I0(x585), .I1(x586), .I2(x587), .I3(n1167), .I4(n1168), .O(n1169));
  LUT3 #(.INIT(8'hE8)) lut_n1170 (.I0(x594), .I1(x595), .I2(x596), .O(n1170));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1171 (.I0(x585), .I1(x586), .I2(x587), .I3(n1167), .I4(n1168), .O(n1171));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1172 (.I0(x591), .I1(x592), .I2(x593), .I3(n1170), .I4(n1171), .O(n1172));
  LUT3 #(.INIT(8'h96)) lut_n1173 (.I0(n1161), .I1(n1164), .I2(n1165), .O(n1173));
  LUT3 #(.INIT(8'hE8)) lut_n1174 (.I0(n1169), .I1(n1172), .I2(n1173), .O(n1174));
  LUT3 #(.INIT(8'h96)) lut_n1175 (.I0(n1142), .I1(n1150), .I2(n1151), .O(n1175));
  LUT3 #(.INIT(8'hE8)) lut_n1176 (.I0(n1166), .I1(n1174), .I2(n1175), .O(n1176));
  LUT3 #(.INIT(8'hE8)) lut_n1177 (.I0(x600), .I1(x601), .I2(x602), .O(n1177));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1178 (.I0(x591), .I1(x592), .I2(x593), .I3(n1170), .I4(n1171), .O(n1178));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1179 (.I0(x597), .I1(x598), .I2(x599), .I3(n1177), .I4(n1178), .O(n1179));
  LUT3 #(.INIT(8'hE8)) lut_n1180 (.I0(x606), .I1(x607), .I2(x608), .O(n1180));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1181 (.I0(x597), .I1(x598), .I2(x599), .I3(n1177), .I4(n1178), .O(n1181));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1182 (.I0(x603), .I1(x604), .I2(x605), .I3(n1180), .I4(n1181), .O(n1182));
  LUT3 #(.INIT(8'h96)) lut_n1183 (.I0(n1169), .I1(n1172), .I2(n1173), .O(n1183));
  LUT3 #(.INIT(8'hE8)) lut_n1184 (.I0(n1179), .I1(n1182), .I2(n1183), .O(n1184));
  LUT3 #(.INIT(8'hE8)) lut_n1185 (.I0(x612), .I1(x613), .I2(x614), .O(n1185));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1186 (.I0(x603), .I1(x604), .I2(x605), .I3(n1180), .I4(n1181), .O(n1186));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1187 (.I0(x609), .I1(x610), .I2(x611), .I3(n1185), .I4(n1186), .O(n1187));
  LUT3 #(.INIT(8'hE8)) lut_n1188 (.I0(x618), .I1(x619), .I2(x620), .O(n1188));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1189 (.I0(x609), .I1(x610), .I2(x611), .I3(n1185), .I4(n1186), .O(n1189));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1190 (.I0(x615), .I1(x616), .I2(x617), .I3(n1188), .I4(n1189), .O(n1190));
  LUT3 #(.INIT(8'h96)) lut_n1191 (.I0(n1179), .I1(n1182), .I2(n1183), .O(n1191));
  LUT3 #(.INIT(8'hE8)) lut_n1192 (.I0(n1187), .I1(n1190), .I2(n1191), .O(n1192));
  LUT3 #(.INIT(8'h96)) lut_n1193 (.I0(n1166), .I1(n1174), .I2(n1175), .O(n1193));
  LUT3 #(.INIT(8'hE8)) lut_n1194 (.I0(n1184), .I1(n1192), .I2(n1193), .O(n1194));
  LUT3 #(.INIT(8'h96)) lut_n1195 (.I0(n1134), .I1(n1152), .I2(n1153), .O(n1195));
  LUT3 #(.INIT(8'hE8)) lut_n1196 (.I0(n1176), .I1(n1194), .I2(n1195), .O(n1196));
  LUT3 #(.INIT(8'hE8)) lut_n1197 (.I0(x624), .I1(x625), .I2(x626), .O(n1197));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1198 (.I0(x615), .I1(x616), .I2(x617), .I3(n1188), .I4(n1189), .O(n1198));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1199 (.I0(x621), .I1(x622), .I2(x623), .I3(n1197), .I4(n1198), .O(n1199));
  LUT3 #(.INIT(8'hE8)) lut_n1200 (.I0(x630), .I1(x631), .I2(x632), .O(n1200));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1201 (.I0(x621), .I1(x622), .I2(x623), .I3(n1197), .I4(n1198), .O(n1201));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1202 (.I0(x627), .I1(x628), .I2(x629), .I3(n1200), .I4(n1201), .O(n1202));
  LUT3 #(.INIT(8'h96)) lut_n1203 (.I0(n1187), .I1(n1190), .I2(n1191), .O(n1203));
  LUT3 #(.INIT(8'hE8)) lut_n1204 (.I0(n1199), .I1(n1202), .I2(n1203), .O(n1204));
  LUT3 #(.INIT(8'hE8)) lut_n1205 (.I0(x636), .I1(x637), .I2(x638), .O(n1205));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1206 (.I0(x627), .I1(x628), .I2(x629), .I3(n1200), .I4(n1201), .O(n1206));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1207 (.I0(x633), .I1(x634), .I2(x635), .I3(n1205), .I4(n1206), .O(n1207));
  LUT3 #(.INIT(8'hE8)) lut_n1208 (.I0(x642), .I1(x643), .I2(x644), .O(n1208));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1209 (.I0(x633), .I1(x634), .I2(x635), .I3(n1205), .I4(n1206), .O(n1209));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1210 (.I0(x639), .I1(x640), .I2(x641), .I3(n1208), .I4(n1209), .O(n1210));
  LUT3 #(.INIT(8'h96)) lut_n1211 (.I0(n1199), .I1(n1202), .I2(n1203), .O(n1211));
  LUT3 #(.INIT(8'hE8)) lut_n1212 (.I0(n1207), .I1(n1210), .I2(n1211), .O(n1212));
  LUT3 #(.INIT(8'h96)) lut_n1213 (.I0(n1184), .I1(n1192), .I2(n1193), .O(n1213));
  LUT3 #(.INIT(8'hE8)) lut_n1214 (.I0(n1204), .I1(n1212), .I2(n1213), .O(n1214));
  LUT3 #(.INIT(8'hE8)) lut_n1215 (.I0(x648), .I1(x649), .I2(x650), .O(n1215));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1216 (.I0(x639), .I1(x640), .I2(x641), .I3(n1208), .I4(n1209), .O(n1216));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1217 (.I0(x645), .I1(x646), .I2(x647), .I3(n1215), .I4(n1216), .O(n1217));
  LUT3 #(.INIT(8'hE8)) lut_n1218 (.I0(x654), .I1(x655), .I2(x656), .O(n1218));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1219 (.I0(x645), .I1(x646), .I2(x647), .I3(n1215), .I4(n1216), .O(n1219));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1220 (.I0(x651), .I1(x652), .I2(x653), .I3(n1218), .I4(n1219), .O(n1220));
  LUT3 #(.INIT(8'h96)) lut_n1221 (.I0(n1207), .I1(n1210), .I2(n1211), .O(n1221));
  LUT3 #(.INIT(8'hE8)) lut_n1222 (.I0(n1217), .I1(n1220), .I2(n1221), .O(n1222));
  LUT3 #(.INIT(8'hE8)) lut_n1223 (.I0(x660), .I1(x661), .I2(x662), .O(n1223));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1224 (.I0(x651), .I1(x652), .I2(x653), .I3(n1218), .I4(n1219), .O(n1224));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1225 (.I0(x657), .I1(x658), .I2(x659), .I3(n1223), .I4(n1224), .O(n1225));
  LUT3 #(.INIT(8'hE8)) lut_n1226 (.I0(x666), .I1(x667), .I2(x668), .O(n1226));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1227 (.I0(x657), .I1(x658), .I2(x659), .I3(n1223), .I4(n1224), .O(n1227));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1228 (.I0(x663), .I1(x664), .I2(x665), .I3(n1226), .I4(n1227), .O(n1228));
  LUT3 #(.INIT(8'h96)) lut_n1229 (.I0(n1217), .I1(n1220), .I2(n1221), .O(n1229));
  LUT3 #(.INIT(8'hE8)) lut_n1230 (.I0(n1225), .I1(n1228), .I2(n1229), .O(n1230));
  LUT3 #(.INIT(8'h96)) lut_n1231 (.I0(n1204), .I1(n1212), .I2(n1213), .O(n1231));
  LUT3 #(.INIT(8'hE8)) lut_n1232 (.I0(n1222), .I1(n1230), .I2(n1231), .O(n1232));
  LUT3 #(.INIT(8'h96)) lut_n1233 (.I0(n1176), .I1(n1194), .I2(n1195), .O(n1233));
  LUT3 #(.INIT(8'hE8)) lut_n1234 (.I0(n1214), .I1(n1232), .I2(n1233), .O(n1234));
  LUT3 #(.INIT(8'h96)) lut_n1235 (.I0(n1116), .I1(n1154), .I2(n1155), .O(n1235));
  LUT3 #(.INIT(8'hE8)) lut_n1236 (.I0(n1196), .I1(n1234), .I2(n1235), .O(n1236));
  LUT3 #(.INIT(8'hE8)) lut_n1237 (.I0(x672), .I1(x673), .I2(x674), .O(n1237));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1238 (.I0(x663), .I1(x664), .I2(x665), .I3(n1226), .I4(n1227), .O(n1238));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1239 (.I0(x669), .I1(x670), .I2(x671), .I3(n1237), .I4(n1238), .O(n1239));
  LUT3 #(.INIT(8'hE8)) lut_n1240 (.I0(x678), .I1(x679), .I2(x680), .O(n1240));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1241 (.I0(x669), .I1(x670), .I2(x671), .I3(n1237), .I4(n1238), .O(n1241));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1242 (.I0(x675), .I1(x676), .I2(x677), .I3(n1240), .I4(n1241), .O(n1242));
  LUT3 #(.INIT(8'h96)) lut_n1243 (.I0(n1225), .I1(n1228), .I2(n1229), .O(n1243));
  LUT3 #(.INIT(8'hE8)) lut_n1244 (.I0(n1239), .I1(n1242), .I2(n1243), .O(n1244));
  LUT3 #(.INIT(8'hE8)) lut_n1245 (.I0(x684), .I1(x685), .I2(x686), .O(n1245));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1246 (.I0(x675), .I1(x676), .I2(x677), .I3(n1240), .I4(n1241), .O(n1246));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1247 (.I0(x681), .I1(x682), .I2(x683), .I3(n1245), .I4(n1246), .O(n1247));
  LUT3 #(.INIT(8'hE8)) lut_n1248 (.I0(x690), .I1(x691), .I2(x692), .O(n1248));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1249 (.I0(x681), .I1(x682), .I2(x683), .I3(n1245), .I4(n1246), .O(n1249));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1250 (.I0(x687), .I1(x688), .I2(x689), .I3(n1248), .I4(n1249), .O(n1250));
  LUT3 #(.INIT(8'h96)) lut_n1251 (.I0(n1239), .I1(n1242), .I2(n1243), .O(n1251));
  LUT3 #(.INIT(8'hE8)) lut_n1252 (.I0(n1247), .I1(n1250), .I2(n1251), .O(n1252));
  LUT3 #(.INIT(8'h96)) lut_n1253 (.I0(n1222), .I1(n1230), .I2(n1231), .O(n1253));
  LUT3 #(.INIT(8'hE8)) lut_n1254 (.I0(n1244), .I1(n1252), .I2(n1253), .O(n1254));
  LUT3 #(.INIT(8'hE8)) lut_n1255 (.I0(x696), .I1(x697), .I2(x698), .O(n1255));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1256 (.I0(x687), .I1(x688), .I2(x689), .I3(n1248), .I4(n1249), .O(n1256));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1257 (.I0(x693), .I1(x694), .I2(x695), .I3(n1255), .I4(n1256), .O(n1257));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1258 (.I0(x693), .I1(x694), .I2(x695), .I3(n1255), .I4(n1256), .O(n1258));
  LUT3 #(.INIT(8'hFE)) lut_n1259 (.I0(x699), .I1(x700), .I2(n1258), .O(n1259));
  LUT3 #(.INIT(8'h96)) lut_n1260 (.I0(n1247), .I1(n1250), .I2(n1251), .O(n1260));
  LUT3 #(.INIT(8'hE8)) lut_n1261 (.I0(n1257), .I1(n1259), .I2(n1260), .O(n1261));
  LUT3 #(.INIT(8'h96)) lut_n1262 (.I0(n1244), .I1(n1252), .I2(n1253), .O(n1262));
  LUT2 #(.INIT(4'hE)) lut_n1263 (.I0(n1261), .I1(n1262), .O(n1263));
  LUT3 #(.INIT(8'h96)) lut_n1264 (.I0(n1214), .I1(n1232), .I2(n1233), .O(n1264));
  LUT3 #(.INIT(8'hE8)) lut_n1265 (.I0(n1254), .I1(n1263), .I2(n1264), .O(n1265));
  LUT3 #(.INIT(8'h96)) lut_n1266 (.I0(n1196), .I1(n1234), .I2(n1235), .O(n1266));
  LUT2 #(.INIT(4'hE)) lut_n1267 (.I0(n1265), .I1(n1266), .O(n1267));
  LUT3 #(.INIT(8'h96)) lut_n1268 (.I0(n1078), .I1(n1156), .I2(n1157), .O(n1268));
  LUT3 #(.INIT(8'hE8)) lut_n1269 (.I0(n1236), .I1(n1267), .I2(n1268), .O(n1269));
  LUT3 #(.INIT(8'h96)) lut_n1270 (.I0(n1236), .I1(n1267), .I2(n1268), .O(n1270));
  LUT3 #(.INIT(8'h96)) lut_n1271 (.I0(x0), .I1(x1), .I2(x2), .O(n1271));
  LUT3 #(.INIT(8'h96)) lut_n1272 (.I0(x6), .I1(x7), .I2(x8), .O(n1272));
  LUT5 #(.INIT(32'hFF969600)) lut_n1273 (.I0(x3), .I1(x4), .I2(x5), .I3(n1271), .I4(n1272), .O(n1273));
  LUT3 #(.INIT(8'h96)) lut_n1274 (.I0(x12), .I1(x13), .I2(x14), .O(n1274));
  LUT5 #(.INIT(32'h96696996)) lut_n1275 (.I0(x3), .I1(x4), .I2(x5), .I3(n1271), .I4(n1272), .O(n1275));
  LUT5 #(.INIT(32'hFF969600)) lut_n1276 (.I0(x9), .I1(x10), .I2(x11), .I3(n1274), .I4(n1275), .O(n1276));
  LUT3 #(.INIT(8'h1E)) lut_n1277 (.I0(x699), .I1(x700), .I2(n1258), .O(n1277));
  LUT3 #(.INIT(8'h8E)) lut_n1278 (.I0(n1273), .I1(n1276), .I2(n1277), .O(n1278));
  LUT3 #(.INIT(8'h96)) lut_n1279 (.I0(n1257), .I1(n1259), .I2(n1260), .O(n1279));
  LUT2 #(.INIT(4'h8)) lut_n1280 (.I0(n1278), .I1(n1279), .O(n1280));
  LUT2 #(.INIT(4'h6)) lut_n1281 (.I0(n1261), .I1(n1262), .O(n1281));
  LUT2 #(.INIT(4'h2)) lut_n1282 (.I0(n1280), .I1(n1281), .O(n1282));
  LUT3 #(.INIT(8'h96)) lut_n1283 (.I0(x18), .I1(x19), .I2(x20), .O(n1283));
  LUT5 #(.INIT(32'h96696996)) lut_n1284 (.I0(x9), .I1(x10), .I2(x11), .I3(n1274), .I4(n1275), .O(n1284));
  LUT5 #(.INIT(32'hFF969600)) lut_n1285 (.I0(x15), .I1(x16), .I2(x17), .I3(n1283), .I4(n1284), .O(n1285));
  LUT3 #(.INIT(8'h96)) lut_n1286 (.I0(x24), .I1(x25), .I2(x26), .O(n1286));
  LUT5 #(.INIT(32'h96696996)) lut_n1287 (.I0(x15), .I1(x16), .I2(x17), .I3(n1283), .I4(n1284), .O(n1287));
  LUT5 #(.INIT(32'hFF969600)) lut_n1288 (.I0(x21), .I1(x22), .I2(x23), .I3(n1286), .I4(n1287), .O(n1288));
  LUT3 #(.INIT(8'h96)) lut_n1289 (.I0(n1273), .I1(n1276), .I2(n1277), .O(n1289));
  LUT3 #(.INIT(8'h8E)) lut_n1290 (.I0(n1285), .I1(n1288), .I2(n1289), .O(n1290));
  LUT3 #(.INIT(8'h96)) lut_n1291 (.I0(x27), .I1(x28), .I2(x29), .O(n1291));
  LUT5 #(.INIT(32'h96696996)) lut_n1292 (.I0(x21), .I1(x22), .I2(x23), .I3(n1286), .I4(n1287), .O(n1292));
  LUT5 #(.INIT(32'hFF969600)) lut_n1293 (.I0(x30), .I1(x31), .I2(x32), .I3(n1291), .I4(n1292), .O(n1293));
  LUT3 #(.INIT(8'h96)) lut_n1294 (.I0(x36), .I1(x37), .I2(x38), .O(n1294));
  LUT5 #(.INIT(32'h96696996)) lut_n1295 (.I0(x30), .I1(x31), .I2(x32), .I3(n1291), .I4(n1292), .O(n1295));
  LUT5 #(.INIT(32'hFF969600)) lut_n1296 (.I0(x33), .I1(x34), .I2(x35), .I3(n1294), .I4(n1295), .O(n1296));
  LUT3 #(.INIT(8'h96)) lut_n1297 (.I0(n1285), .I1(n1288), .I2(n1289), .O(n1297));
  LUT3 #(.INIT(8'h8E)) lut_n1298 (.I0(n1293), .I1(n1296), .I2(n1297), .O(n1298));
  LUT2 #(.INIT(4'h6)) lut_n1299 (.I0(n1278), .I1(n1279), .O(n1299));
  LUT3 #(.INIT(8'hE8)) lut_n1300 (.I0(n1290), .I1(n1298), .I2(n1299), .O(n1300));
  LUT3 #(.INIT(8'h96)) lut_n1301 (.I0(x42), .I1(x43), .I2(x44), .O(n1301));
  LUT5 #(.INIT(32'h96696996)) lut_n1302 (.I0(x33), .I1(x34), .I2(x35), .I3(n1294), .I4(n1295), .O(n1302));
  LUT5 #(.INIT(32'hFF969600)) lut_n1303 (.I0(x39), .I1(x40), .I2(x41), .I3(n1301), .I4(n1302), .O(n1303));
  LUT3 #(.INIT(8'h96)) lut_n1304 (.I0(x48), .I1(x49), .I2(x50), .O(n1304));
  LUT5 #(.INIT(32'h96696996)) lut_n1305 (.I0(x39), .I1(x40), .I2(x41), .I3(n1301), .I4(n1302), .O(n1305));
  LUT5 #(.INIT(32'hFF969600)) lut_n1306 (.I0(x45), .I1(x46), .I2(x47), .I3(n1304), .I4(n1305), .O(n1306));
  LUT3 #(.INIT(8'h96)) lut_n1307 (.I0(n1293), .I1(n1296), .I2(n1297), .O(n1307));
  LUT3 #(.INIT(8'h8E)) lut_n1308 (.I0(n1303), .I1(n1306), .I2(n1307), .O(n1308));
  LUT3 #(.INIT(8'h96)) lut_n1309 (.I0(x54), .I1(x55), .I2(x56), .O(n1309));
  LUT5 #(.INIT(32'h96696996)) lut_n1310 (.I0(x45), .I1(x46), .I2(x47), .I3(n1304), .I4(n1305), .O(n1310));
  LUT5 #(.INIT(32'hFF969600)) lut_n1311 (.I0(x51), .I1(x52), .I2(x53), .I3(n1309), .I4(n1310), .O(n1311));
  LUT3 #(.INIT(8'h96)) lut_n1312 (.I0(x60), .I1(x61), .I2(x62), .O(n1312));
  LUT5 #(.INIT(32'h96696996)) lut_n1313 (.I0(x51), .I1(x52), .I2(x53), .I3(n1309), .I4(n1310), .O(n1313));
  LUT5 #(.INIT(32'hFF969600)) lut_n1314 (.I0(x57), .I1(x58), .I2(x59), .I3(n1312), .I4(n1313), .O(n1314));
  LUT3 #(.INIT(8'h96)) lut_n1315 (.I0(n1303), .I1(n1306), .I2(n1307), .O(n1315));
  LUT3 #(.INIT(8'h8E)) lut_n1316 (.I0(n1311), .I1(n1314), .I2(n1315), .O(n1316));
  LUT3 #(.INIT(8'h96)) lut_n1317 (.I0(n1290), .I1(n1298), .I2(n1299), .O(n1317));
  LUT3 #(.INIT(8'hE8)) lut_n1318 (.I0(n1308), .I1(n1316), .I2(n1317), .O(n1318));
  LUT2 #(.INIT(4'h6)) lut_n1319 (.I0(n1280), .I1(n1281), .O(n1319));
  LUT3 #(.INIT(8'h8E)) lut_n1320 (.I0(n1300), .I1(n1318), .I2(n1319), .O(n1320));
  LUT3 #(.INIT(8'h96)) lut_n1321 (.I0(n1254), .I1(n1263), .I2(n1264), .O(n1321));
  LUT3 #(.INIT(8'hE8)) lut_n1322 (.I0(n1282), .I1(n1320), .I2(n1321), .O(n1322));
  LUT2 #(.INIT(4'h6)) lut_n1323 (.I0(n1265), .I1(n1266), .O(n1323));
  LUT2 #(.INIT(4'h2)) lut_n1324 (.I0(n1322), .I1(n1323), .O(n1324));
  LUT3 #(.INIT(8'h96)) lut_n1325 (.I0(x66), .I1(x67), .I2(x68), .O(n1325));
  LUT5 #(.INIT(32'h96696996)) lut_n1326 (.I0(x57), .I1(x58), .I2(x59), .I3(n1312), .I4(n1313), .O(n1326));
  LUT5 #(.INIT(32'hFF969600)) lut_n1327 (.I0(x63), .I1(x64), .I2(x65), .I3(n1325), .I4(n1326), .O(n1327));
  LUT3 #(.INIT(8'h96)) lut_n1328 (.I0(x72), .I1(x73), .I2(x74), .O(n1328));
  LUT5 #(.INIT(32'h96696996)) lut_n1329 (.I0(x63), .I1(x64), .I2(x65), .I3(n1325), .I4(n1326), .O(n1329));
  LUT5 #(.INIT(32'hFF969600)) lut_n1330 (.I0(x69), .I1(x70), .I2(x71), .I3(n1328), .I4(n1329), .O(n1330));
  LUT3 #(.INIT(8'h96)) lut_n1331 (.I0(n1311), .I1(n1314), .I2(n1315), .O(n1331));
  LUT3 #(.INIT(8'h8E)) lut_n1332 (.I0(n1327), .I1(n1330), .I2(n1331), .O(n1332));
  LUT3 #(.INIT(8'h96)) lut_n1333 (.I0(x78), .I1(x79), .I2(x80), .O(n1333));
  LUT5 #(.INIT(32'h96696996)) lut_n1334 (.I0(x69), .I1(x70), .I2(x71), .I3(n1328), .I4(n1329), .O(n1334));
  LUT5 #(.INIT(32'hFF969600)) lut_n1335 (.I0(x75), .I1(x76), .I2(x77), .I3(n1333), .I4(n1334), .O(n1335));
  LUT3 #(.INIT(8'h96)) lut_n1336 (.I0(x84), .I1(x85), .I2(x86), .O(n1336));
  LUT5 #(.INIT(32'h96696996)) lut_n1337 (.I0(x75), .I1(x76), .I2(x77), .I3(n1333), .I4(n1334), .O(n1337));
  LUT5 #(.INIT(32'hFF969600)) lut_n1338 (.I0(x81), .I1(x82), .I2(x83), .I3(n1336), .I4(n1337), .O(n1338));
  LUT3 #(.INIT(8'h96)) lut_n1339 (.I0(n1327), .I1(n1330), .I2(n1331), .O(n1339));
  LUT3 #(.INIT(8'h8E)) lut_n1340 (.I0(n1335), .I1(n1338), .I2(n1339), .O(n1340));
  LUT3 #(.INIT(8'h96)) lut_n1341 (.I0(n1308), .I1(n1316), .I2(n1317), .O(n1341));
  LUT3 #(.INIT(8'hE8)) lut_n1342 (.I0(n1332), .I1(n1340), .I2(n1341), .O(n1342));
  LUT3 #(.INIT(8'h96)) lut_n1343 (.I0(x90), .I1(x91), .I2(x92), .O(n1343));
  LUT5 #(.INIT(32'h96696996)) lut_n1344 (.I0(x81), .I1(x82), .I2(x83), .I3(n1336), .I4(n1337), .O(n1344));
  LUT5 #(.INIT(32'hFF969600)) lut_n1345 (.I0(x87), .I1(x88), .I2(x89), .I3(n1343), .I4(n1344), .O(n1345));
  LUT3 #(.INIT(8'h96)) lut_n1346 (.I0(x96), .I1(x97), .I2(x98), .O(n1346));
  LUT5 #(.INIT(32'h96696996)) lut_n1347 (.I0(x87), .I1(x88), .I2(x89), .I3(n1343), .I4(n1344), .O(n1347));
  LUT5 #(.INIT(32'hFF969600)) lut_n1348 (.I0(x93), .I1(x94), .I2(x95), .I3(n1346), .I4(n1347), .O(n1348));
  LUT3 #(.INIT(8'h96)) lut_n1349 (.I0(n1335), .I1(n1338), .I2(n1339), .O(n1349));
  LUT3 #(.INIT(8'h8E)) lut_n1350 (.I0(n1345), .I1(n1348), .I2(n1349), .O(n1350));
  LUT3 #(.INIT(8'h96)) lut_n1351 (.I0(x102), .I1(x103), .I2(x104), .O(n1351));
  LUT5 #(.INIT(32'h96696996)) lut_n1352 (.I0(x93), .I1(x94), .I2(x95), .I3(n1346), .I4(n1347), .O(n1352));
  LUT5 #(.INIT(32'hFF969600)) lut_n1353 (.I0(x99), .I1(x100), .I2(x101), .I3(n1351), .I4(n1352), .O(n1353));
  LUT3 #(.INIT(8'h96)) lut_n1354 (.I0(x108), .I1(x109), .I2(x110), .O(n1354));
  LUT5 #(.INIT(32'h96696996)) lut_n1355 (.I0(x99), .I1(x100), .I2(x101), .I3(n1351), .I4(n1352), .O(n1355));
  LUT5 #(.INIT(32'hFF969600)) lut_n1356 (.I0(x105), .I1(x106), .I2(x107), .I3(n1354), .I4(n1355), .O(n1356));
  LUT3 #(.INIT(8'h96)) lut_n1357 (.I0(n1345), .I1(n1348), .I2(n1349), .O(n1357));
  LUT3 #(.INIT(8'h8E)) lut_n1358 (.I0(n1353), .I1(n1356), .I2(n1357), .O(n1358));
  LUT3 #(.INIT(8'h96)) lut_n1359 (.I0(n1332), .I1(n1340), .I2(n1341), .O(n1359));
  LUT3 #(.INIT(8'hE8)) lut_n1360 (.I0(n1350), .I1(n1358), .I2(n1359), .O(n1360));
  LUT3 #(.INIT(8'h96)) lut_n1361 (.I0(n1300), .I1(n1318), .I2(n1319), .O(n1361));
  LUT3 #(.INIT(8'h8E)) lut_n1362 (.I0(n1342), .I1(n1360), .I2(n1361), .O(n1362));
  LUT3 #(.INIT(8'h96)) lut_n1363 (.I0(x114), .I1(x115), .I2(x116), .O(n1363));
  LUT5 #(.INIT(32'h96696996)) lut_n1364 (.I0(x105), .I1(x106), .I2(x107), .I3(n1354), .I4(n1355), .O(n1364));
  LUT5 #(.INIT(32'hFF969600)) lut_n1365 (.I0(x111), .I1(x112), .I2(x113), .I3(n1363), .I4(n1364), .O(n1365));
  LUT3 #(.INIT(8'h96)) lut_n1366 (.I0(x120), .I1(x121), .I2(x122), .O(n1366));
  LUT5 #(.INIT(32'h96696996)) lut_n1367 (.I0(x111), .I1(x112), .I2(x113), .I3(n1363), .I4(n1364), .O(n1367));
  LUT5 #(.INIT(32'hFF969600)) lut_n1368 (.I0(x117), .I1(x118), .I2(x119), .I3(n1366), .I4(n1367), .O(n1368));
  LUT3 #(.INIT(8'h96)) lut_n1369 (.I0(n1353), .I1(n1356), .I2(n1357), .O(n1369));
  LUT3 #(.INIT(8'h8E)) lut_n1370 (.I0(n1365), .I1(n1368), .I2(n1369), .O(n1370));
  LUT3 #(.INIT(8'h96)) lut_n1371 (.I0(x126), .I1(x127), .I2(x128), .O(n1371));
  LUT5 #(.INIT(32'h96696996)) lut_n1372 (.I0(x117), .I1(x118), .I2(x119), .I3(n1366), .I4(n1367), .O(n1372));
  LUT5 #(.INIT(32'hFF969600)) lut_n1373 (.I0(x123), .I1(x124), .I2(x125), .I3(n1371), .I4(n1372), .O(n1373));
  LUT3 #(.INIT(8'h96)) lut_n1374 (.I0(x132), .I1(x133), .I2(x134), .O(n1374));
  LUT5 #(.INIT(32'h96696996)) lut_n1375 (.I0(x123), .I1(x124), .I2(x125), .I3(n1371), .I4(n1372), .O(n1375));
  LUT5 #(.INIT(32'hFF969600)) lut_n1376 (.I0(x129), .I1(x130), .I2(x131), .I3(n1374), .I4(n1375), .O(n1376));
  LUT3 #(.INIT(8'h96)) lut_n1377 (.I0(n1365), .I1(n1368), .I2(n1369), .O(n1377));
  LUT3 #(.INIT(8'h8E)) lut_n1378 (.I0(n1373), .I1(n1376), .I2(n1377), .O(n1378));
  LUT3 #(.INIT(8'h96)) lut_n1379 (.I0(n1350), .I1(n1358), .I2(n1359), .O(n1379));
  LUT3 #(.INIT(8'hE8)) lut_n1380 (.I0(n1370), .I1(n1378), .I2(n1379), .O(n1380));
  LUT3 #(.INIT(8'h96)) lut_n1381 (.I0(x138), .I1(x139), .I2(x140), .O(n1381));
  LUT5 #(.INIT(32'h96696996)) lut_n1382 (.I0(x129), .I1(x130), .I2(x131), .I3(n1374), .I4(n1375), .O(n1382));
  LUT5 #(.INIT(32'hFF969600)) lut_n1383 (.I0(x135), .I1(x136), .I2(x137), .I3(n1381), .I4(n1382), .O(n1383));
  LUT3 #(.INIT(8'h96)) lut_n1384 (.I0(x144), .I1(x145), .I2(x146), .O(n1384));
  LUT5 #(.INIT(32'h96696996)) lut_n1385 (.I0(x135), .I1(x136), .I2(x137), .I3(n1381), .I4(n1382), .O(n1385));
  LUT5 #(.INIT(32'hFF969600)) lut_n1386 (.I0(x141), .I1(x142), .I2(x143), .I3(n1384), .I4(n1385), .O(n1386));
  LUT3 #(.INIT(8'h96)) lut_n1387 (.I0(n1373), .I1(n1376), .I2(n1377), .O(n1387));
  LUT3 #(.INIT(8'h8E)) lut_n1388 (.I0(n1383), .I1(n1386), .I2(n1387), .O(n1388));
  LUT3 #(.INIT(8'h96)) lut_n1389 (.I0(x150), .I1(x151), .I2(x152), .O(n1389));
  LUT5 #(.INIT(32'h96696996)) lut_n1390 (.I0(x141), .I1(x142), .I2(x143), .I3(n1384), .I4(n1385), .O(n1390));
  LUT5 #(.INIT(32'hFF969600)) lut_n1391 (.I0(x147), .I1(x148), .I2(x149), .I3(n1389), .I4(n1390), .O(n1391));
  LUT3 #(.INIT(8'h96)) lut_n1392 (.I0(x156), .I1(x157), .I2(x158), .O(n1392));
  LUT5 #(.INIT(32'h96696996)) lut_n1393 (.I0(x147), .I1(x148), .I2(x149), .I3(n1389), .I4(n1390), .O(n1393));
  LUT5 #(.INIT(32'hFF969600)) lut_n1394 (.I0(x153), .I1(x154), .I2(x155), .I3(n1392), .I4(n1393), .O(n1394));
  LUT3 #(.INIT(8'h96)) lut_n1395 (.I0(n1383), .I1(n1386), .I2(n1387), .O(n1395));
  LUT3 #(.INIT(8'h8E)) lut_n1396 (.I0(n1391), .I1(n1394), .I2(n1395), .O(n1396));
  LUT3 #(.INIT(8'h96)) lut_n1397 (.I0(n1370), .I1(n1378), .I2(n1379), .O(n1397));
  LUT3 #(.INIT(8'hE8)) lut_n1398 (.I0(n1388), .I1(n1396), .I2(n1397), .O(n1398));
  LUT3 #(.INIT(8'h96)) lut_n1399 (.I0(n1342), .I1(n1360), .I2(n1361), .O(n1399));
  LUT3 #(.INIT(8'h8E)) lut_n1400 (.I0(n1380), .I1(n1398), .I2(n1399), .O(n1400));
  LUT3 #(.INIT(8'h96)) lut_n1401 (.I0(n1282), .I1(n1320), .I2(n1321), .O(n1401));
  LUT3 #(.INIT(8'hE8)) lut_n1402 (.I0(n1362), .I1(n1400), .I2(n1401), .O(n1402));
  LUT3 #(.INIT(8'h96)) lut_n1403 (.I0(x162), .I1(x163), .I2(x164), .O(n1403));
  LUT5 #(.INIT(32'h96696996)) lut_n1404 (.I0(x153), .I1(x154), .I2(x155), .I3(n1392), .I4(n1393), .O(n1404));
  LUT5 #(.INIT(32'hFF969600)) lut_n1405 (.I0(x159), .I1(x160), .I2(x161), .I3(n1403), .I4(n1404), .O(n1405));
  LUT3 #(.INIT(8'h96)) lut_n1406 (.I0(x168), .I1(x169), .I2(x170), .O(n1406));
  LUT5 #(.INIT(32'h96696996)) lut_n1407 (.I0(x159), .I1(x160), .I2(x161), .I3(n1403), .I4(n1404), .O(n1407));
  LUT5 #(.INIT(32'hFF969600)) lut_n1408 (.I0(x165), .I1(x166), .I2(x167), .I3(n1406), .I4(n1407), .O(n1408));
  LUT3 #(.INIT(8'h96)) lut_n1409 (.I0(n1391), .I1(n1394), .I2(n1395), .O(n1409));
  LUT3 #(.INIT(8'h8E)) lut_n1410 (.I0(n1405), .I1(n1408), .I2(n1409), .O(n1410));
  LUT3 #(.INIT(8'h96)) lut_n1411 (.I0(x174), .I1(x175), .I2(x176), .O(n1411));
  LUT5 #(.INIT(32'h96696996)) lut_n1412 (.I0(x165), .I1(x166), .I2(x167), .I3(n1406), .I4(n1407), .O(n1412));
  LUT5 #(.INIT(32'hFF969600)) lut_n1413 (.I0(x171), .I1(x172), .I2(x173), .I3(n1411), .I4(n1412), .O(n1413));
  LUT3 #(.INIT(8'h96)) lut_n1414 (.I0(x180), .I1(x181), .I2(x182), .O(n1414));
  LUT5 #(.INIT(32'h96696996)) lut_n1415 (.I0(x171), .I1(x172), .I2(x173), .I3(n1411), .I4(n1412), .O(n1415));
  LUT5 #(.INIT(32'hFF969600)) lut_n1416 (.I0(x177), .I1(x178), .I2(x179), .I3(n1414), .I4(n1415), .O(n1416));
  LUT3 #(.INIT(8'h96)) lut_n1417 (.I0(n1405), .I1(n1408), .I2(n1409), .O(n1417));
  LUT3 #(.INIT(8'h8E)) lut_n1418 (.I0(n1413), .I1(n1416), .I2(n1417), .O(n1418));
  LUT3 #(.INIT(8'h96)) lut_n1419 (.I0(n1388), .I1(n1396), .I2(n1397), .O(n1419));
  LUT3 #(.INIT(8'hE8)) lut_n1420 (.I0(n1410), .I1(n1418), .I2(n1419), .O(n1420));
  LUT3 #(.INIT(8'h96)) lut_n1421 (.I0(x186), .I1(x187), .I2(x188), .O(n1421));
  LUT5 #(.INIT(32'h96696996)) lut_n1422 (.I0(x177), .I1(x178), .I2(x179), .I3(n1414), .I4(n1415), .O(n1422));
  LUT5 #(.INIT(32'hFF969600)) lut_n1423 (.I0(x183), .I1(x184), .I2(x185), .I3(n1421), .I4(n1422), .O(n1423));
  LUT3 #(.INIT(8'h96)) lut_n1424 (.I0(x192), .I1(x193), .I2(x194), .O(n1424));
  LUT5 #(.INIT(32'h96696996)) lut_n1425 (.I0(x183), .I1(x184), .I2(x185), .I3(n1421), .I4(n1422), .O(n1425));
  LUT5 #(.INIT(32'hFF969600)) lut_n1426 (.I0(x189), .I1(x190), .I2(x191), .I3(n1424), .I4(n1425), .O(n1426));
  LUT3 #(.INIT(8'h96)) lut_n1427 (.I0(n1413), .I1(n1416), .I2(n1417), .O(n1427));
  LUT3 #(.INIT(8'h8E)) lut_n1428 (.I0(n1423), .I1(n1426), .I2(n1427), .O(n1428));
  LUT3 #(.INIT(8'h96)) lut_n1429 (.I0(x198), .I1(x199), .I2(x200), .O(n1429));
  LUT5 #(.INIT(32'h96696996)) lut_n1430 (.I0(x189), .I1(x190), .I2(x191), .I3(n1424), .I4(n1425), .O(n1430));
  LUT5 #(.INIT(32'hFF969600)) lut_n1431 (.I0(x195), .I1(x196), .I2(x197), .I3(n1429), .I4(n1430), .O(n1431));
  LUT3 #(.INIT(8'h96)) lut_n1432 (.I0(x204), .I1(x205), .I2(x206), .O(n1432));
  LUT5 #(.INIT(32'h96696996)) lut_n1433 (.I0(x195), .I1(x196), .I2(x197), .I3(n1429), .I4(n1430), .O(n1433));
  LUT5 #(.INIT(32'hFF969600)) lut_n1434 (.I0(x201), .I1(x202), .I2(x203), .I3(n1432), .I4(n1433), .O(n1434));
  LUT3 #(.INIT(8'h96)) lut_n1435 (.I0(n1423), .I1(n1426), .I2(n1427), .O(n1435));
  LUT3 #(.INIT(8'h8E)) lut_n1436 (.I0(n1431), .I1(n1434), .I2(n1435), .O(n1436));
  LUT3 #(.INIT(8'h96)) lut_n1437 (.I0(n1410), .I1(n1418), .I2(n1419), .O(n1437));
  LUT3 #(.INIT(8'hE8)) lut_n1438 (.I0(n1428), .I1(n1436), .I2(n1437), .O(n1438));
  LUT3 #(.INIT(8'h96)) lut_n1439 (.I0(n1380), .I1(n1398), .I2(n1399), .O(n1439));
  LUT3 #(.INIT(8'h8E)) lut_n1440 (.I0(n1420), .I1(n1438), .I2(n1439), .O(n1440));
  LUT3 #(.INIT(8'h96)) lut_n1441 (.I0(x210), .I1(x211), .I2(x212), .O(n1441));
  LUT5 #(.INIT(32'h96696996)) lut_n1442 (.I0(x201), .I1(x202), .I2(x203), .I3(n1432), .I4(n1433), .O(n1442));
  LUT5 #(.INIT(32'hFF969600)) lut_n1443 (.I0(x207), .I1(x208), .I2(x209), .I3(n1441), .I4(n1442), .O(n1443));
  LUT3 #(.INIT(8'h96)) lut_n1444 (.I0(x216), .I1(x217), .I2(x218), .O(n1444));
  LUT5 #(.INIT(32'h96696996)) lut_n1445 (.I0(x207), .I1(x208), .I2(x209), .I3(n1441), .I4(n1442), .O(n1445));
  LUT5 #(.INIT(32'hFF969600)) lut_n1446 (.I0(x213), .I1(x214), .I2(x215), .I3(n1444), .I4(n1445), .O(n1446));
  LUT3 #(.INIT(8'h96)) lut_n1447 (.I0(n1431), .I1(n1434), .I2(n1435), .O(n1447));
  LUT3 #(.INIT(8'h8E)) lut_n1448 (.I0(n1443), .I1(n1446), .I2(n1447), .O(n1448));
  LUT3 #(.INIT(8'h96)) lut_n1449 (.I0(x222), .I1(x223), .I2(x224), .O(n1449));
  LUT5 #(.INIT(32'h96696996)) lut_n1450 (.I0(x213), .I1(x214), .I2(x215), .I3(n1444), .I4(n1445), .O(n1450));
  LUT5 #(.INIT(32'hFF969600)) lut_n1451 (.I0(x219), .I1(x220), .I2(x221), .I3(n1449), .I4(n1450), .O(n1451));
  LUT3 #(.INIT(8'h96)) lut_n1452 (.I0(x228), .I1(x229), .I2(x230), .O(n1452));
  LUT5 #(.INIT(32'h96696996)) lut_n1453 (.I0(x219), .I1(x220), .I2(x221), .I3(n1449), .I4(n1450), .O(n1453));
  LUT5 #(.INIT(32'hFF969600)) lut_n1454 (.I0(x225), .I1(x226), .I2(x227), .I3(n1452), .I4(n1453), .O(n1454));
  LUT3 #(.INIT(8'h96)) lut_n1455 (.I0(n1443), .I1(n1446), .I2(n1447), .O(n1455));
  LUT3 #(.INIT(8'h8E)) lut_n1456 (.I0(n1451), .I1(n1454), .I2(n1455), .O(n1456));
  LUT3 #(.INIT(8'h96)) lut_n1457 (.I0(n1428), .I1(n1436), .I2(n1437), .O(n1457));
  LUT3 #(.INIT(8'hE8)) lut_n1458 (.I0(n1448), .I1(n1456), .I2(n1457), .O(n1458));
  LUT3 #(.INIT(8'h96)) lut_n1459 (.I0(x234), .I1(x235), .I2(x236), .O(n1459));
  LUT5 #(.INIT(32'h96696996)) lut_n1460 (.I0(x225), .I1(x226), .I2(x227), .I3(n1452), .I4(n1453), .O(n1460));
  LUT5 #(.INIT(32'hFF969600)) lut_n1461 (.I0(x231), .I1(x232), .I2(x233), .I3(n1459), .I4(n1460), .O(n1461));
  LUT3 #(.INIT(8'h96)) lut_n1462 (.I0(x240), .I1(x241), .I2(x242), .O(n1462));
  LUT5 #(.INIT(32'h96696996)) lut_n1463 (.I0(x231), .I1(x232), .I2(x233), .I3(n1459), .I4(n1460), .O(n1463));
  LUT5 #(.INIT(32'hFF969600)) lut_n1464 (.I0(x237), .I1(x238), .I2(x239), .I3(n1462), .I4(n1463), .O(n1464));
  LUT3 #(.INIT(8'h96)) lut_n1465 (.I0(n1451), .I1(n1454), .I2(n1455), .O(n1465));
  LUT3 #(.INIT(8'h8E)) lut_n1466 (.I0(n1461), .I1(n1464), .I2(n1465), .O(n1466));
  LUT3 #(.INIT(8'h96)) lut_n1467 (.I0(x246), .I1(x247), .I2(x248), .O(n1467));
  LUT5 #(.INIT(32'h96696996)) lut_n1468 (.I0(x237), .I1(x238), .I2(x239), .I3(n1462), .I4(n1463), .O(n1468));
  LUT5 #(.INIT(32'hFF969600)) lut_n1469 (.I0(x243), .I1(x244), .I2(x245), .I3(n1467), .I4(n1468), .O(n1469));
  LUT3 #(.INIT(8'h96)) lut_n1470 (.I0(x252), .I1(x253), .I2(x254), .O(n1470));
  LUT5 #(.INIT(32'h96696996)) lut_n1471 (.I0(x243), .I1(x244), .I2(x245), .I3(n1467), .I4(n1468), .O(n1471));
  LUT5 #(.INIT(32'hFF969600)) lut_n1472 (.I0(x249), .I1(x250), .I2(x251), .I3(n1470), .I4(n1471), .O(n1472));
  LUT3 #(.INIT(8'h96)) lut_n1473 (.I0(n1461), .I1(n1464), .I2(n1465), .O(n1473));
  LUT3 #(.INIT(8'h8E)) lut_n1474 (.I0(n1469), .I1(n1472), .I2(n1473), .O(n1474));
  LUT3 #(.INIT(8'h96)) lut_n1475 (.I0(n1448), .I1(n1456), .I2(n1457), .O(n1475));
  LUT3 #(.INIT(8'hE8)) lut_n1476 (.I0(n1466), .I1(n1474), .I2(n1475), .O(n1476));
  LUT3 #(.INIT(8'h96)) lut_n1477 (.I0(n1420), .I1(n1438), .I2(n1439), .O(n1477));
  LUT3 #(.INIT(8'h8E)) lut_n1478 (.I0(n1458), .I1(n1476), .I2(n1477), .O(n1478));
  LUT3 #(.INIT(8'h96)) lut_n1479 (.I0(n1362), .I1(n1400), .I2(n1401), .O(n1479));
  LUT3 #(.INIT(8'hE8)) lut_n1480 (.I0(n1440), .I1(n1478), .I2(n1479), .O(n1480));
  LUT2 #(.INIT(4'h6)) lut_n1481 (.I0(n1322), .I1(n1323), .O(n1481));
  LUT3 #(.INIT(8'h8E)) lut_n1482 (.I0(n1402), .I1(n1480), .I2(n1481), .O(n1482));
  LUT3 #(.INIT(8'hD4)) lut_n1483 (.I0(n1270), .I1(n1324), .I2(n1482), .O(n1483));
  LUT3 #(.INIT(8'h96)) lut_n1484 (.I0(n1000), .I1(n1158), .I2(n1269), .O(n1484));
  LUT3 #(.INIT(8'hE8)) lut_n1485 (.I0(n1270), .I1(n1483), .I2(n1484), .O(n1485));
  LUT3 #(.INIT(8'h96)) lut_n1486 (.I0(x258), .I1(x259), .I2(x260), .O(n1486));
  LUT5 #(.INIT(32'h96696996)) lut_n1487 (.I0(x249), .I1(x250), .I2(x251), .I3(n1470), .I4(n1471), .O(n1487));
  LUT5 #(.INIT(32'hFF969600)) lut_n1488 (.I0(x255), .I1(x256), .I2(x257), .I3(n1486), .I4(n1487), .O(n1488));
  LUT3 #(.INIT(8'h96)) lut_n1489 (.I0(x264), .I1(x265), .I2(x266), .O(n1489));
  LUT5 #(.INIT(32'h96696996)) lut_n1490 (.I0(x255), .I1(x256), .I2(x257), .I3(n1486), .I4(n1487), .O(n1490));
  LUT5 #(.INIT(32'hFF969600)) lut_n1491 (.I0(x261), .I1(x262), .I2(x263), .I3(n1489), .I4(n1490), .O(n1491));
  LUT3 #(.INIT(8'h96)) lut_n1492 (.I0(n1469), .I1(n1472), .I2(n1473), .O(n1492));
  LUT3 #(.INIT(8'h8E)) lut_n1493 (.I0(n1488), .I1(n1491), .I2(n1492), .O(n1493));
  LUT3 #(.INIT(8'h96)) lut_n1494 (.I0(x270), .I1(x271), .I2(x272), .O(n1494));
  LUT5 #(.INIT(32'h96696996)) lut_n1495 (.I0(x261), .I1(x262), .I2(x263), .I3(n1489), .I4(n1490), .O(n1495));
  LUT5 #(.INIT(32'hFF969600)) lut_n1496 (.I0(x267), .I1(x268), .I2(x269), .I3(n1494), .I4(n1495), .O(n1496));
  LUT3 #(.INIT(8'h96)) lut_n1497 (.I0(x276), .I1(x277), .I2(x278), .O(n1497));
  LUT5 #(.INIT(32'h96696996)) lut_n1498 (.I0(x267), .I1(x268), .I2(x269), .I3(n1494), .I4(n1495), .O(n1498));
  LUT5 #(.INIT(32'hFF969600)) lut_n1499 (.I0(x273), .I1(x274), .I2(x275), .I3(n1497), .I4(n1498), .O(n1499));
  LUT3 #(.INIT(8'h96)) lut_n1500 (.I0(n1488), .I1(n1491), .I2(n1492), .O(n1500));
  LUT3 #(.INIT(8'h8E)) lut_n1501 (.I0(n1496), .I1(n1499), .I2(n1500), .O(n1501));
  LUT3 #(.INIT(8'h96)) lut_n1502 (.I0(n1466), .I1(n1474), .I2(n1475), .O(n1502));
  LUT3 #(.INIT(8'hE8)) lut_n1503 (.I0(n1493), .I1(n1501), .I2(n1502), .O(n1503));
  LUT3 #(.INIT(8'h96)) lut_n1504 (.I0(x282), .I1(x283), .I2(x284), .O(n1504));
  LUT5 #(.INIT(32'h96696996)) lut_n1505 (.I0(x273), .I1(x274), .I2(x275), .I3(n1497), .I4(n1498), .O(n1505));
  LUT5 #(.INIT(32'hFF969600)) lut_n1506 (.I0(x279), .I1(x280), .I2(x281), .I3(n1504), .I4(n1505), .O(n1506));
  LUT3 #(.INIT(8'h96)) lut_n1507 (.I0(x288), .I1(x289), .I2(x290), .O(n1507));
  LUT5 #(.INIT(32'h96696996)) lut_n1508 (.I0(x279), .I1(x280), .I2(x281), .I3(n1504), .I4(n1505), .O(n1508));
  LUT5 #(.INIT(32'hFF969600)) lut_n1509 (.I0(x285), .I1(x286), .I2(x287), .I3(n1507), .I4(n1508), .O(n1509));
  LUT3 #(.INIT(8'h96)) lut_n1510 (.I0(n1496), .I1(n1499), .I2(n1500), .O(n1510));
  LUT3 #(.INIT(8'h8E)) lut_n1511 (.I0(n1506), .I1(n1509), .I2(n1510), .O(n1511));
  LUT3 #(.INIT(8'h96)) lut_n1512 (.I0(x294), .I1(x295), .I2(x296), .O(n1512));
  LUT5 #(.INIT(32'h96696996)) lut_n1513 (.I0(x285), .I1(x286), .I2(x287), .I3(n1507), .I4(n1508), .O(n1513));
  LUT5 #(.INIT(32'hFF969600)) lut_n1514 (.I0(x291), .I1(x292), .I2(x293), .I3(n1512), .I4(n1513), .O(n1514));
  LUT3 #(.INIT(8'h96)) lut_n1515 (.I0(x297), .I1(x298), .I2(x299), .O(n1515));
  LUT5 #(.INIT(32'h96696996)) lut_n1516 (.I0(x291), .I1(x292), .I2(x293), .I3(n1512), .I4(n1513), .O(n1516));
  LUT5 #(.INIT(32'hFF969600)) lut_n1517 (.I0(x300), .I1(x301), .I2(x302), .I3(n1515), .I4(n1516), .O(n1517));
  LUT3 #(.INIT(8'h96)) lut_n1518 (.I0(n1506), .I1(n1509), .I2(n1510), .O(n1518));
  LUT3 #(.INIT(8'h8E)) lut_n1519 (.I0(n1514), .I1(n1517), .I2(n1518), .O(n1519));
  LUT3 #(.INIT(8'h96)) lut_n1520 (.I0(n1493), .I1(n1501), .I2(n1502), .O(n1520));
  LUT3 #(.INIT(8'hE8)) lut_n1521 (.I0(n1511), .I1(n1519), .I2(n1520), .O(n1521));
  LUT3 #(.INIT(8'h96)) lut_n1522 (.I0(n1458), .I1(n1476), .I2(n1477), .O(n1522));
  LUT3 #(.INIT(8'h8E)) lut_n1523 (.I0(n1503), .I1(n1521), .I2(n1522), .O(n1523));
  LUT3 #(.INIT(8'h96)) lut_n1524 (.I0(x306), .I1(x307), .I2(x308), .O(n1524));
  LUT5 #(.INIT(32'h96696996)) lut_n1525 (.I0(x300), .I1(x301), .I2(x302), .I3(n1515), .I4(n1516), .O(n1525));
  LUT5 #(.INIT(32'hFF969600)) lut_n1526 (.I0(x303), .I1(x304), .I2(x305), .I3(n1524), .I4(n1525), .O(n1526));
  LUT3 #(.INIT(8'h96)) lut_n1527 (.I0(x312), .I1(x313), .I2(x314), .O(n1527));
  LUT5 #(.INIT(32'h96696996)) lut_n1528 (.I0(x303), .I1(x304), .I2(x305), .I3(n1524), .I4(n1525), .O(n1528));
  LUT5 #(.INIT(32'hFF969600)) lut_n1529 (.I0(x309), .I1(x310), .I2(x311), .I3(n1527), .I4(n1528), .O(n1529));
  LUT3 #(.INIT(8'h96)) lut_n1530 (.I0(n1514), .I1(n1517), .I2(n1518), .O(n1530));
  LUT3 #(.INIT(8'h8E)) lut_n1531 (.I0(n1526), .I1(n1529), .I2(n1530), .O(n1531));
  LUT3 #(.INIT(8'h96)) lut_n1532 (.I0(x318), .I1(x319), .I2(x320), .O(n1532));
  LUT5 #(.INIT(32'h96696996)) lut_n1533 (.I0(x309), .I1(x310), .I2(x311), .I3(n1527), .I4(n1528), .O(n1533));
  LUT5 #(.INIT(32'hFF969600)) lut_n1534 (.I0(x315), .I1(x316), .I2(x317), .I3(n1532), .I4(n1533), .O(n1534));
  LUT3 #(.INIT(8'h96)) lut_n1535 (.I0(x324), .I1(x325), .I2(x326), .O(n1535));
  LUT5 #(.INIT(32'h96696996)) lut_n1536 (.I0(x315), .I1(x316), .I2(x317), .I3(n1532), .I4(n1533), .O(n1536));
  LUT5 #(.INIT(32'hFF969600)) lut_n1537 (.I0(x321), .I1(x322), .I2(x323), .I3(n1535), .I4(n1536), .O(n1537));
  LUT3 #(.INIT(8'h96)) lut_n1538 (.I0(n1526), .I1(n1529), .I2(n1530), .O(n1538));
  LUT3 #(.INIT(8'h8E)) lut_n1539 (.I0(n1534), .I1(n1537), .I2(n1538), .O(n1539));
  LUT3 #(.INIT(8'h96)) lut_n1540 (.I0(n1511), .I1(n1519), .I2(n1520), .O(n1540));
  LUT3 #(.INIT(8'hE8)) lut_n1541 (.I0(n1531), .I1(n1539), .I2(n1540), .O(n1541));
  LUT3 #(.INIT(8'h96)) lut_n1542 (.I0(x330), .I1(x331), .I2(x332), .O(n1542));
  LUT5 #(.INIT(32'h96696996)) lut_n1543 (.I0(x321), .I1(x322), .I2(x323), .I3(n1535), .I4(n1536), .O(n1543));
  LUT5 #(.INIT(32'hFF969600)) lut_n1544 (.I0(x327), .I1(x328), .I2(x329), .I3(n1542), .I4(n1543), .O(n1544));
  LUT3 #(.INIT(8'h96)) lut_n1545 (.I0(x336), .I1(x337), .I2(x338), .O(n1545));
  LUT5 #(.INIT(32'h96696996)) lut_n1546 (.I0(x327), .I1(x328), .I2(x329), .I3(n1542), .I4(n1543), .O(n1546));
  LUT5 #(.INIT(32'hFF969600)) lut_n1547 (.I0(x333), .I1(x334), .I2(x335), .I3(n1545), .I4(n1546), .O(n1547));
  LUT3 #(.INIT(8'h96)) lut_n1548 (.I0(n1534), .I1(n1537), .I2(n1538), .O(n1548));
  LUT3 #(.INIT(8'h8E)) lut_n1549 (.I0(n1544), .I1(n1547), .I2(n1548), .O(n1549));
  LUT3 #(.INIT(8'h96)) lut_n1550 (.I0(x342), .I1(x343), .I2(x344), .O(n1550));
  LUT5 #(.INIT(32'h96696996)) lut_n1551 (.I0(x333), .I1(x334), .I2(x335), .I3(n1545), .I4(n1546), .O(n1551));
  LUT5 #(.INIT(32'hFF969600)) lut_n1552 (.I0(x339), .I1(x340), .I2(x341), .I3(n1550), .I4(n1551), .O(n1552));
  LUT3 #(.INIT(8'h96)) lut_n1553 (.I0(x348), .I1(x349), .I2(x350), .O(n1553));
  LUT5 #(.INIT(32'h96696996)) lut_n1554 (.I0(x339), .I1(x340), .I2(x341), .I3(n1550), .I4(n1551), .O(n1554));
  LUT5 #(.INIT(32'hFF969600)) lut_n1555 (.I0(x345), .I1(x346), .I2(x347), .I3(n1553), .I4(n1554), .O(n1555));
  LUT3 #(.INIT(8'h96)) lut_n1556 (.I0(n1544), .I1(n1547), .I2(n1548), .O(n1556));
  LUT3 #(.INIT(8'h8E)) lut_n1557 (.I0(n1552), .I1(n1555), .I2(n1556), .O(n1557));
  LUT3 #(.INIT(8'h96)) lut_n1558 (.I0(n1531), .I1(n1539), .I2(n1540), .O(n1558));
  LUT3 #(.INIT(8'hE8)) lut_n1559 (.I0(n1549), .I1(n1557), .I2(n1558), .O(n1559));
  LUT3 #(.INIT(8'h96)) lut_n1560 (.I0(n1503), .I1(n1521), .I2(n1522), .O(n1560));
  LUT3 #(.INIT(8'h8E)) lut_n1561 (.I0(n1541), .I1(n1559), .I2(n1560), .O(n1561));
  LUT3 #(.INIT(8'h96)) lut_n1562 (.I0(n1440), .I1(n1478), .I2(n1479), .O(n1562));
  LUT3 #(.INIT(8'hE8)) lut_n1563 (.I0(n1523), .I1(n1561), .I2(n1562), .O(n1563));
  LUT3 #(.INIT(8'h96)) lut_n1564 (.I0(x354), .I1(x355), .I2(x356), .O(n1564));
  LUT5 #(.INIT(32'h96696996)) lut_n1565 (.I0(x345), .I1(x346), .I2(x347), .I3(n1553), .I4(n1554), .O(n1565));
  LUT5 #(.INIT(32'hFF969600)) lut_n1566 (.I0(x351), .I1(x352), .I2(x353), .I3(n1564), .I4(n1565), .O(n1566));
  LUT3 #(.INIT(8'h96)) lut_n1567 (.I0(x360), .I1(x361), .I2(x362), .O(n1567));
  LUT5 #(.INIT(32'h96696996)) lut_n1568 (.I0(x351), .I1(x352), .I2(x353), .I3(n1564), .I4(n1565), .O(n1568));
  LUT5 #(.INIT(32'hFF969600)) lut_n1569 (.I0(x357), .I1(x358), .I2(x359), .I3(n1567), .I4(n1568), .O(n1569));
  LUT3 #(.INIT(8'h96)) lut_n1570 (.I0(n1552), .I1(n1555), .I2(n1556), .O(n1570));
  LUT3 #(.INIT(8'h8E)) lut_n1571 (.I0(n1566), .I1(n1569), .I2(n1570), .O(n1571));
  LUT3 #(.INIT(8'h96)) lut_n1572 (.I0(x366), .I1(x367), .I2(x368), .O(n1572));
  LUT5 #(.INIT(32'h96696996)) lut_n1573 (.I0(x357), .I1(x358), .I2(x359), .I3(n1567), .I4(n1568), .O(n1573));
  LUT5 #(.INIT(32'hFF969600)) lut_n1574 (.I0(x363), .I1(x364), .I2(x365), .I3(n1572), .I4(n1573), .O(n1574));
  LUT3 #(.INIT(8'h96)) lut_n1575 (.I0(x372), .I1(x373), .I2(x374), .O(n1575));
  LUT5 #(.INIT(32'h96696996)) lut_n1576 (.I0(x363), .I1(x364), .I2(x365), .I3(n1572), .I4(n1573), .O(n1576));
  LUT5 #(.INIT(32'hFF969600)) lut_n1577 (.I0(x369), .I1(x370), .I2(x371), .I3(n1575), .I4(n1576), .O(n1577));
  LUT3 #(.INIT(8'h96)) lut_n1578 (.I0(n1566), .I1(n1569), .I2(n1570), .O(n1578));
  LUT3 #(.INIT(8'h8E)) lut_n1579 (.I0(n1574), .I1(n1577), .I2(n1578), .O(n1579));
  LUT3 #(.INIT(8'h96)) lut_n1580 (.I0(n1549), .I1(n1557), .I2(n1558), .O(n1580));
  LUT3 #(.INIT(8'hE8)) lut_n1581 (.I0(n1571), .I1(n1579), .I2(n1580), .O(n1581));
  LUT3 #(.INIT(8'h96)) lut_n1582 (.I0(x378), .I1(x379), .I2(x380), .O(n1582));
  LUT5 #(.INIT(32'h96696996)) lut_n1583 (.I0(x369), .I1(x370), .I2(x371), .I3(n1575), .I4(n1576), .O(n1583));
  LUT5 #(.INIT(32'hFF969600)) lut_n1584 (.I0(x375), .I1(x376), .I2(x377), .I3(n1582), .I4(n1583), .O(n1584));
  LUT3 #(.INIT(8'h96)) lut_n1585 (.I0(x384), .I1(x385), .I2(x386), .O(n1585));
  LUT5 #(.INIT(32'h96696996)) lut_n1586 (.I0(x375), .I1(x376), .I2(x377), .I3(n1582), .I4(n1583), .O(n1586));
  LUT5 #(.INIT(32'hFF969600)) lut_n1587 (.I0(x381), .I1(x382), .I2(x383), .I3(n1585), .I4(n1586), .O(n1587));
  LUT3 #(.INIT(8'h96)) lut_n1588 (.I0(n1574), .I1(n1577), .I2(n1578), .O(n1588));
  LUT3 #(.INIT(8'h8E)) lut_n1589 (.I0(n1584), .I1(n1587), .I2(n1588), .O(n1589));
  LUT3 #(.INIT(8'h96)) lut_n1590 (.I0(x390), .I1(x391), .I2(x392), .O(n1590));
  LUT5 #(.INIT(32'h96696996)) lut_n1591 (.I0(x381), .I1(x382), .I2(x383), .I3(n1585), .I4(n1586), .O(n1591));
  LUT5 #(.INIT(32'hFF969600)) lut_n1592 (.I0(x387), .I1(x388), .I2(x389), .I3(n1590), .I4(n1591), .O(n1592));
  LUT3 #(.INIT(8'h96)) lut_n1593 (.I0(x396), .I1(x397), .I2(x398), .O(n1593));
  LUT5 #(.INIT(32'h96696996)) lut_n1594 (.I0(x387), .I1(x388), .I2(x389), .I3(n1590), .I4(n1591), .O(n1594));
  LUT5 #(.INIT(32'hFF969600)) lut_n1595 (.I0(x393), .I1(x394), .I2(x395), .I3(n1593), .I4(n1594), .O(n1595));
  LUT3 #(.INIT(8'h96)) lut_n1596 (.I0(n1584), .I1(n1587), .I2(n1588), .O(n1596));
  LUT3 #(.INIT(8'h8E)) lut_n1597 (.I0(n1592), .I1(n1595), .I2(n1596), .O(n1597));
  LUT3 #(.INIT(8'h96)) lut_n1598 (.I0(n1571), .I1(n1579), .I2(n1580), .O(n1598));
  LUT3 #(.INIT(8'hE8)) lut_n1599 (.I0(n1589), .I1(n1597), .I2(n1598), .O(n1599));
  LUT3 #(.INIT(8'h96)) lut_n1600 (.I0(n1541), .I1(n1559), .I2(n1560), .O(n1600));
  LUT3 #(.INIT(8'h8E)) lut_n1601 (.I0(n1581), .I1(n1599), .I2(n1600), .O(n1601));
  LUT3 #(.INIT(8'h96)) lut_n1602 (.I0(x402), .I1(x403), .I2(x404), .O(n1602));
  LUT5 #(.INIT(32'h96696996)) lut_n1603 (.I0(x393), .I1(x394), .I2(x395), .I3(n1593), .I4(n1594), .O(n1603));
  LUT5 #(.INIT(32'hFF969600)) lut_n1604 (.I0(x399), .I1(x400), .I2(x401), .I3(n1602), .I4(n1603), .O(n1604));
  LUT3 #(.INIT(8'h96)) lut_n1605 (.I0(x408), .I1(x409), .I2(x410), .O(n1605));
  LUT5 #(.INIT(32'h96696996)) lut_n1606 (.I0(x399), .I1(x400), .I2(x401), .I3(n1602), .I4(n1603), .O(n1606));
  LUT5 #(.INIT(32'hFF969600)) lut_n1607 (.I0(x405), .I1(x406), .I2(x407), .I3(n1605), .I4(n1606), .O(n1607));
  LUT3 #(.INIT(8'h96)) lut_n1608 (.I0(n1592), .I1(n1595), .I2(n1596), .O(n1608));
  LUT3 #(.INIT(8'h8E)) lut_n1609 (.I0(n1604), .I1(n1607), .I2(n1608), .O(n1609));
  LUT3 #(.INIT(8'h96)) lut_n1610 (.I0(x414), .I1(x415), .I2(x416), .O(n1610));
  LUT5 #(.INIT(32'h96696996)) lut_n1611 (.I0(x405), .I1(x406), .I2(x407), .I3(n1605), .I4(n1606), .O(n1611));
  LUT5 #(.INIT(32'hFF969600)) lut_n1612 (.I0(x411), .I1(x412), .I2(x413), .I3(n1610), .I4(n1611), .O(n1612));
  LUT3 #(.INIT(8'h96)) lut_n1613 (.I0(x420), .I1(x421), .I2(x422), .O(n1613));
  LUT5 #(.INIT(32'h96696996)) lut_n1614 (.I0(x411), .I1(x412), .I2(x413), .I3(n1610), .I4(n1611), .O(n1614));
  LUT5 #(.INIT(32'hFF969600)) lut_n1615 (.I0(x417), .I1(x418), .I2(x419), .I3(n1613), .I4(n1614), .O(n1615));
  LUT3 #(.INIT(8'h96)) lut_n1616 (.I0(n1604), .I1(n1607), .I2(n1608), .O(n1616));
  LUT3 #(.INIT(8'h8E)) lut_n1617 (.I0(n1612), .I1(n1615), .I2(n1616), .O(n1617));
  LUT3 #(.INIT(8'h96)) lut_n1618 (.I0(n1589), .I1(n1597), .I2(n1598), .O(n1618));
  LUT3 #(.INIT(8'hE8)) lut_n1619 (.I0(n1609), .I1(n1617), .I2(n1618), .O(n1619));
  LUT3 #(.INIT(8'h96)) lut_n1620 (.I0(x426), .I1(x427), .I2(x428), .O(n1620));
  LUT5 #(.INIT(32'h96696996)) lut_n1621 (.I0(x417), .I1(x418), .I2(x419), .I3(n1613), .I4(n1614), .O(n1621));
  LUT5 #(.INIT(32'hFF969600)) lut_n1622 (.I0(x423), .I1(x424), .I2(x425), .I3(n1620), .I4(n1621), .O(n1622));
  LUT3 #(.INIT(8'h96)) lut_n1623 (.I0(x432), .I1(x433), .I2(x434), .O(n1623));
  LUT5 #(.INIT(32'h96696996)) lut_n1624 (.I0(x423), .I1(x424), .I2(x425), .I3(n1620), .I4(n1621), .O(n1624));
  LUT5 #(.INIT(32'hFF969600)) lut_n1625 (.I0(x429), .I1(x430), .I2(x431), .I3(n1623), .I4(n1624), .O(n1625));
  LUT3 #(.INIT(8'h96)) lut_n1626 (.I0(n1612), .I1(n1615), .I2(n1616), .O(n1626));
  LUT3 #(.INIT(8'h8E)) lut_n1627 (.I0(n1622), .I1(n1625), .I2(n1626), .O(n1627));
  LUT3 #(.INIT(8'h96)) lut_n1628 (.I0(x438), .I1(x439), .I2(x440), .O(n1628));
  LUT5 #(.INIT(32'h96696996)) lut_n1629 (.I0(x429), .I1(x430), .I2(x431), .I3(n1623), .I4(n1624), .O(n1629));
  LUT5 #(.INIT(32'hFF969600)) lut_n1630 (.I0(x435), .I1(x436), .I2(x437), .I3(n1628), .I4(n1629), .O(n1630));
  LUT3 #(.INIT(8'h96)) lut_n1631 (.I0(x444), .I1(x445), .I2(x446), .O(n1631));
  LUT5 #(.INIT(32'h96696996)) lut_n1632 (.I0(x435), .I1(x436), .I2(x437), .I3(n1628), .I4(n1629), .O(n1632));
  LUT5 #(.INIT(32'hFF969600)) lut_n1633 (.I0(x441), .I1(x442), .I2(x443), .I3(n1631), .I4(n1632), .O(n1633));
  LUT3 #(.INIT(8'h96)) lut_n1634 (.I0(n1622), .I1(n1625), .I2(n1626), .O(n1634));
  LUT3 #(.INIT(8'h8E)) lut_n1635 (.I0(n1630), .I1(n1633), .I2(n1634), .O(n1635));
  LUT3 #(.INIT(8'h96)) lut_n1636 (.I0(n1609), .I1(n1617), .I2(n1618), .O(n1636));
  LUT3 #(.INIT(8'hE8)) lut_n1637 (.I0(n1627), .I1(n1635), .I2(n1636), .O(n1637));
  LUT3 #(.INIT(8'h96)) lut_n1638 (.I0(n1581), .I1(n1599), .I2(n1600), .O(n1638));
  LUT3 #(.INIT(8'h8E)) lut_n1639 (.I0(n1619), .I1(n1637), .I2(n1638), .O(n1639));
  LUT3 #(.INIT(8'h96)) lut_n1640 (.I0(n1523), .I1(n1561), .I2(n1562), .O(n1640));
  LUT3 #(.INIT(8'hE8)) lut_n1641 (.I0(n1601), .I1(n1639), .I2(n1640), .O(n1641));
  LUT3 #(.INIT(8'h96)) lut_n1642 (.I0(n1402), .I1(n1480), .I2(n1481), .O(n1642));
  LUT3 #(.INIT(8'h8E)) lut_n1643 (.I0(n1563), .I1(n1641), .I2(n1642), .O(n1643));
  LUT3 #(.INIT(8'h96)) lut_n1644 (.I0(x450), .I1(x451), .I2(x452), .O(n1644));
  LUT5 #(.INIT(32'h96696996)) lut_n1645 (.I0(x441), .I1(x442), .I2(x443), .I3(n1631), .I4(n1632), .O(n1645));
  LUT5 #(.INIT(32'hFF969600)) lut_n1646 (.I0(x447), .I1(x448), .I2(x449), .I3(n1644), .I4(n1645), .O(n1646));
  LUT3 #(.INIT(8'h96)) lut_n1647 (.I0(x456), .I1(x457), .I2(x458), .O(n1647));
  LUT5 #(.INIT(32'h96696996)) lut_n1648 (.I0(x447), .I1(x448), .I2(x449), .I3(n1644), .I4(n1645), .O(n1648));
  LUT5 #(.INIT(32'hFF969600)) lut_n1649 (.I0(x453), .I1(x454), .I2(x455), .I3(n1647), .I4(n1648), .O(n1649));
  LUT3 #(.INIT(8'h96)) lut_n1650 (.I0(n1630), .I1(n1633), .I2(n1634), .O(n1650));
  LUT3 #(.INIT(8'h8E)) lut_n1651 (.I0(n1646), .I1(n1649), .I2(n1650), .O(n1651));
  LUT3 #(.INIT(8'h96)) lut_n1652 (.I0(x462), .I1(x463), .I2(x464), .O(n1652));
  LUT5 #(.INIT(32'h96696996)) lut_n1653 (.I0(x453), .I1(x454), .I2(x455), .I3(n1647), .I4(n1648), .O(n1653));
  LUT5 #(.INIT(32'hFF969600)) lut_n1654 (.I0(x459), .I1(x460), .I2(x461), .I3(n1652), .I4(n1653), .O(n1654));
  LUT3 #(.INIT(8'h96)) lut_n1655 (.I0(x468), .I1(x469), .I2(x470), .O(n1655));
  LUT5 #(.INIT(32'h96696996)) lut_n1656 (.I0(x459), .I1(x460), .I2(x461), .I3(n1652), .I4(n1653), .O(n1656));
  LUT5 #(.INIT(32'hFF969600)) lut_n1657 (.I0(x465), .I1(x466), .I2(x467), .I3(n1655), .I4(n1656), .O(n1657));
  LUT3 #(.INIT(8'h96)) lut_n1658 (.I0(n1646), .I1(n1649), .I2(n1650), .O(n1658));
  LUT3 #(.INIT(8'h8E)) lut_n1659 (.I0(n1654), .I1(n1657), .I2(n1658), .O(n1659));
  LUT3 #(.INIT(8'h96)) lut_n1660 (.I0(n1627), .I1(n1635), .I2(n1636), .O(n1660));
  LUT3 #(.INIT(8'hE8)) lut_n1661 (.I0(n1651), .I1(n1659), .I2(n1660), .O(n1661));
  LUT3 #(.INIT(8'h96)) lut_n1662 (.I0(x474), .I1(x475), .I2(x476), .O(n1662));
  LUT5 #(.INIT(32'h96696996)) lut_n1663 (.I0(x465), .I1(x466), .I2(x467), .I3(n1655), .I4(n1656), .O(n1663));
  LUT5 #(.INIT(32'hFF969600)) lut_n1664 (.I0(x471), .I1(x472), .I2(x473), .I3(n1662), .I4(n1663), .O(n1664));
  LUT3 #(.INIT(8'h96)) lut_n1665 (.I0(x480), .I1(x481), .I2(x482), .O(n1665));
  LUT5 #(.INIT(32'h96696996)) lut_n1666 (.I0(x471), .I1(x472), .I2(x473), .I3(n1662), .I4(n1663), .O(n1666));
  LUT5 #(.INIT(32'hFF969600)) lut_n1667 (.I0(x477), .I1(x478), .I2(x479), .I3(n1665), .I4(n1666), .O(n1667));
  LUT3 #(.INIT(8'h96)) lut_n1668 (.I0(n1654), .I1(n1657), .I2(n1658), .O(n1668));
  LUT3 #(.INIT(8'h8E)) lut_n1669 (.I0(n1664), .I1(n1667), .I2(n1668), .O(n1669));
  LUT3 #(.INIT(8'h96)) lut_n1670 (.I0(x486), .I1(x487), .I2(x488), .O(n1670));
  LUT5 #(.INIT(32'h96696996)) lut_n1671 (.I0(x477), .I1(x478), .I2(x479), .I3(n1665), .I4(n1666), .O(n1671));
  LUT5 #(.INIT(32'hFF969600)) lut_n1672 (.I0(x483), .I1(x484), .I2(x485), .I3(n1670), .I4(n1671), .O(n1672));
  LUT3 #(.INIT(8'h96)) lut_n1673 (.I0(x492), .I1(x493), .I2(x494), .O(n1673));
  LUT5 #(.INIT(32'h96696996)) lut_n1674 (.I0(x483), .I1(x484), .I2(x485), .I3(n1670), .I4(n1671), .O(n1674));
  LUT5 #(.INIT(32'hFF969600)) lut_n1675 (.I0(x489), .I1(x490), .I2(x491), .I3(n1673), .I4(n1674), .O(n1675));
  LUT3 #(.INIT(8'h96)) lut_n1676 (.I0(n1664), .I1(n1667), .I2(n1668), .O(n1676));
  LUT3 #(.INIT(8'h8E)) lut_n1677 (.I0(n1672), .I1(n1675), .I2(n1676), .O(n1677));
  LUT3 #(.INIT(8'h96)) lut_n1678 (.I0(n1651), .I1(n1659), .I2(n1660), .O(n1678));
  LUT3 #(.INIT(8'hE8)) lut_n1679 (.I0(n1669), .I1(n1677), .I2(n1678), .O(n1679));
  LUT3 #(.INIT(8'h96)) lut_n1680 (.I0(n1619), .I1(n1637), .I2(n1638), .O(n1680));
  LUT3 #(.INIT(8'h8E)) lut_n1681 (.I0(n1661), .I1(n1679), .I2(n1680), .O(n1681));
  LUT3 #(.INIT(8'h96)) lut_n1682 (.I0(x498), .I1(x499), .I2(x500), .O(n1682));
  LUT5 #(.INIT(32'h96696996)) lut_n1683 (.I0(x489), .I1(x490), .I2(x491), .I3(n1673), .I4(n1674), .O(n1683));
  LUT5 #(.INIT(32'hFF969600)) lut_n1684 (.I0(x495), .I1(x496), .I2(x497), .I3(n1682), .I4(n1683), .O(n1684));
  LUT3 #(.INIT(8'h96)) lut_n1685 (.I0(x504), .I1(x505), .I2(x506), .O(n1685));
  LUT5 #(.INIT(32'h96696996)) lut_n1686 (.I0(x495), .I1(x496), .I2(x497), .I3(n1682), .I4(n1683), .O(n1686));
  LUT5 #(.INIT(32'hFF969600)) lut_n1687 (.I0(x501), .I1(x502), .I2(x503), .I3(n1685), .I4(n1686), .O(n1687));
  LUT3 #(.INIT(8'h96)) lut_n1688 (.I0(n1672), .I1(n1675), .I2(n1676), .O(n1688));
  LUT3 #(.INIT(8'h8E)) lut_n1689 (.I0(n1684), .I1(n1687), .I2(n1688), .O(n1689));
  LUT3 #(.INIT(8'h96)) lut_n1690 (.I0(x510), .I1(x511), .I2(x512), .O(n1690));
  LUT5 #(.INIT(32'h96696996)) lut_n1691 (.I0(x501), .I1(x502), .I2(x503), .I3(n1685), .I4(n1686), .O(n1691));
  LUT5 #(.INIT(32'hFF969600)) lut_n1692 (.I0(x507), .I1(x508), .I2(x509), .I3(n1690), .I4(n1691), .O(n1692));
  LUT3 #(.INIT(8'h96)) lut_n1693 (.I0(x516), .I1(x517), .I2(x518), .O(n1693));
  LUT5 #(.INIT(32'h96696996)) lut_n1694 (.I0(x507), .I1(x508), .I2(x509), .I3(n1690), .I4(n1691), .O(n1694));
  LUT5 #(.INIT(32'hFF969600)) lut_n1695 (.I0(x513), .I1(x514), .I2(x515), .I3(n1693), .I4(n1694), .O(n1695));
  LUT3 #(.INIT(8'h96)) lut_n1696 (.I0(n1684), .I1(n1687), .I2(n1688), .O(n1696));
  LUT3 #(.INIT(8'h8E)) lut_n1697 (.I0(n1692), .I1(n1695), .I2(n1696), .O(n1697));
  LUT3 #(.INIT(8'h96)) lut_n1698 (.I0(n1669), .I1(n1677), .I2(n1678), .O(n1698));
  LUT3 #(.INIT(8'hE8)) lut_n1699 (.I0(n1689), .I1(n1697), .I2(n1698), .O(n1699));
  LUT3 #(.INIT(8'h96)) lut_n1700 (.I0(x522), .I1(x523), .I2(x524), .O(n1700));
  LUT5 #(.INIT(32'h96696996)) lut_n1701 (.I0(x513), .I1(x514), .I2(x515), .I3(n1693), .I4(n1694), .O(n1701));
  LUT5 #(.INIT(32'hFF969600)) lut_n1702 (.I0(x519), .I1(x520), .I2(x521), .I3(n1700), .I4(n1701), .O(n1702));
  LUT3 #(.INIT(8'h96)) lut_n1703 (.I0(x528), .I1(x529), .I2(x530), .O(n1703));
  LUT5 #(.INIT(32'h96696996)) lut_n1704 (.I0(x519), .I1(x520), .I2(x521), .I3(n1700), .I4(n1701), .O(n1704));
  LUT5 #(.INIT(32'hFF969600)) lut_n1705 (.I0(x525), .I1(x526), .I2(x527), .I3(n1703), .I4(n1704), .O(n1705));
  LUT3 #(.INIT(8'h96)) lut_n1706 (.I0(n1692), .I1(n1695), .I2(n1696), .O(n1706));
  LUT3 #(.INIT(8'h8E)) lut_n1707 (.I0(n1702), .I1(n1705), .I2(n1706), .O(n1707));
  LUT3 #(.INIT(8'h96)) lut_n1708 (.I0(x534), .I1(x535), .I2(x536), .O(n1708));
  LUT5 #(.INIT(32'h96696996)) lut_n1709 (.I0(x525), .I1(x526), .I2(x527), .I3(n1703), .I4(n1704), .O(n1709));
  LUT5 #(.INIT(32'hFF969600)) lut_n1710 (.I0(x531), .I1(x532), .I2(x533), .I3(n1708), .I4(n1709), .O(n1710));
  LUT3 #(.INIT(8'h96)) lut_n1711 (.I0(x540), .I1(x541), .I2(x542), .O(n1711));
  LUT5 #(.INIT(32'h96696996)) lut_n1712 (.I0(x531), .I1(x532), .I2(x533), .I3(n1708), .I4(n1709), .O(n1712));
  LUT5 #(.INIT(32'hFF969600)) lut_n1713 (.I0(x537), .I1(x538), .I2(x539), .I3(n1711), .I4(n1712), .O(n1713));
  LUT3 #(.INIT(8'h96)) lut_n1714 (.I0(n1702), .I1(n1705), .I2(n1706), .O(n1714));
  LUT3 #(.INIT(8'h8E)) lut_n1715 (.I0(n1710), .I1(n1713), .I2(n1714), .O(n1715));
  LUT3 #(.INIT(8'h96)) lut_n1716 (.I0(n1689), .I1(n1697), .I2(n1698), .O(n1716));
  LUT3 #(.INIT(8'hE8)) lut_n1717 (.I0(n1707), .I1(n1715), .I2(n1716), .O(n1717));
  LUT3 #(.INIT(8'h96)) lut_n1718 (.I0(n1661), .I1(n1679), .I2(n1680), .O(n1718));
  LUT3 #(.INIT(8'h8E)) lut_n1719 (.I0(n1699), .I1(n1717), .I2(n1718), .O(n1719));
  LUT3 #(.INIT(8'h96)) lut_n1720 (.I0(n1601), .I1(n1639), .I2(n1640), .O(n1720));
  LUT3 #(.INIT(8'hE8)) lut_n1721 (.I0(n1681), .I1(n1719), .I2(n1720), .O(n1721));
  LUT3 #(.INIT(8'h96)) lut_n1722 (.I0(x546), .I1(x547), .I2(x548), .O(n1722));
  LUT5 #(.INIT(32'h96696996)) lut_n1723 (.I0(x537), .I1(x538), .I2(x539), .I3(n1711), .I4(n1712), .O(n1723));
  LUT5 #(.INIT(32'hFF969600)) lut_n1724 (.I0(x543), .I1(x544), .I2(x545), .I3(n1722), .I4(n1723), .O(n1724));
  LUT3 #(.INIT(8'h96)) lut_n1725 (.I0(x552), .I1(x553), .I2(x554), .O(n1725));
  LUT5 #(.INIT(32'h96696996)) lut_n1726 (.I0(x543), .I1(x544), .I2(x545), .I3(n1722), .I4(n1723), .O(n1726));
  LUT5 #(.INIT(32'hFF969600)) lut_n1727 (.I0(x549), .I1(x550), .I2(x551), .I3(n1725), .I4(n1726), .O(n1727));
  LUT3 #(.INIT(8'h96)) lut_n1728 (.I0(n1710), .I1(n1713), .I2(n1714), .O(n1728));
  LUT3 #(.INIT(8'h8E)) lut_n1729 (.I0(n1724), .I1(n1727), .I2(n1728), .O(n1729));
  LUT3 #(.INIT(8'h96)) lut_n1730 (.I0(x558), .I1(x559), .I2(x560), .O(n1730));
  LUT5 #(.INIT(32'h96696996)) lut_n1731 (.I0(x549), .I1(x550), .I2(x551), .I3(n1725), .I4(n1726), .O(n1731));
  LUT5 #(.INIT(32'hFF969600)) lut_n1732 (.I0(x555), .I1(x556), .I2(x557), .I3(n1730), .I4(n1731), .O(n1732));
  LUT3 #(.INIT(8'h96)) lut_n1733 (.I0(x564), .I1(x565), .I2(x566), .O(n1733));
  LUT5 #(.INIT(32'h96696996)) lut_n1734 (.I0(x555), .I1(x556), .I2(x557), .I3(n1730), .I4(n1731), .O(n1734));
  LUT5 #(.INIT(32'hFF969600)) lut_n1735 (.I0(x561), .I1(x562), .I2(x563), .I3(n1733), .I4(n1734), .O(n1735));
  LUT3 #(.INIT(8'h96)) lut_n1736 (.I0(n1724), .I1(n1727), .I2(n1728), .O(n1736));
  LUT3 #(.INIT(8'h8E)) lut_n1737 (.I0(n1732), .I1(n1735), .I2(n1736), .O(n1737));
  LUT3 #(.INIT(8'h96)) lut_n1738 (.I0(n1707), .I1(n1715), .I2(n1716), .O(n1738));
  LUT3 #(.INIT(8'hE8)) lut_n1739 (.I0(n1729), .I1(n1737), .I2(n1738), .O(n1739));
  LUT3 #(.INIT(8'h96)) lut_n1740 (.I0(x570), .I1(x571), .I2(x572), .O(n1740));
  LUT5 #(.INIT(32'h96696996)) lut_n1741 (.I0(x561), .I1(x562), .I2(x563), .I3(n1733), .I4(n1734), .O(n1741));
  LUT5 #(.INIT(32'hFF969600)) lut_n1742 (.I0(x567), .I1(x568), .I2(x569), .I3(n1740), .I4(n1741), .O(n1742));
  LUT3 #(.INIT(8'h96)) lut_n1743 (.I0(x576), .I1(x577), .I2(x578), .O(n1743));
  LUT5 #(.INIT(32'h96696996)) lut_n1744 (.I0(x567), .I1(x568), .I2(x569), .I3(n1740), .I4(n1741), .O(n1744));
  LUT5 #(.INIT(32'hFF969600)) lut_n1745 (.I0(x573), .I1(x574), .I2(x575), .I3(n1743), .I4(n1744), .O(n1745));
  LUT3 #(.INIT(8'h96)) lut_n1746 (.I0(n1732), .I1(n1735), .I2(n1736), .O(n1746));
  LUT3 #(.INIT(8'h8E)) lut_n1747 (.I0(n1742), .I1(n1745), .I2(n1746), .O(n1747));
  LUT3 #(.INIT(8'h96)) lut_n1748 (.I0(x582), .I1(x583), .I2(x584), .O(n1748));
  LUT5 #(.INIT(32'h96696996)) lut_n1749 (.I0(x573), .I1(x574), .I2(x575), .I3(n1743), .I4(n1744), .O(n1749));
  LUT5 #(.INIT(32'hFF969600)) lut_n1750 (.I0(x579), .I1(x580), .I2(x581), .I3(n1748), .I4(n1749), .O(n1750));
  LUT3 #(.INIT(8'h96)) lut_n1751 (.I0(x588), .I1(x589), .I2(x590), .O(n1751));
  LUT5 #(.INIT(32'h96696996)) lut_n1752 (.I0(x579), .I1(x580), .I2(x581), .I3(n1748), .I4(n1749), .O(n1752));
  LUT5 #(.INIT(32'hFF969600)) lut_n1753 (.I0(x585), .I1(x586), .I2(x587), .I3(n1751), .I4(n1752), .O(n1753));
  LUT3 #(.INIT(8'h96)) lut_n1754 (.I0(n1742), .I1(n1745), .I2(n1746), .O(n1754));
  LUT3 #(.INIT(8'h8E)) lut_n1755 (.I0(n1750), .I1(n1753), .I2(n1754), .O(n1755));
  LUT3 #(.INIT(8'h96)) lut_n1756 (.I0(n1729), .I1(n1737), .I2(n1738), .O(n1756));
  LUT3 #(.INIT(8'hE8)) lut_n1757 (.I0(n1747), .I1(n1755), .I2(n1756), .O(n1757));
  LUT3 #(.INIT(8'h96)) lut_n1758 (.I0(n1699), .I1(n1717), .I2(n1718), .O(n1758));
  LUT3 #(.INIT(8'h8E)) lut_n1759 (.I0(n1739), .I1(n1757), .I2(n1758), .O(n1759));
  LUT3 #(.INIT(8'h96)) lut_n1760 (.I0(x594), .I1(x595), .I2(x596), .O(n1760));
  LUT5 #(.INIT(32'h96696996)) lut_n1761 (.I0(x585), .I1(x586), .I2(x587), .I3(n1751), .I4(n1752), .O(n1761));
  LUT5 #(.INIT(32'hFF969600)) lut_n1762 (.I0(x591), .I1(x592), .I2(x593), .I3(n1760), .I4(n1761), .O(n1762));
  LUT3 #(.INIT(8'h96)) lut_n1763 (.I0(x600), .I1(x601), .I2(x602), .O(n1763));
  LUT5 #(.INIT(32'h96696996)) lut_n1764 (.I0(x591), .I1(x592), .I2(x593), .I3(n1760), .I4(n1761), .O(n1764));
  LUT5 #(.INIT(32'hFF969600)) lut_n1765 (.I0(x597), .I1(x598), .I2(x599), .I3(n1763), .I4(n1764), .O(n1765));
  LUT3 #(.INIT(8'h96)) lut_n1766 (.I0(n1750), .I1(n1753), .I2(n1754), .O(n1766));
  LUT3 #(.INIT(8'h8E)) lut_n1767 (.I0(n1762), .I1(n1765), .I2(n1766), .O(n1767));
  LUT3 #(.INIT(8'h96)) lut_n1768 (.I0(x606), .I1(x607), .I2(x608), .O(n1768));
  LUT5 #(.INIT(32'h96696996)) lut_n1769 (.I0(x597), .I1(x598), .I2(x599), .I3(n1763), .I4(n1764), .O(n1769));
  LUT5 #(.INIT(32'hFF969600)) lut_n1770 (.I0(x603), .I1(x604), .I2(x605), .I3(n1768), .I4(n1769), .O(n1770));
  LUT3 #(.INIT(8'h96)) lut_n1771 (.I0(x612), .I1(x613), .I2(x614), .O(n1771));
  LUT5 #(.INIT(32'h96696996)) lut_n1772 (.I0(x603), .I1(x604), .I2(x605), .I3(n1768), .I4(n1769), .O(n1772));
  LUT5 #(.INIT(32'hFF969600)) lut_n1773 (.I0(x609), .I1(x610), .I2(x611), .I3(n1771), .I4(n1772), .O(n1773));
  LUT3 #(.INIT(8'h96)) lut_n1774 (.I0(n1762), .I1(n1765), .I2(n1766), .O(n1774));
  LUT3 #(.INIT(8'h8E)) lut_n1775 (.I0(n1770), .I1(n1773), .I2(n1774), .O(n1775));
  LUT3 #(.INIT(8'h96)) lut_n1776 (.I0(n1747), .I1(n1755), .I2(n1756), .O(n1776));
  LUT3 #(.INIT(8'hE8)) lut_n1777 (.I0(n1767), .I1(n1775), .I2(n1776), .O(n1777));
  LUT3 #(.INIT(8'h96)) lut_n1778 (.I0(x618), .I1(x619), .I2(x620), .O(n1778));
  LUT5 #(.INIT(32'h96696996)) lut_n1779 (.I0(x609), .I1(x610), .I2(x611), .I3(n1771), .I4(n1772), .O(n1779));
  LUT5 #(.INIT(32'hFF969600)) lut_n1780 (.I0(x615), .I1(x616), .I2(x617), .I3(n1778), .I4(n1779), .O(n1780));
  LUT3 #(.INIT(8'h96)) lut_n1781 (.I0(x624), .I1(x625), .I2(x626), .O(n1781));
  LUT5 #(.INIT(32'h96696996)) lut_n1782 (.I0(x615), .I1(x616), .I2(x617), .I3(n1778), .I4(n1779), .O(n1782));
  LUT5 #(.INIT(32'hFF969600)) lut_n1783 (.I0(x621), .I1(x622), .I2(x623), .I3(n1781), .I4(n1782), .O(n1783));
  LUT3 #(.INIT(8'h96)) lut_n1784 (.I0(n1770), .I1(n1773), .I2(n1774), .O(n1784));
  LUT3 #(.INIT(8'h8E)) lut_n1785 (.I0(n1780), .I1(n1783), .I2(n1784), .O(n1785));
  LUT3 #(.INIT(8'h96)) lut_n1786 (.I0(x630), .I1(x631), .I2(x632), .O(n1786));
  LUT5 #(.INIT(32'h96696996)) lut_n1787 (.I0(x621), .I1(x622), .I2(x623), .I3(n1781), .I4(n1782), .O(n1787));
  LUT5 #(.INIT(32'hFF969600)) lut_n1788 (.I0(x627), .I1(x628), .I2(x629), .I3(n1786), .I4(n1787), .O(n1788));
  LUT3 #(.INIT(8'h96)) lut_n1789 (.I0(x636), .I1(x637), .I2(x638), .O(n1789));
  LUT5 #(.INIT(32'h96696996)) lut_n1790 (.I0(x627), .I1(x628), .I2(x629), .I3(n1786), .I4(n1787), .O(n1790));
  LUT5 #(.INIT(32'hFF969600)) lut_n1791 (.I0(x633), .I1(x634), .I2(x635), .I3(n1789), .I4(n1790), .O(n1791));
  LUT3 #(.INIT(8'h96)) lut_n1792 (.I0(n1780), .I1(n1783), .I2(n1784), .O(n1792));
  LUT3 #(.INIT(8'h8E)) lut_n1793 (.I0(n1788), .I1(n1791), .I2(n1792), .O(n1793));
  LUT3 #(.INIT(8'h96)) lut_n1794 (.I0(n1767), .I1(n1775), .I2(n1776), .O(n1794));
  LUT3 #(.INIT(8'hE8)) lut_n1795 (.I0(n1785), .I1(n1793), .I2(n1794), .O(n1795));
  LUT3 #(.INIT(8'h96)) lut_n1796 (.I0(n1739), .I1(n1757), .I2(n1758), .O(n1796));
  LUT3 #(.INIT(8'h8E)) lut_n1797 (.I0(n1777), .I1(n1795), .I2(n1796), .O(n1797));
  LUT3 #(.INIT(8'h96)) lut_n1798 (.I0(n1681), .I1(n1719), .I2(n1720), .O(n1798));
  LUT3 #(.INIT(8'hE8)) lut_n1799 (.I0(n1759), .I1(n1797), .I2(n1798), .O(n1799));
  LUT3 #(.INIT(8'h96)) lut_n1800 (.I0(n1563), .I1(n1641), .I2(n1642), .O(n1800));
  LUT3 #(.INIT(8'h8E)) lut_n1801 (.I0(n1721), .I1(n1799), .I2(n1800), .O(n1801));
  LUT3 #(.INIT(8'h96)) lut_n1802 (.I0(n1270), .I1(n1324), .I2(n1482), .O(n1802));
  LUT3 #(.INIT(8'h8E)) lut_n1803 (.I0(n1643), .I1(n1801), .I2(n1802), .O(n1803));
  LUT3 #(.INIT(8'h96)) lut_n1804 (.I0(x642), .I1(x643), .I2(x644), .O(n1804));
  LUT5 #(.INIT(32'h96696996)) lut_n1805 (.I0(x633), .I1(x634), .I2(x635), .I3(n1789), .I4(n1790), .O(n1805));
  LUT5 #(.INIT(32'hFF969600)) lut_n1806 (.I0(x639), .I1(x640), .I2(x641), .I3(n1804), .I4(n1805), .O(n1806));
  LUT3 #(.INIT(8'h96)) lut_n1807 (.I0(x648), .I1(x649), .I2(x650), .O(n1807));
  LUT5 #(.INIT(32'h96696996)) lut_n1808 (.I0(x639), .I1(x640), .I2(x641), .I3(n1804), .I4(n1805), .O(n1808));
  LUT5 #(.INIT(32'hFF969600)) lut_n1809 (.I0(x645), .I1(x646), .I2(x647), .I3(n1807), .I4(n1808), .O(n1809));
  LUT3 #(.INIT(8'h96)) lut_n1810 (.I0(n1788), .I1(n1791), .I2(n1792), .O(n1810));
  LUT3 #(.INIT(8'h8E)) lut_n1811 (.I0(n1806), .I1(n1809), .I2(n1810), .O(n1811));
  LUT3 #(.INIT(8'h96)) lut_n1812 (.I0(x654), .I1(x655), .I2(x656), .O(n1812));
  LUT5 #(.INIT(32'h96696996)) lut_n1813 (.I0(x645), .I1(x646), .I2(x647), .I3(n1807), .I4(n1808), .O(n1813));
  LUT5 #(.INIT(32'hFF969600)) lut_n1814 (.I0(x651), .I1(x652), .I2(x653), .I3(n1812), .I4(n1813), .O(n1814));
  LUT3 #(.INIT(8'h96)) lut_n1815 (.I0(x660), .I1(x661), .I2(x662), .O(n1815));
  LUT5 #(.INIT(32'h96696996)) lut_n1816 (.I0(x651), .I1(x652), .I2(x653), .I3(n1812), .I4(n1813), .O(n1816));
  LUT5 #(.INIT(32'hFF969600)) lut_n1817 (.I0(x657), .I1(x658), .I2(x659), .I3(n1815), .I4(n1816), .O(n1817));
  LUT3 #(.INIT(8'h96)) lut_n1818 (.I0(n1806), .I1(n1809), .I2(n1810), .O(n1818));
  LUT3 #(.INIT(8'h8E)) lut_n1819 (.I0(n1814), .I1(n1817), .I2(n1818), .O(n1819));
  LUT3 #(.INIT(8'h96)) lut_n1820 (.I0(n1785), .I1(n1793), .I2(n1794), .O(n1820));
  LUT3 #(.INIT(8'hE8)) lut_n1821 (.I0(n1811), .I1(n1819), .I2(n1820), .O(n1821));
  LUT3 #(.INIT(8'h96)) lut_n1822 (.I0(x666), .I1(x667), .I2(x668), .O(n1822));
  LUT5 #(.INIT(32'h96696996)) lut_n1823 (.I0(x657), .I1(x658), .I2(x659), .I3(n1815), .I4(n1816), .O(n1823));
  LUT5 #(.INIT(32'hFF969600)) lut_n1824 (.I0(x663), .I1(x664), .I2(x665), .I3(n1822), .I4(n1823), .O(n1824));
  LUT3 #(.INIT(8'h96)) lut_n1825 (.I0(x672), .I1(x673), .I2(x674), .O(n1825));
  LUT5 #(.INIT(32'h96696996)) lut_n1826 (.I0(x663), .I1(x664), .I2(x665), .I3(n1822), .I4(n1823), .O(n1826));
  LUT5 #(.INIT(32'hFF969600)) lut_n1827 (.I0(x669), .I1(x670), .I2(x671), .I3(n1825), .I4(n1826), .O(n1827));
  LUT3 #(.INIT(8'h96)) lut_n1828 (.I0(n1814), .I1(n1817), .I2(n1818), .O(n1828));
  LUT3 #(.INIT(8'h8E)) lut_n1829 (.I0(n1824), .I1(n1827), .I2(n1828), .O(n1829));
  LUT3 #(.INIT(8'h96)) lut_n1830 (.I0(x678), .I1(x679), .I2(x680), .O(n1830));
  LUT5 #(.INIT(32'h96696996)) lut_n1831 (.I0(x669), .I1(x670), .I2(x671), .I3(n1825), .I4(n1826), .O(n1831));
  LUT5 #(.INIT(32'hFF969600)) lut_n1832 (.I0(x675), .I1(x676), .I2(x677), .I3(n1830), .I4(n1831), .O(n1832));
  LUT3 #(.INIT(8'h96)) lut_n1833 (.I0(x684), .I1(x685), .I2(x686), .O(n1833));
  LUT5 #(.INIT(32'h96696996)) lut_n1834 (.I0(x675), .I1(x676), .I2(x677), .I3(n1830), .I4(n1831), .O(n1834));
  LUT5 #(.INIT(32'hFF969600)) lut_n1835 (.I0(x681), .I1(x682), .I2(x683), .I3(n1833), .I4(n1834), .O(n1835));
  LUT3 #(.INIT(8'h96)) lut_n1836 (.I0(n1824), .I1(n1827), .I2(n1828), .O(n1836));
  LUT3 #(.INIT(8'h8E)) lut_n1837 (.I0(n1832), .I1(n1835), .I2(n1836), .O(n1837));
  LUT3 #(.INIT(8'h96)) lut_n1838 (.I0(n1811), .I1(n1819), .I2(n1820), .O(n1838));
  LUT3 #(.INIT(8'hE8)) lut_n1839 (.I0(n1829), .I1(n1837), .I2(n1838), .O(n1839));
  LUT3 #(.INIT(8'h96)) lut_n1840 (.I0(n1777), .I1(n1795), .I2(n1796), .O(n1840));
  LUT3 #(.INIT(8'h8E)) lut_n1841 (.I0(n1821), .I1(n1839), .I2(n1840), .O(n1841));
  LUT3 #(.INIT(8'h96)) lut_n1842 (.I0(x690), .I1(x691), .I2(x692), .O(n1842));
  LUT5 #(.INIT(32'h96696996)) lut_n1843 (.I0(x681), .I1(x682), .I2(x683), .I3(n1833), .I4(n1834), .O(n1843));
  LUT5 #(.INIT(32'hFF969600)) lut_n1844 (.I0(x687), .I1(x688), .I2(x689), .I3(n1842), .I4(n1843), .O(n1844));
  LUT3 #(.INIT(8'h96)) lut_n1845 (.I0(x696), .I1(x697), .I2(x698), .O(n1845));
  LUT5 #(.INIT(32'h96696996)) lut_n1846 (.I0(x687), .I1(x688), .I2(x689), .I3(n1842), .I4(n1843), .O(n1846));
  LUT5 #(.INIT(32'hFF969600)) lut_n1847 (.I0(x693), .I1(x694), .I2(x695), .I3(n1845), .I4(n1846), .O(n1847));
  LUT3 #(.INIT(8'h96)) lut_n1848 (.I0(n1832), .I1(n1835), .I2(n1836), .O(n1848));
  LUT3 #(.INIT(8'h8E)) lut_n1849 (.I0(n1844), .I1(n1847), .I2(n1848), .O(n1849));
  LUT2 #(.INIT(4'h6)) lut_n1850 (.I0(x699), .I1(x700), .O(n1850));
  LUT5 #(.INIT(32'h96696996)) lut_n1851 (.I0(x693), .I1(x694), .I2(x695), .I3(n1845), .I4(n1846), .O(n1851));
  LUT3 #(.INIT(8'h96)) lut_n1852 (.I0(n1844), .I1(n1847), .I2(n1848), .O(n1852));
  LUT3 #(.INIT(8'h96)) lut_n1853 (.I0(n1829), .I1(n1837), .I2(n1838), .O(n1853));
  LUT3 #(.INIT(8'h96)) lut_n1854 (.I0(n1821), .I1(n1839), .I2(n1840), .O(n1854));
  LUT6 #(.INIT(64'h04005D5500000000)) lut_n1855 (.I0(n1849), .I1(n1850), .I2(n1851), .I3(n1852), .I4(n1853), .I5(n1854), .O(n1855));
  LUT3 #(.INIT(8'h96)) lut_n1856 (.I0(n1759), .I1(n1797), .I2(n1798), .O(n1856));
  LUT3 #(.INIT(8'h96)) lut_n1857 (.I0(n1721), .I1(n1799), .I2(n1800), .O(n1857));
  LUT6 #(.INIT(64'hDB55A2AA00004500)) lut_n1858 (.I0(n1849), .I1(n1850), .I2(n1851), .I3(n1852), .I4(n1853), .I5(n1854), .O(n1858));
  LUT3 #(.INIT(8'h96)) lut_n1859 (.I0(n1643), .I1(n1801), .I2(n1802), .O(n1859));
  LUT6 #(.INIT(64'hFFFFFFDF4D000400)) lut_n1860 (.I0(n1841), .I1(n1855), .I2(n1856), .I3(n1857), .I4(n1858), .I5(n1859), .O(n1860));
  LUT5 #(.INIT(32'h9600FF96)) lut_n1861 (.I0(n1270), .I1(n1483), .I2(n1484), .I3(n1803), .I4(n1860), .O(n1861));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1862 (.I0(n1000), .I1(n1158), .I2(n1269), .I3(n1485), .I4(n1861), .O(n1862));
  assign y0 = n1862;
endmodule
