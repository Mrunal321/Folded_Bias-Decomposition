`timescale 1ns/1ps
`default_nettype none

module tb_top;
  // 1015-bit input vector
  reg  [1014:0] x = 1015'b0;
  wire       y0;
  reg  [63:0] idx;

  // DUT instantiation
  top dut (
    .x0(x[0]), .x1(x[1]), .x2(x[2]), .x3(x[3]), .x4(x[4]), .x5(x[5]), .x6(x[6]), .x7(x[7]), .x8(x[8]), .x9(x[9]), .x10(x[10]), .x11(x[11]), .x12(x[12]), .x13(x[13]), .x14(x[14]), .x15(x[15]), .x16(x[16]), .x17(x[17]), .x18(x[18]), .x19(x[19]), .x20(x[20]), .x21(x[21]), .x22(x[22]), .x23(x[23]), .x24(x[24]), .x25(x[25]), .x26(x[26]), .x27(x[27]), .x28(x[28]), .x29(x[29]), .x30(x[30]), .x31(x[31]), .x32(x[32]), .x33(x[33]), .x34(x[34]), .x35(x[35]), .x36(x[36]), .x37(x[37]), .x38(x[38]), .x39(x[39]), .x40(x[40]), .x41(x[41]), .x42(x[42]), .x43(x[43]), .x44(x[44]), .x45(x[45]), .x46(x[46]), .x47(x[47]), .x48(x[48]), .x49(x[49]), .x50(x[50]), .x51(x[51]), .x52(x[52]), .x53(x[53]), .x54(x[54]), .x55(x[55]), .x56(x[56]), .x57(x[57]), .x58(x[58]), .x59(x[59]), .x60(x[60]), .x61(x[61]), .x62(x[62]), .x63(x[63]), .x64(x[64]), .x65(x[65]), .x66(x[66]), .x67(x[67]), .x68(x[68]), .x69(x[69]), .x70(x[70]), .x71(x[71]), .x72(x[72]), .x73(x[73]), .x74(x[74]), .x75(x[75]), .x76(x[76]), .x77(x[77]), .x78(x[78]), .x79(x[79]), .x80(x[80]), .x81(x[81]), .x82(x[82]), .x83(x[83]), .x84(x[84]), .x85(x[85]), .x86(x[86]), .x87(x[87]), .x88(x[88]), .x89(x[89]), .x90(x[90]), .x91(x[91]), .x92(x[92]), .x93(x[93]), .x94(x[94]), .x95(x[95]), .x96(x[96]), .x97(x[97]), .x98(x[98]), .x99(x[99]), .x100(x[100]), .x101(x[101]), .x102(x[102]), .x103(x[103]), .x104(x[104]), .x105(x[105]), .x106(x[106]), .x107(x[107]), .x108(x[108]), .x109(x[109]), .x110(x[110]), .x111(x[111]), .x112(x[112]), .x113(x[113]), .x114(x[114]), .x115(x[115]), .x116(x[116]), .x117(x[117]), .x118(x[118]), .x119(x[119]), .x120(x[120]), .x121(x[121]), .x122(x[122]), .x123(x[123]), .x124(x[124]), .x125(x[125]), .x126(x[126]), .x127(x[127]), .x128(x[128]), .x129(x[129]), .x130(x[130]), .x131(x[131]), .x132(x[132]), .x133(x[133]), .x134(x[134]), .x135(x[135]), .x136(x[136]), .x137(x[137]), .x138(x[138]), .x139(x[139]), .x140(x[140]), .x141(x[141]), .x142(x[142]), .x143(x[143]), .x144(x[144]), .x145(x[145]), .x146(x[146]), .x147(x[147]), .x148(x[148]), .x149(x[149]), .x150(x[150]), .x151(x[151]), .x152(x[152]), .x153(x[153]), .x154(x[154]), .x155(x[155]), .x156(x[156]), .x157(x[157]), .x158(x[158]), .x159(x[159]), .x160(x[160]), .x161(x[161]), .x162(x[162]), .x163(x[163]), .x164(x[164]), .x165(x[165]), .x166(x[166]), .x167(x[167]), .x168(x[168]), .x169(x[169]), .x170(x[170]), .x171(x[171]), .x172(x[172]), .x173(x[173]), .x174(x[174]), .x175(x[175]), .x176(x[176]), .x177(x[177]), .x178(x[178]), .x179(x[179]), .x180(x[180]), .x181(x[181]), .x182(x[182]), .x183(x[183]), .x184(x[184]), .x185(x[185]), .x186(x[186]), .x187(x[187]), .x188(x[188]), .x189(x[189]), .x190(x[190]), .x191(x[191]), .x192(x[192]), .x193(x[193]), .x194(x[194]), .x195(x[195]), .x196(x[196]), .x197(x[197]), .x198(x[198]), .x199(x[199]), .x200(x[200]), .x201(x[201]), .x202(x[202]), .x203(x[203]), .x204(x[204]), .x205(x[205]), .x206(x[206]), .x207(x[207]), .x208(x[208]), .x209(x[209]), .x210(x[210]), .x211(x[211]), .x212(x[212]), .x213(x[213]), .x214(x[214]), .x215(x[215]), .x216(x[216]), .x217(x[217]), .x218(x[218]), .x219(x[219]), .x220(x[220]), .x221(x[221]), .x222(x[222]), .x223(x[223]), .x224(x[224]), .x225(x[225]), .x226(x[226]), .x227(x[227]), .x228(x[228]), .x229(x[229]), .x230(x[230]), .x231(x[231]), .x232(x[232]), .x233(x[233]), .x234(x[234]), .x235(x[235]), .x236(x[236]), .x237(x[237]), .x238(x[238]), .x239(x[239]), .x240(x[240]), .x241(x[241]), .x242(x[242]), .x243(x[243]), .x244(x[244]), .x245(x[245]), .x246(x[246]), .x247(x[247]), .x248(x[248]), .x249(x[249]), .x250(x[250]), .x251(x[251]), .x252(x[252]), .x253(x[253]), .x254(x[254]), .x255(x[255]), .x256(x[256]), .x257(x[257]), .x258(x[258]), .x259(x[259]), .x260(x[260]), .x261(x[261]), .x262(x[262]), .x263(x[263]), .x264(x[264]), .x265(x[265]), .x266(x[266]), .x267(x[267]), .x268(x[268]), .x269(x[269]), .x270(x[270]), .x271(x[271]), .x272(x[272]), .x273(x[273]), .x274(x[274]), .x275(x[275]), .x276(x[276]), .x277(x[277]), .x278(x[278]), .x279(x[279]), .x280(x[280]), .x281(x[281]), .x282(x[282]), .x283(x[283]), .x284(x[284]), .x285(x[285]), .x286(x[286]), .x287(x[287]), .x288(x[288]), .x289(x[289]), .x290(x[290]), .x291(x[291]), .x292(x[292]), .x293(x[293]), .x294(x[294]), .x295(x[295]), .x296(x[296]), .x297(x[297]), .x298(x[298]), .x299(x[299]), .x300(x[300]), .x301(x[301]), .x302(x[302]), .x303(x[303]), .x304(x[304]), .x305(x[305]), .x306(x[306]), .x307(x[307]), .x308(x[308]), .x309(x[309]), .x310(x[310]), .x311(x[311]), .x312(x[312]), .x313(x[313]), .x314(x[314]), .x315(x[315]), .x316(x[316]), .x317(x[317]), .x318(x[318]), .x319(x[319]), .x320(x[320]), .x321(x[321]), .x322(x[322]), .x323(x[323]), .x324(x[324]), .x325(x[325]), .x326(x[326]), .x327(x[327]), .x328(x[328]), .x329(x[329]), .x330(x[330]), .x331(x[331]), .x332(x[332]), .x333(x[333]), .x334(x[334]), .x335(x[335]), .x336(x[336]), .x337(x[337]), .x338(x[338]), .x339(x[339]), .x340(x[340]), .x341(x[341]), .x342(x[342]), .x343(x[343]), .x344(x[344]), .x345(x[345]), .x346(x[346]), .x347(x[347]), .x348(x[348]), .x349(x[349]), .x350(x[350]), .x351(x[351]), .x352(x[352]), .x353(x[353]), .x354(x[354]), .x355(x[355]), .x356(x[356]), .x357(x[357]), .x358(x[358]), .x359(x[359]), .x360(x[360]), .x361(x[361]), .x362(x[362]), .x363(x[363]), .x364(x[364]), .x365(x[365]), .x366(x[366]), .x367(x[367]), .x368(x[368]), .x369(x[369]), .x370(x[370]), .x371(x[371]), .x372(x[372]), .x373(x[373]), .x374(x[374]), .x375(x[375]), .x376(x[376]), .x377(x[377]), .x378(x[378]), .x379(x[379]), .x380(x[380]), .x381(x[381]), .x382(x[382]), .x383(x[383]), .x384(x[384]), .x385(x[385]), .x386(x[386]), .x387(x[387]), .x388(x[388]), .x389(x[389]), .x390(x[390]), .x391(x[391]), .x392(x[392]), .x393(x[393]), .x394(x[394]), .x395(x[395]), .x396(x[396]), .x397(x[397]), .x398(x[398]), .x399(x[399]), .x400(x[400]), .x401(x[401]), .x402(x[402]), .x403(x[403]), .x404(x[404]), .x405(x[405]), .x406(x[406]), .x407(x[407]), .x408(x[408]), .x409(x[409]), .x410(x[410]), .x411(x[411]), .x412(x[412]), .x413(x[413]), .x414(x[414]), .x415(x[415]), .x416(x[416]), .x417(x[417]), .x418(x[418]), .x419(x[419]), .x420(x[420]), .x421(x[421]), .x422(x[422]), .x423(x[423]), .x424(x[424]), .x425(x[425]), .x426(x[426]), .x427(x[427]), .x428(x[428]), .x429(x[429]), .x430(x[430]), .x431(x[431]), .x432(x[432]), .x433(x[433]), .x434(x[434]), .x435(x[435]), .x436(x[436]), .x437(x[437]), .x438(x[438]), .x439(x[439]), .x440(x[440]), .x441(x[441]), .x442(x[442]), .x443(x[443]), .x444(x[444]), .x445(x[445]), .x446(x[446]), .x447(x[447]), .x448(x[448]), .x449(x[449]), .x450(x[450]), .x451(x[451]), .x452(x[452]), .x453(x[453]), .x454(x[454]), .x455(x[455]), .x456(x[456]), .x457(x[457]), .x458(x[458]), .x459(x[459]), .x460(x[460]), .x461(x[461]), .x462(x[462]), .x463(x[463]), .x464(x[464]), .x465(x[465]), .x466(x[466]), .x467(x[467]), .x468(x[468]), .x469(x[469]), .x470(x[470]), .x471(x[471]), .x472(x[472]), .x473(x[473]), .x474(x[474]), .x475(x[475]), .x476(x[476]), .x477(x[477]), .x478(x[478]), .x479(x[479]), .x480(x[480]), .x481(x[481]), .x482(x[482]), .x483(x[483]), .x484(x[484]), .x485(x[485]), .x486(x[486]), .x487(x[487]), .x488(x[488]), .x489(x[489]), .x490(x[490]), .x491(x[491]), .x492(x[492]), .x493(x[493]), .x494(x[494]), .x495(x[495]), .x496(x[496]), .x497(x[497]), .x498(x[498]), .x499(x[499]), .x500(x[500]), .x501(x[501]), .x502(x[502]), .x503(x[503]), .x504(x[504]), .x505(x[505]), .x506(x[506]), .x507(x[507]), .x508(x[508]), .x509(x[509]), .x510(x[510]), .x511(x[511]), .x512(x[512]), .x513(x[513]), .x514(x[514]), .x515(x[515]), .x516(x[516]), .x517(x[517]), .x518(x[518]), .x519(x[519]), .x520(x[520]), .x521(x[521]), .x522(x[522]), .x523(x[523]), .x524(x[524]), .x525(x[525]), .x526(x[526]), .x527(x[527]), .x528(x[528]), .x529(x[529]), .x530(x[530]), .x531(x[531]), .x532(x[532]), .x533(x[533]), .x534(x[534]), .x535(x[535]), .x536(x[536]), .x537(x[537]), .x538(x[538]), .x539(x[539]), .x540(x[540]), .x541(x[541]), .x542(x[542]), .x543(x[543]), .x544(x[544]), .x545(x[545]), .x546(x[546]), .x547(x[547]), .x548(x[548]), .x549(x[549]), .x550(x[550]), .x551(x[551]), .x552(x[552]), .x553(x[553]), .x554(x[554]), .x555(x[555]), .x556(x[556]), .x557(x[557]), .x558(x[558]), .x559(x[559]), .x560(x[560]), .x561(x[561]), .x562(x[562]), .x563(x[563]), .x564(x[564]), .x565(x[565]), .x566(x[566]), .x567(x[567]), .x568(x[568]), .x569(x[569]), .x570(x[570]), .x571(x[571]), .x572(x[572]), .x573(x[573]), .x574(x[574]), .x575(x[575]), .x576(x[576]), .x577(x[577]), .x578(x[578]), .x579(x[579]), .x580(x[580]), .x581(x[581]), .x582(x[582]), .x583(x[583]), .x584(x[584]), .x585(x[585]), .x586(x[586]), .x587(x[587]), .x588(x[588]), .x589(x[589]), .x590(x[590]), .x591(x[591]), .x592(x[592]), .x593(x[593]), .x594(x[594]), .x595(x[595]), .x596(x[596]), .x597(x[597]), .x598(x[598]), .x599(x[599]), .x600(x[600]), .x601(x[601]), .x602(x[602]), .x603(x[603]), .x604(x[604]), .x605(x[605]), .x606(x[606]), .x607(x[607]), .x608(x[608]), .x609(x[609]), .x610(x[610]), .x611(x[611]), .x612(x[612]), .x613(x[613]), .x614(x[614]), .x615(x[615]), .x616(x[616]), .x617(x[617]), .x618(x[618]), .x619(x[619]), .x620(x[620]), .x621(x[621]), .x622(x[622]), .x623(x[623]), .x624(x[624]), .x625(x[625]), .x626(x[626]), .x627(x[627]), .x628(x[628]), .x629(x[629]), .x630(x[630]), .x631(x[631]), .x632(x[632]), .x633(x[633]), .x634(x[634]), .x635(x[635]), .x636(x[636]), .x637(x[637]), .x638(x[638]), .x639(x[639]), .x640(x[640]), .x641(x[641]), .x642(x[642]), .x643(x[643]), .x644(x[644]), .x645(x[645]), .x646(x[646]), .x647(x[647]), .x648(x[648]), .x649(x[649]), .x650(x[650]), .x651(x[651]), .x652(x[652]), .x653(x[653]), .x654(x[654]), .x655(x[655]), .x656(x[656]), .x657(x[657]), .x658(x[658]), .x659(x[659]), .x660(x[660]), .x661(x[661]), .x662(x[662]), .x663(x[663]), .x664(x[664]), .x665(x[665]), .x666(x[666]), .x667(x[667]), .x668(x[668]), .x669(x[669]), .x670(x[670]), .x671(x[671]), .x672(x[672]), .x673(x[673]), .x674(x[674]), .x675(x[675]), .x676(x[676]), .x677(x[677]), .x678(x[678]), .x679(x[679]), .x680(x[680]), .x681(x[681]), .x682(x[682]), .x683(x[683]), .x684(x[684]), .x685(x[685]), .x686(x[686]), .x687(x[687]), .x688(x[688]), .x689(x[689]), .x690(x[690]), .x691(x[691]), .x692(x[692]), .x693(x[693]), .x694(x[694]), .x695(x[695]), .x696(x[696]), .x697(x[697]), .x698(x[698]), .x699(x[699]), .x700(x[700]), .x701(x[701]), .x702(x[702]), .x703(x[703]), .x704(x[704]), .x705(x[705]), .x706(x[706]), .x707(x[707]), .x708(x[708]), .x709(x[709]), .x710(x[710]), .x711(x[711]), .x712(x[712]), .x713(x[713]), .x714(x[714]), .x715(x[715]), .x716(x[716]), .x717(x[717]), .x718(x[718]), .x719(x[719]), .x720(x[720]), .x721(x[721]), .x722(x[722]), .x723(x[723]), .x724(x[724]), .x725(x[725]), .x726(x[726]), .x727(x[727]), .x728(x[728]), .x729(x[729]), .x730(x[730]), .x731(x[731]), .x732(x[732]), .x733(x[733]), .x734(x[734]), .x735(x[735]), .x736(x[736]), .x737(x[737]), .x738(x[738]), .x739(x[739]), .x740(x[740]), .x741(x[741]), .x742(x[742]), .x743(x[743]), .x744(x[744]), .x745(x[745]), .x746(x[746]), .x747(x[747]), .x748(x[748]), .x749(x[749]), .x750(x[750]), .x751(x[751]), .x752(x[752]), .x753(x[753]), .x754(x[754]), .x755(x[755]), .x756(x[756]), .x757(x[757]), .x758(x[758]), .x759(x[759]), .x760(x[760]), .x761(x[761]), .x762(x[762]), .x763(x[763]), .x764(x[764]), .x765(x[765]), .x766(x[766]), .x767(x[767]), .x768(x[768]), .x769(x[769]), .x770(x[770]), .x771(x[771]), .x772(x[772]), .x773(x[773]), .x774(x[774]), .x775(x[775]), .x776(x[776]), .x777(x[777]), .x778(x[778]), .x779(x[779]), .x780(x[780]), .x781(x[781]), .x782(x[782]), .x783(x[783]), .x784(x[784]), .x785(x[785]), .x786(x[786]), .x787(x[787]), .x788(x[788]), .x789(x[789]), .x790(x[790]), .x791(x[791]), .x792(x[792]), .x793(x[793]), .x794(x[794]), .x795(x[795]), .x796(x[796]), .x797(x[797]), .x798(x[798]), .x799(x[799]), .x800(x[800]), .x801(x[801]), .x802(x[802]), .x803(x[803]), .x804(x[804]), .x805(x[805]), .x806(x[806]), .x807(x[807]), .x808(x[808]), .x809(x[809]), .x810(x[810]), .x811(x[811]), .x812(x[812]), .x813(x[813]), .x814(x[814]), .x815(x[815]), .x816(x[816]), .x817(x[817]), .x818(x[818]), .x819(x[819]), .x820(x[820]), .x821(x[821]), .x822(x[822]), .x823(x[823]), .x824(x[824]), .x825(x[825]), .x826(x[826]), .x827(x[827]), .x828(x[828]), .x829(x[829]), .x830(x[830]), .x831(x[831]), .x832(x[832]), .x833(x[833]), .x834(x[834]), .x835(x[835]), .x836(x[836]), .x837(x[837]), .x838(x[838]), .x839(x[839]), .x840(x[840]), .x841(x[841]), .x842(x[842]), .x843(x[843]), .x844(x[844]), .x845(x[845]), .x846(x[846]), .x847(x[847]), .x848(x[848]), .x849(x[849]), .x850(x[850]), .x851(x[851]), .x852(x[852]), .x853(x[853]), .x854(x[854]), .x855(x[855]), .x856(x[856]), .x857(x[857]), .x858(x[858]), .x859(x[859]), .x860(x[860]), .x861(x[861]), .x862(x[862]), .x863(x[863]), .x864(x[864]), .x865(x[865]), .x866(x[866]), .x867(x[867]), .x868(x[868]), .x869(x[869]), .x870(x[870]), .x871(x[871]), .x872(x[872]), .x873(x[873]), .x874(x[874]), .x875(x[875]), .x876(x[876]), .x877(x[877]), .x878(x[878]), .x879(x[879]), .x880(x[880]), .x881(x[881]), .x882(x[882]), .x883(x[883]), .x884(x[884]), .x885(x[885]), .x886(x[886]), .x887(x[887]), .x888(x[888]), .x889(x[889]), .x890(x[890]), .x891(x[891]), .x892(x[892]), .x893(x[893]), .x894(x[894]), .x895(x[895]), .x896(x[896]), .x897(x[897]), .x898(x[898]), .x899(x[899]), .x900(x[900]), .x901(x[901]), .x902(x[902]), .x903(x[903]), .x904(x[904]), .x905(x[905]), .x906(x[906]), .x907(x[907]), .x908(x[908]), .x909(x[909]), .x910(x[910]), .x911(x[911]), .x912(x[912]), .x913(x[913]), .x914(x[914]), .x915(x[915]), .x916(x[916]), .x917(x[917]), .x918(x[918]), .x919(x[919]), .x920(x[920]), .x921(x[921]), .x922(x[922]), .x923(x[923]), .x924(x[924]), .x925(x[925]), .x926(x[926]), .x927(x[927]), .x928(x[928]), .x929(x[929]), .x930(x[930]), .x931(x[931]), .x932(x[932]), .x933(x[933]), .x934(x[934]), .x935(x[935]), .x936(x[936]), .x937(x[937]), .x938(x[938]), .x939(x[939]), .x940(x[940]), .x941(x[941]), .x942(x[942]), .x943(x[943]), .x944(x[944]), .x945(x[945]), .x946(x[946]), .x947(x[947]), .x948(x[948]), .x949(x[949]), .x950(x[950]), .x951(x[951]), .x952(x[952]), .x953(x[953]), .x954(x[954]), .x955(x[955]), .x956(x[956]), .x957(x[957]), .x958(x[958]), .x959(x[959]), .x960(x[960]), .x961(x[961]), .x962(x[962]), .x963(x[963]), .x964(x[964]), .x965(x[965]), .x966(x[966]), .x967(x[967]), .x968(x[968]), .x969(x[969]), .x970(x[970]), .x971(x[971]), .x972(x[972]), .x973(x[973]), .x974(x[974]), .x975(x[975]), .x976(x[976]), .x977(x[977]), .x978(x[978]), .x979(x[979]), .x980(x[980]), .x981(x[981]), .x982(x[982]), .x983(x[983]), .x984(x[984]), .x985(x[985]), .x986(x[986]), .x987(x[987]), .x988(x[988]), .x989(x[989]), .x990(x[990]), .x991(x[991]), .x992(x[992]), .x993(x[993]), .x994(x[994]), .x995(x[995]), .x996(x[996]), .x997(x[997]), .x998(x[998]), .x999(x[999]), .x1000(x[1000]), .x1001(x[1001]), .x1002(x[1002]), .x1003(x[1003]), .x1004(x[1004]), .x1005(x[1005]), .x1006(x[1006]), .x1007(x[1007]), .x1008(x[1008]), .x1009(x[1009]), .x1010(x[1010]), .x1011(x[1011]), .x1012(x[1012]), .x1013(x[1013]), .x1014(x[1014]),
    .y0(y0)
  );

  // Optional reference function (majority reference for sanity check)
  function [9:0] popcount(input [1014:0] v);
    integer i; reg [9:0] c;
    begin
      c = 0;
      for (i = 0; i < 1015; i = i + 1)
        c = c + v[i];
      popcount = c;
    end
  endfunction

  // Reference majority: at least 508 ones
  wire y_ref = (popcount(x) >= 508);

  localparam [63:0] TOTAL_VECTORS = 64'd351111940402796075728379920075981393284761128699669252487168127261196632432619068618571244770327218791250222421623815151677323767215657465806342637967722899175327916845440400930277772658683777577056802640791026892262013051450122815378736544025053197584668966180832613749896964723593195907881555331297312768;

  initial begin
    $display("Time | x1014 x1013 x1012 x1011 x1010 x1009 x1008 x1007 x1006 x1005 x1004 x1003 x1002 x1001 x1000 x999 x998 x997 x996 x995 x994 x993 x992 x991 x990 x989 x988 x987 x986 x985 x984 x983 x982 x981 x980 x979 x978 x977 x976 x975 x974 x973 x972 x971 x970 x969 x968 x967 x966 x965 x964 x963 x962 x961 x960 x959 x958 x957 x956 x955 x954 x953 x952 x951 x950 x949 x948 x947 x946 x945 x944 x943 x942 x941 x940 x939 x938 x937 x936 x935 x934 x933 x932 x931 x930 x929 x928 x927 x926 x925 x924 x923 x922 x921 x920 x919 x918 x917 x916 x915 x914 x913 x912 x911 x910 x909 x908 x907 x906 x905 x904 x903 x902 x901 x900 x899 x898 x897 x896 x895 x894 x893 x892 x891 x890 x889 x888 x887 x886 x885 x884 x883 x882 x881 x880 x879 x878 x877 x876 x875 x874 x873 x872 x871 x870 x869 x868 x867 x866 x865 x864 x863 x862 x861 x860 x859 x858 x857 x856 x855 x854 x853 x852 x851 x850 x849 x848 x847 x846 x845 x844 x843 x842 x841 x840 x839 x838 x837 x836 x835 x834 x833 x832 x831 x830 x829 x828 x827 x826 x825 x824 x823 x822 x821 x820 x819 x818 x817 x816 x815 x814 x813 x812 x811 x810 x809 x808 x807 x806 x805 x804 x803 x802 x801 x800 x799 x798 x797 x796 x795 x794 x793 x792 x791 x790 x789 x788 x787 x786 x785 x784 x783 x782 x781 x780 x779 x778 x777 x776 x775 x774 x773 x772 x771 x770 x769 x768 x767 x766 x765 x764 x763 x762 x761 x760 x759 x758 x757 x756 x755 x754 x753 x752 x751 x750 x749 x748 x747 x746 x745 x744 x743 x742 x741 x740 x739 x738 x737 x736 x735 x734 x733 x732 x731 x730 x729 x728 x727 x726 x725 x724 x723 x722 x721 x720 x719 x718 x717 x716 x715 x714 x713 x712 x711 x710 x709 x708 x707 x706 x705 x704 x703 x702 x701 x700 x699 x698 x697 x696 x695 x694 x693 x692 x691 x690 x689 x688 x687 x686 x685 x684 x683 x682 x681 x680 x679 x678 x677 x676 x675 x674 x673 x672 x671 x670 x669 x668 x667 x666 x665 x664 x663 x662 x661 x660 x659 x658 x657 x656 x655 x654 x653 x652 x651 x650 x649 x648 x647 x646 x645 x644 x643 x642 x641 x640 x639 x638 x637 x636 x635 x634 x633 x632 x631 x630 x629 x628 x627 x626 x625 x624 x623 x622 x621 x620 x619 x618 x617 x616 x615 x614 x613 x612 x611 x610 x609 x608 x607 x606 x605 x604 x603 x602 x601 x600 x599 x598 x597 x596 x595 x594 x593 x592 x591 x590 x589 x588 x587 x586 x585 x584 x583 x582 x581 x580 x579 x578 x577 x576 x575 x574 x573 x572 x571 x570 x569 x568 x567 x566 x565 x564 x563 x562 x561 x560 x559 x558 x557 x556 x555 x554 x553 x552 x551 x550 x549 x548 x547 x546 x545 x544 x543 x542 x541 x540 x539 x538 x537 x536 x535 x534 x533 x532 x531 x530 x529 x528 x527 x526 x525 x524 x523 x522 x521 x520 x519 x518 x517 x516 x515 x514 x513 x512 x511 x510 x509 x508 x507 x506 x505 x504 x503 x502 x501 x500 x499 x498 x497 x496 x495 x494 x493 x492 x491 x490 x489 x488 x487 x486 x485 x484 x483 x482 x481 x480 x479 x478 x477 x476 x475 x474 x473 x472 x471 x470 x469 x468 x467 x466 x465 x464 x463 x462 x461 x460 x459 x458 x457 x456 x455 x454 x453 x452 x451 x450 x449 x448 x447 x446 x445 x444 x443 x442 x441 x440 x439 x438 x437 x436 x435 x434 x433 x432 x431 x430 x429 x428 x427 x426 x425 x424 x423 x422 x421 x420 x419 x418 x417 x416 x415 x414 x413 x412 x411 x410 x409 x408 x407 x406 x405 x404 x403 x402 x401 x400 x399 x398 x397 x396 x395 x394 x393 x392 x391 x390 x389 x388 x387 x386 x385 x384 x383 x382 x381 x380 x379 x378 x377 x376 x375 x374 x373 x372 x371 x370 x369 x368 x367 x366 x365 x364 x363 x362 x361 x360 x359 x358 x357 x356 x355 x354 x353 x352 x351 x350 x349 x348 x347 x346 x345 x344 x343 x342 x341 x340 x339 x338 x337 x336 x335 x334 x333 x332 x331 x330 x329 x328 x327 x326 x325 x324 x323 x322 x321 x320 x319 x318 x317 x316 x315 x314 x313 x312 x311 x310 x309 x308 x307 x306 x305 x304 x303 x302 x301 x300 x299 x298 x297 x296 x295 x294 x293 x292 x291 x290 x289 x288 x287 x286 x285 x284 x283 x282 x281 x280 x279 x278 x277 x276 x275 x274 x273 x272 x271 x270 x269 x268 x267 x266 x265 x264 x263 x262 x261 x260 x259 x258 x257 x256 x255 x254 x253 x252 x251 x250 x249 x248 x247 x246 x245 x244 x243 x242 x241 x240 x239 x238 x237 x236 x235 x234 x233 x232 x231 x230 x229 x228 x227 x226 x225 x224 x223 x222 x221 x220 x219 x218 x217 x216 x215 x214 x213 x212 x211 x210 x209 x208 x207 x206 x205 x204 x203 x202 x201 x200 x199 x198 x197 x196 x195 x194 x193 x192 x191 x190 x189 x188 x187 x186 x185 x184 x183 x182 x181 x180 x179 x178 x177 x176 x175 x174 x173 x172 x171 x170 x169 x168 x167 x166 x165 x164 x163 x162 x161 x160 x159 x158 x157 x156 x155 x154 x153 x152 x151 x150 x149 x148 x147 x146 x145 x144 x143 x142 x141 x140 x139 x138 x137 x136 x135 x134 x133 x132 x131 x130 x129 x128 x127 x126 x125 x124 x123 x122 x121 x120 x119 x118 x117 x116 x115 x114 x113 x112 x111 x110 x109 x108 x107 x106 x105 x104 x103 x102 x101 x100 x99 x98 x97 x96 x95 x94 x93 x92 x91 x90 x89 x88 x87 x86 x85 x84 x83 x82 x81 x80 x79 x78 x77 x76 x75 x74 x73 x72 x71 x70 x69 x68 x67 x66 x65 x64 x63 x62 x61 x60 x59 x58 x57 x56 x55 x54 x53 x52 x51 x50 x49 x48 x47 x46 x45 x44 x43 x42 x41 x40 x39 x38 x37 x36 x35 x34 x33 x32 x31 x30 x29 x28 x27 x26 x25 x24 x23 x22 x21 x20 x19 x18 x17 x16 x15 x14 x13 x12 x11 x10 x9 x8 x7 x6 x5 x4 x3 x2 x1 x0 | y0 (DUT) y_ref (Maj1015)");
    $display("---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------");
    // Loop through all 351111940402796075728379920075981393284761128699669252487168127261196632432619068618571244770327218791250222421623815151677323767215657465806342637967722899175327916845440400930277772658683777577056802640791026892262013051450122815378736544025053197584668966180832613749896964723593195907881555331297312768 combinations
    for (idx = 0; idx < TOTAL_VECTORS; idx = idx + 1) begin
      x = idx[1014:0];
      #10 $display("%4t |  %b  |   %b       %b",
                   $time, x, y0, y_ref);
    end
    #10 $finish;
  end

  // Optional mismatch check
  always #1 if (^x !== 1'bx && y0 !== y_ref)
    $display("Mismatch at t=%0t x=%b HW=%0d y0=%0b ref=%0b",
             $time, x, popcount(x), y0, y_ref);

endmodule

`default_nettype wire
