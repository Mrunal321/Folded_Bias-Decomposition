module top (x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255, x256, x257, x258, x259, x260, x261, x262, x263, x264, x265, x266, x267, x268, x269, x270, x271, x272, x273, x274, x275, x276, x277, x278, x279, x280, x281, x282, x283, x284, x285, x286, x287, x288, x289, x290, x291, x292, x293, x294, x295, x296, x297, x298, x299, x300, x301, x302, x303, x304, x305, x306, x307, x308, x309, x310, x311, x312, x313, x314, x315, x316, x317, x318, x319, x320, x321, x322, x323, x324, x325, x326, x327, x328, x329, x330, x331, x332, x333, x334, x335, x336, x337, x338, x339, x340, x341, x342, x343, x344, x345, x346, x347, x348, x349, x350, x351, x352, x353, x354, x355, x356, x357, x358, x359, x360, x361, x362, x363, x364, x365, x366, x367, x368, x369, x370, x371, x372, x373, x374, x375, x376, x377, x378, x379, x380, x381, x382, x383, x384, x385, x386, x387, x388, x389, x390, x391, x392, x393, x394, x395, x396, x397, x398, x399, x400, x401, x402, x403, x404, x405, x406, x407, x408, x409, x410, x411, x412, x413, x414, x415, x416, x417, x418, x419, x420, x421, x422, x423, x424, x425, x426, x427, x428, x429, x430, x431, x432, x433, x434, x435, x436, x437, x438, x439, x440, x441, x442, x443, x444, x445, x446, x447, x448, x449, x450, x451, x452, x453, x454, x455, x456, x457, x458, x459, x460, x461, x462, x463, x464, x465, x466, x467, x468, x469, x470, x471, x472, x473, x474, x475, x476, x477, x478, x479, x480, x481, x482, x483, x484, x485, x486, x487, x488, x489, x490, x491, x492, x493, x494, x495, x496, x497, x498, x499, x500, x501, x502, x503, x504, x505, x506, x507, x508, x509, x510, x511, x512, x513, x514, x515, x516, x517, x518, x519, x520, x521, x522, x523, x524, x525, x526, x527, x528, x529, x530, x531, x532, x533, x534, x535, x536, x537, x538, x539, x540, x541, x542, x543, x544, x545, x546, x547, x548, x549, x550, x551, x552, x553, x554, x555, x556, x557, x558, x559, x560, x561, x562, x563, x564, x565, x566, x567, x568, x569, x570, x571, x572, x573, x574, x575, x576, x577, x578, x579, x580, x581, x582, x583, x584, x585, x586, x587, x588, x589, x590, x591, x592, x593, x594, x595, x596, x597, x598, x599, x600, x601, x602, x603, x604, x605, x606, x607, x608, x609, x610, x611, x612, x613, x614, x615, x616, x617, x618, x619, x620, x621, x622, x623, x624, x625, x626, x627, x628, x629, x630, x631, x632, x633, x634, x635, x636, x637, x638, x639, x640, x641, x642, x643, x644, x645, x646, x647, x648, x649, x650, x651, x652, x653, x654, x655, x656, x657, x658, x659, x660, x661, x662, x663, x664, x665, x666, x667, x668, x669, x670, x671, x672, x673, x674, x675, x676, x677, x678, x679, x680, x681, x682, x683, x684, x685, x686, x687, x688, x689, x690, x691, x692, x693, x694, x695, x696, x697, x698, x699, x700, x701, x702, x703, x704, x705, x706, x707, x708, x709, x710, x711, x712, x713, x714, x715, x716, x717, x718, x719, x720, x721, x722, x723, x724, x725, x726, x727, x728, x729, x730, x731, x732, x733, x734, x735, x736, x737, x738, x739, x740, x741, x742, x743, x744, x745, x746, x747, x748, x749, x750, x751, x752, x753, x754, x755, x756, x757, x758, x759, x760, x761, x762, x763, x764, x765, x766, x767, x768, x769, x770, x771, x772, x773, x774, x775, x776, x777, x778, x779, x780, x781, x782, x783, x784, x785, x786, x787, x788, x789, x790, x791, x792, x793, x794, x795, x796, x797, x798, x799, x800, x801, x802, x803, x804, x805, x806, x807, x808, x809, x810, x811, x812, x813, x814, x815, x816, x817, x818, x819, x820, x821, x822, x823, x824, x825, x826, x827, x828, x829, x830, x831, x832, x833, x834, x835, x836, x837, x838, x839, x840, x841, x842, x843, x844, x845, x846, x847, x848, x849, x850, x851, x852, x853, x854, x855, x856, x857, x858, x859, x860, x861, x862, x863, x864, x865, x866, x867, x868, x869, x870, x871, x872, x873, x874, x875, x876, x877, x878, x879, x880, x881, x882, x883, x884, x885, x886, x887, x888, x889, x890, x891, x892, x893, x894, x895, x896, x897, x898, x899, x900, x901, x902, x903, x904, x905, x906, x907, x908, x909, x910, x911, x912, x913, x914, x915, x916, x917, x918, x919, x920, x921, x922, x923, x924, x925, x926, x927, x928, x929, x930, x931, x932, x933, x934, x935, x936, x937, x938, x939, x940, x941, x942, x943, x944, x945, x946, x947, x948, x949, x950, x951, x952, x953, x954, x955, x956, x957, x958, x959, x960, x961, x962, x963, x964, x965, x966, x967, x968, x969, x970, x971, x972, x973, x974, x975, x976, x977, x978, x979, x980, x981, x982, x983, x984, x985, x986, x987, x988, x989, x990, x991, x992, x993, x994, x995, x996, x997, x998, x999, x1000, x1001, x1002, x1003, x1004, x1005, x1006, x1007, x1008, x1009, x1010, x1011, x1012, x1013, x1014, y0);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, x39, x40, x41, x42, x43, x44, x45, x46, x47, x48, x49, x50, x51, x52, x53, x54, x55, x56, x57, x58, x59, x60, x61, x62, x63, x64, x65, x66, x67, x68, x69, x70, x71, x72, x73, x74, x75, x76, x77, x78, x79, x80, x81, x82, x83, x84, x85, x86, x87, x88, x89, x90, x91, x92, x93, x94, x95, x96, x97, x98, x99, x100, x101, x102, x103, x104, x105, x106, x107, x108, x109, x110, x111, x112, x113, x114, x115, x116, x117, x118, x119, x120, x121, x122, x123, x124, x125, x126, x127, x128, x129, x130, x131, x132, x133, x134, x135, x136, x137, x138, x139, x140, x141, x142, x143, x144, x145, x146, x147, x148, x149, x150, x151, x152, x153, x154, x155, x156, x157, x158, x159, x160, x161, x162, x163, x164, x165, x166, x167, x168, x169, x170, x171, x172, x173, x174, x175, x176, x177, x178, x179, x180, x181, x182, x183, x184, x185, x186, x187, x188, x189, x190, x191, x192, x193, x194, x195, x196, x197, x198, x199, x200, x201, x202, x203, x204, x205, x206, x207, x208, x209, x210, x211, x212, x213, x214, x215, x216, x217, x218, x219, x220, x221, x222, x223, x224, x225, x226, x227, x228, x229, x230, x231, x232, x233, x234, x235, x236, x237, x238, x239, x240, x241, x242, x243, x244, x245, x246, x247, x248, x249, x250, x251, x252, x253, x254, x255, x256, x257, x258, x259, x260, x261, x262, x263, x264, x265, x266, x267, x268, x269, x270, x271, x272, x273, x274, x275, x276, x277, x278, x279, x280, x281, x282, x283, x284, x285, x286, x287, x288, x289, x290, x291, x292, x293, x294, x295, x296, x297, x298, x299, x300, x301, x302, x303, x304, x305, x306, x307, x308, x309, x310, x311, x312, x313, x314, x315, x316, x317, x318, x319, x320, x321, x322, x323, x324, x325, x326, x327, x328, x329, x330, x331, x332, x333, x334, x335, x336, x337, x338, x339, x340, x341, x342, x343, x344, x345, x346, x347, x348, x349, x350, x351, x352, x353, x354, x355, x356, x357, x358, x359, x360, x361, x362, x363, x364, x365, x366, x367, x368, x369, x370, x371, x372, x373, x374, x375, x376, x377, x378, x379, x380, x381, x382, x383, x384, x385, x386, x387, x388, x389, x390, x391, x392, x393, x394, x395, x396, x397, x398, x399, x400, x401, x402, x403, x404, x405, x406, x407, x408, x409, x410, x411, x412, x413, x414, x415, x416, x417, x418, x419, x420, x421, x422, x423, x424, x425, x426, x427, x428, x429, x430, x431, x432, x433, x434, x435, x436, x437, x438, x439, x440, x441, x442, x443, x444, x445, x446, x447, x448, x449, x450, x451, x452, x453, x454, x455, x456, x457, x458, x459, x460, x461, x462, x463, x464, x465, x466, x467, x468, x469, x470, x471, x472, x473, x474, x475, x476, x477, x478, x479, x480, x481, x482, x483, x484, x485, x486, x487, x488, x489, x490, x491, x492, x493, x494, x495, x496, x497, x498, x499, x500, x501, x502, x503, x504, x505, x506, x507, x508, x509, x510, x511, x512, x513, x514, x515, x516, x517, x518, x519, x520, x521, x522, x523, x524, x525, x526, x527, x528, x529, x530, x531, x532, x533, x534, x535, x536, x537, x538, x539, x540, x541, x542, x543, x544, x545, x546, x547, x548, x549, x550, x551, x552, x553, x554, x555, x556, x557, x558, x559, x560, x561, x562, x563, x564, x565, x566, x567, x568, x569, x570, x571, x572, x573, x574, x575, x576, x577, x578, x579, x580, x581, x582, x583, x584, x585, x586, x587, x588, x589, x590, x591, x592, x593, x594, x595, x596, x597, x598, x599, x600, x601, x602, x603, x604, x605, x606, x607, x608, x609, x610, x611, x612, x613, x614, x615, x616, x617, x618, x619, x620, x621, x622, x623, x624, x625, x626, x627, x628, x629, x630, x631, x632, x633, x634, x635, x636, x637, x638, x639, x640, x641, x642, x643, x644, x645, x646, x647, x648, x649, x650, x651, x652, x653, x654, x655, x656, x657, x658, x659, x660, x661, x662, x663, x664, x665, x666, x667, x668, x669, x670, x671, x672, x673, x674, x675, x676, x677, x678, x679, x680, x681, x682, x683, x684, x685, x686, x687, x688, x689, x690, x691, x692, x693, x694, x695, x696, x697, x698, x699, x700, x701, x702, x703, x704, x705, x706, x707, x708, x709, x710, x711, x712, x713, x714, x715, x716, x717, x718, x719, x720, x721, x722, x723, x724, x725, x726, x727, x728, x729, x730, x731, x732, x733, x734, x735, x736, x737, x738, x739, x740, x741, x742, x743, x744, x745, x746, x747, x748, x749, x750, x751, x752, x753, x754, x755, x756, x757, x758, x759, x760, x761, x762, x763, x764, x765, x766, x767, x768, x769, x770, x771, x772, x773, x774, x775, x776, x777, x778, x779, x780, x781, x782, x783, x784, x785, x786, x787, x788, x789, x790, x791, x792, x793, x794, x795, x796, x797, x798, x799, x800, x801, x802, x803, x804, x805, x806, x807, x808, x809, x810, x811, x812, x813, x814, x815, x816, x817, x818, x819, x820, x821, x822, x823, x824, x825, x826, x827, x828, x829, x830, x831, x832, x833, x834, x835, x836, x837, x838, x839, x840, x841, x842, x843, x844, x845, x846, x847, x848, x849, x850, x851, x852, x853, x854, x855, x856, x857, x858, x859, x860, x861, x862, x863, x864, x865, x866, x867, x868, x869, x870, x871, x872, x873, x874, x875, x876, x877, x878, x879, x880, x881, x882, x883, x884, x885, x886, x887, x888, x889, x890, x891, x892, x893, x894, x895, x896, x897, x898, x899, x900, x901, x902, x903, x904, x905, x906, x907, x908, x909, x910, x911, x912, x913, x914, x915, x916, x917, x918, x919, x920, x921, x922, x923, x924, x925, x926, x927, x928, x929, x930, x931, x932, x933, x934, x935, x936, x937, x938, x939, x940, x941, x942, x943, x944, x945, x946, x947, x948, x949, x950, x951, x952, x953, x954, x955, x956, x957, x958, x959, x960, x961, x962, x963, x964, x965, x966, x967, x968, x969, x970, x971, x972, x973, x974, x975, x976, x977, x978, x979, x980, x981, x982, x983, x984, x985, x986, x987, x988, x989, x990, x991, x992, x993, x994, x995, x996, x997, x998, x999, x1000, x1001, x1002, x1003, x1004, x1005, x1006, x1007, x1008, x1009, x1010, x1011, x1012, x1013, x1014;
  output y0;
  wire n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674;
  LUT3 #(.INIT(8'hE8)) lut_n1017 (.I0(x0), .I1(x1), .I2(x2), .O(n1017));
  LUT3 #(.INIT(8'hE8)) lut_n1018 (.I0(x6), .I1(x7), .I2(x8), .O(n1018));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1019 (.I0(x3), .I1(x4), .I2(x5), .I3(n1017), .I4(n1018), .O(n1019));
  LUT3 #(.INIT(8'hE8)) lut_n1020 (.I0(x12), .I1(x13), .I2(x14), .O(n1020));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1021 (.I0(x3), .I1(x4), .I2(x5), .I3(n1017), .I4(n1018), .O(n1021));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1022 (.I0(x9), .I1(x10), .I2(x11), .I3(n1020), .I4(n1021), .O(n1022));
  LUT3 #(.INIT(8'hE8)) lut_n1023 (.I0(x18), .I1(x19), .I2(x20), .O(n1023));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1024 (.I0(x9), .I1(x10), .I2(x11), .I3(n1020), .I4(n1021), .O(n1024));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1025 (.I0(x15), .I1(x16), .I2(x17), .I3(n1023), .I4(n1024), .O(n1025));
  LUT3 #(.INIT(8'hE8)) lut_n1026 (.I0(n1019), .I1(n1022), .I2(n1025), .O(n1026));
  LUT3 #(.INIT(8'hE8)) lut_n1027 (.I0(x24), .I1(x25), .I2(x26), .O(n1027));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1028 (.I0(x15), .I1(x16), .I2(x17), .I3(n1023), .I4(n1024), .O(n1028));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1029 (.I0(x21), .I1(x22), .I2(x23), .I3(n1027), .I4(n1028), .O(n1029));
  LUT3 #(.INIT(8'hE8)) lut_n1030 (.I0(x27), .I1(x28), .I2(x29), .O(n1030));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1031 (.I0(x21), .I1(x22), .I2(x23), .I3(n1027), .I4(n1028), .O(n1031));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1032 (.I0(x30), .I1(x31), .I2(x32), .I3(n1030), .I4(n1031), .O(n1032));
  LUT3 #(.INIT(8'h96)) lut_n1033 (.I0(n1019), .I1(n1022), .I2(n1025), .O(n1033));
  LUT3 #(.INIT(8'hE8)) lut_n1034 (.I0(n1029), .I1(n1032), .I2(n1033), .O(n1034));
  LUT3 #(.INIT(8'hE8)) lut_n1035 (.I0(x36), .I1(x37), .I2(x38), .O(n1035));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1036 (.I0(x30), .I1(x31), .I2(x32), .I3(n1030), .I4(n1031), .O(n1036));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1037 (.I0(x33), .I1(x34), .I2(x35), .I3(n1035), .I4(n1036), .O(n1037));
  LUT3 #(.INIT(8'hE8)) lut_n1038 (.I0(x42), .I1(x43), .I2(x44), .O(n1038));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1039 (.I0(x33), .I1(x34), .I2(x35), .I3(n1035), .I4(n1036), .O(n1039));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1040 (.I0(x39), .I1(x40), .I2(x41), .I3(n1038), .I4(n1039), .O(n1040));
  LUT3 #(.INIT(8'h96)) lut_n1041 (.I0(n1029), .I1(n1032), .I2(n1033), .O(n1041));
  LUT3 #(.INIT(8'hE8)) lut_n1042 (.I0(n1037), .I1(n1040), .I2(n1041), .O(n1042));
  LUT3 #(.INIT(8'hE8)) lut_n1043 (.I0(n1026), .I1(n1034), .I2(n1042), .O(n1043));
  LUT3 #(.INIT(8'hE8)) lut_n1044 (.I0(x48), .I1(x49), .I2(x50), .O(n1044));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1045 (.I0(x39), .I1(x40), .I2(x41), .I3(n1038), .I4(n1039), .O(n1045));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1046 (.I0(x45), .I1(x46), .I2(x47), .I3(n1044), .I4(n1045), .O(n1046));
  LUT3 #(.INIT(8'hE8)) lut_n1047 (.I0(x54), .I1(x55), .I2(x56), .O(n1047));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1048 (.I0(x45), .I1(x46), .I2(x47), .I3(n1044), .I4(n1045), .O(n1048));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1049 (.I0(x51), .I1(x52), .I2(x53), .I3(n1047), .I4(n1048), .O(n1049));
  LUT3 #(.INIT(8'h96)) lut_n1050 (.I0(n1037), .I1(n1040), .I2(n1041), .O(n1050));
  LUT3 #(.INIT(8'hE8)) lut_n1051 (.I0(n1046), .I1(n1049), .I2(n1050), .O(n1051));
  LUT3 #(.INIT(8'hE8)) lut_n1052 (.I0(x60), .I1(x61), .I2(x62), .O(n1052));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1053 (.I0(x51), .I1(x52), .I2(x53), .I3(n1047), .I4(n1048), .O(n1053));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1054 (.I0(x57), .I1(x58), .I2(x59), .I3(n1052), .I4(n1053), .O(n1054));
  LUT3 #(.INIT(8'hE8)) lut_n1055 (.I0(x66), .I1(x67), .I2(x68), .O(n1055));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1056 (.I0(x57), .I1(x58), .I2(x59), .I3(n1052), .I4(n1053), .O(n1056));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1057 (.I0(x63), .I1(x64), .I2(x65), .I3(n1055), .I4(n1056), .O(n1057));
  LUT3 #(.INIT(8'h96)) lut_n1058 (.I0(n1046), .I1(n1049), .I2(n1050), .O(n1058));
  LUT3 #(.INIT(8'hE8)) lut_n1059 (.I0(n1054), .I1(n1057), .I2(n1058), .O(n1059));
  LUT3 #(.INIT(8'h96)) lut_n1060 (.I0(n1026), .I1(n1034), .I2(n1042), .O(n1060));
  LUT3 #(.INIT(8'hE8)) lut_n1061 (.I0(n1051), .I1(n1059), .I2(n1060), .O(n1061));
  LUT3 #(.INIT(8'hE8)) lut_n1062 (.I0(x72), .I1(x73), .I2(x74), .O(n1062));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1063 (.I0(x63), .I1(x64), .I2(x65), .I3(n1055), .I4(n1056), .O(n1063));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1064 (.I0(x69), .I1(x70), .I2(x71), .I3(n1062), .I4(n1063), .O(n1064));
  LUT3 #(.INIT(8'hE8)) lut_n1065 (.I0(x78), .I1(x79), .I2(x80), .O(n1065));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1066 (.I0(x69), .I1(x70), .I2(x71), .I3(n1062), .I4(n1063), .O(n1066));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1067 (.I0(x75), .I1(x76), .I2(x77), .I3(n1065), .I4(n1066), .O(n1067));
  LUT3 #(.INIT(8'h96)) lut_n1068 (.I0(n1054), .I1(n1057), .I2(n1058), .O(n1068));
  LUT3 #(.INIT(8'hE8)) lut_n1069 (.I0(n1064), .I1(n1067), .I2(n1068), .O(n1069));
  LUT3 #(.INIT(8'hE8)) lut_n1070 (.I0(x84), .I1(x85), .I2(x86), .O(n1070));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1071 (.I0(x75), .I1(x76), .I2(x77), .I3(n1065), .I4(n1066), .O(n1071));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1072 (.I0(x81), .I1(x82), .I2(x83), .I3(n1070), .I4(n1071), .O(n1072));
  LUT3 #(.INIT(8'hE8)) lut_n1073 (.I0(x90), .I1(x91), .I2(x92), .O(n1073));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1074 (.I0(x81), .I1(x82), .I2(x83), .I3(n1070), .I4(n1071), .O(n1074));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1075 (.I0(x87), .I1(x88), .I2(x89), .I3(n1073), .I4(n1074), .O(n1075));
  LUT3 #(.INIT(8'h96)) lut_n1076 (.I0(n1064), .I1(n1067), .I2(n1068), .O(n1076));
  LUT3 #(.INIT(8'hE8)) lut_n1077 (.I0(n1072), .I1(n1075), .I2(n1076), .O(n1077));
  LUT3 #(.INIT(8'h96)) lut_n1078 (.I0(n1051), .I1(n1059), .I2(n1060), .O(n1078));
  LUT3 #(.INIT(8'hE8)) lut_n1079 (.I0(n1069), .I1(n1077), .I2(n1078), .O(n1079));
  LUT3 #(.INIT(8'hE8)) lut_n1080 (.I0(n1043), .I1(n1061), .I2(n1079), .O(n1080));
  LUT3 #(.INIT(8'hE8)) lut_n1081 (.I0(x96), .I1(x97), .I2(x98), .O(n1081));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1082 (.I0(x87), .I1(x88), .I2(x89), .I3(n1073), .I4(n1074), .O(n1082));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1083 (.I0(x93), .I1(x94), .I2(x95), .I3(n1081), .I4(n1082), .O(n1083));
  LUT3 #(.INIT(8'hE8)) lut_n1084 (.I0(x102), .I1(x103), .I2(x104), .O(n1084));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1085 (.I0(x93), .I1(x94), .I2(x95), .I3(n1081), .I4(n1082), .O(n1085));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1086 (.I0(x99), .I1(x100), .I2(x101), .I3(n1084), .I4(n1085), .O(n1086));
  LUT3 #(.INIT(8'h96)) lut_n1087 (.I0(n1072), .I1(n1075), .I2(n1076), .O(n1087));
  LUT3 #(.INIT(8'hE8)) lut_n1088 (.I0(n1083), .I1(n1086), .I2(n1087), .O(n1088));
  LUT3 #(.INIT(8'hE8)) lut_n1089 (.I0(x108), .I1(x109), .I2(x110), .O(n1089));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1090 (.I0(x99), .I1(x100), .I2(x101), .I3(n1084), .I4(n1085), .O(n1090));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1091 (.I0(x105), .I1(x106), .I2(x107), .I3(n1089), .I4(n1090), .O(n1091));
  LUT3 #(.INIT(8'hE8)) lut_n1092 (.I0(x114), .I1(x115), .I2(x116), .O(n1092));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1093 (.I0(x105), .I1(x106), .I2(x107), .I3(n1089), .I4(n1090), .O(n1093));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1094 (.I0(x111), .I1(x112), .I2(x113), .I3(n1092), .I4(n1093), .O(n1094));
  LUT3 #(.INIT(8'h96)) lut_n1095 (.I0(n1083), .I1(n1086), .I2(n1087), .O(n1095));
  LUT3 #(.INIT(8'hE8)) lut_n1096 (.I0(n1091), .I1(n1094), .I2(n1095), .O(n1096));
  LUT3 #(.INIT(8'h96)) lut_n1097 (.I0(n1069), .I1(n1077), .I2(n1078), .O(n1097));
  LUT3 #(.INIT(8'hE8)) lut_n1098 (.I0(n1088), .I1(n1096), .I2(n1097), .O(n1098));
  LUT3 #(.INIT(8'hE8)) lut_n1099 (.I0(x120), .I1(x121), .I2(x122), .O(n1099));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1100 (.I0(x111), .I1(x112), .I2(x113), .I3(n1092), .I4(n1093), .O(n1100));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1101 (.I0(x117), .I1(x118), .I2(x119), .I3(n1099), .I4(n1100), .O(n1101));
  LUT3 #(.INIT(8'hE8)) lut_n1102 (.I0(x126), .I1(x127), .I2(x128), .O(n1102));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1103 (.I0(x117), .I1(x118), .I2(x119), .I3(n1099), .I4(n1100), .O(n1103));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1104 (.I0(x123), .I1(x124), .I2(x125), .I3(n1102), .I4(n1103), .O(n1104));
  LUT3 #(.INIT(8'h96)) lut_n1105 (.I0(n1091), .I1(n1094), .I2(n1095), .O(n1105));
  LUT3 #(.INIT(8'hE8)) lut_n1106 (.I0(n1101), .I1(n1104), .I2(n1105), .O(n1106));
  LUT3 #(.INIT(8'hE8)) lut_n1107 (.I0(x132), .I1(x133), .I2(x134), .O(n1107));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1108 (.I0(x123), .I1(x124), .I2(x125), .I3(n1102), .I4(n1103), .O(n1108));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1109 (.I0(x129), .I1(x130), .I2(x131), .I3(n1107), .I4(n1108), .O(n1109));
  LUT3 #(.INIT(8'hE8)) lut_n1110 (.I0(x138), .I1(x139), .I2(x140), .O(n1110));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1111 (.I0(x129), .I1(x130), .I2(x131), .I3(n1107), .I4(n1108), .O(n1111));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1112 (.I0(x135), .I1(x136), .I2(x137), .I3(n1110), .I4(n1111), .O(n1112));
  LUT3 #(.INIT(8'h96)) lut_n1113 (.I0(n1101), .I1(n1104), .I2(n1105), .O(n1113));
  LUT3 #(.INIT(8'hE8)) lut_n1114 (.I0(n1109), .I1(n1112), .I2(n1113), .O(n1114));
  LUT3 #(.INIT(8'h96)) lut_n1115 (.I0(n1088), .I1(n1096), .I2(n1097), .O(n1115));
  LUT3 #(.INIT(8'hE8)) lut_n1116 (.I0(n1106), .I1(n1114), .I2(n1115), .O(n1116));
  LUT3 #(.INIT(8'h96)) lut_n1117 (.I0(n1043), .I1(n1061), .I2(n1079), .O(n1117));
  LUT3 #(.INIT(8'hE8)) lut_n1118 (.I0(n1098), .I1(n1116), .I2(n1117), .O(n1118));
  LUT3 #(.INIT(8'hE8)) lut_n1119 (.I0(x144), .I1(x145), .I2(x146), .O(n1119));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1120 (.I0(x135), .I1(x136), .I2(x137), .I3(n1110), .I4(n1111), .O(n1120));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1121 (.I0(x141), .I1(x142), .I2(x143), .I3(n1119), .I4(n1120), .O(n1121));
  LUT3 #(.INIT(8'hE8)) lut_n1122 (.I0(x150), .I1(x151), .I2(x152), .O(n1122));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1123 (.I0(x141), .I1(x142), .I2(x143), .I3(n1119), .I4(n1120), .O(n1123));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1124 (.I0(x147), .I1(x148), .I2(x149), .I3(n1122), .I4(n1123), .O(n1124));
  LUT3 #(.INIT(8'h96)) lut_n1125 (.I0(n1109), .I1(n1112), .I2(n1113), .O(n1125));
  LUT3 #(.INIT(8'hE8)) lut_n1126 (.I0(n1121), .I1(n1124), .I2(n1125), .O(n1126));
  LUT3 #(.INIT(8'hE8)) lut_n1127 (.I0(x156), .I1(x157), .I2(x158), .O(n1127));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1128 (.I0(x147), .I1(x148), .I2(x149), .I3(n1122), .I4(n1123), .O(n1128));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1129 (.I0(x153), .I1(x154), .I2(x155), .I3(n1127), .I4(n1128), .O(n1129));
  LUT3 #(.INIT(8'hE8)) lut_n1130 (.I0(x162), .I1(x163), .I2(x164), .O(n1130));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1131 (.I0(x153), .I1(x154), .I2(x155), .I3(n1127), .I4(n1128), .O(n1131));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1132 (.I0(x159), .I1(x160), .I2(x161), .I3(n1130), .I4(n1131), .O(n1132));
  LUT3 #(.INIT(8'h96)) lut_n1133 (.I0(n1121), .I1(n1124), .I2(n1125), .O(n1133));
  LUT3 #(.INIT(8'hE8)) lut_n1134 (.I0(n1129), .I1(n1132), .I2(n1133), .O(n1134));
  LUT3 #(.INIT(8'h96)) lut_n1135 (.I0(n1106), .I1(n1114), .I2(n1115), .O(n1135));
  LUT3 #(.INIT(8'hE8)) lut_n1136 (.I0(n1126), .I1(n1134), .I2(n1135), .O(n1136));
  LUT3 #(.INIT(8'hE8)) lut_n1137 (.I0(x168), .I1(x169), .I2(x170), .O(n1137));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1138 (.I0(x159), .I1(x160), .I2(x161), .I3(n1130), .I4(n1131), .O(n1138));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1139 (.I0(x165), .I1(x166), .I2(x167), .I3(n1137), .I4(n1138), .O(n1139));
  LUT3 #(.INIT(8'hE8)) lut_n1140 (.I0(x174), .I1(x175), .I2(x176), .O(n1140));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1141 (.I0(x165), .I1(x166), .I2(x167), .I3(n1137), .I4(n1138), .O(n1141));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1142 (.I0(x171), .I1(x172), .I2(x173), .I3(n1140), .I4(n1141), .O(n1142));
  LUT3 #(.INIT(8'h96)) lut_n1143 (.I0(n1129), .I1(n1132), .I2(n1133), .O(n1143));
  LUT3 #(.INIT(8'hE8)) lut_n1144 (.I0(n1139), .I1(n1142), .I2(n1143), .O(n1144));
  LUT3 #(.INIT(8'hE8)) lut_n1145 (.I0(x180), .I1(x181), .I2(x182), .O(n1145));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1146 (.I0(x171), .I1(x172), .I2(x173), .I3(n1140), .I4(n1141), .O(n1146));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1147 (.I0(x177), .I1(x178), .I2(x179), .I3(n1145), .I4(n1146), .O(n1147));
  LUT3 #(.INIT(8'hE8)) lut_n1148 (.I0(x186), .I1(x187), .I2(x188), .O(n1148));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1149 (.I0(x177), .I1(x178), .I2(x179), .I3(n1145), .I4(n1146), .O(n1149));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1150 (.I0(x183), .I1(x184), .I2(x185), .I3(n1148), .I4(n1149), .O(n1150));
  LUT3 #(.INIT(8'h96)) lut_n1151 (.I0(n1139), .I1(n1142), .I2(n1143), .O(n1151));
  LUT3 #(.INIT(8'hE8)) lut_n1152 (.I0(n1147), .I1(n1150), .I2(n1151), .O(n1152));
  LUT3 #(.INIT(8'h96)) lut_n1153 (.I0(n1126), .I1(n1134), .I2(n1135), .O(n1153));
  LUT3 #(.INIT(8'hE8)) lut_n1154 (.I0(n1144), .I1(n1152), .I2(n1153), .O(n1154));
  LUT3 #(.INIT(8'h96)) lut_n1155 (.I0(n1098), .I1(n1116), .I2(n1117), .O(n1155));
  LUT3 #(.INIT(8'hE8)) lut_n1156 (.I0(n1136), .I1(n1154), .I2(n1155), .O(n1156));
  LUT3 #(.INIT(8'hE8)) lut_n1157 (.I0(n1080), .I1(n1118), .I2(n1156), .O(n1157));
  LUT3 #(.INIT(8'hE8)) lut_n1158 (.I0(x192), .I1(x193), .I2(x194), .O(n1158));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1159 (.I0(x183), .I1(x184), .I2(x185), .I3(n1148), .I4(n1149), .O(n1159));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1160 (.I0(x189), .I1(x190), .I2(x191), .I3(n1158), .I4(n1159), .O(n1160));
  LUT3 #(.INIT(8'hE8)) lut_n1161 (.I0(x198), .I1(x199), .I2(x200), .O(n1161));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1162 (.I0(x189), .I1(x190), .I2(x191), .I3(n1158), .I4(n1159), .O(n1162));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1163 (.I0(x195), .I1(x196), .I2(x197), .I3(n1161), .I4(n1162), .O(n1163));
  LUT3 #(.INIT(8'h96)) lut_n1164 (.I0(n1147), .I1(n1150), .I2(n1151), .O(n1164));
  LUT3 #(.INIT(8'hE8)) lut_n1165 (.I0(n1160), .I1(n1163), .I2(n1164), .O(n1165));
  LUT3 #(.INIT(8'hE8)) lut_n1166 (.I0(x204), .I1(x205), .I2(x206), .O(n1166));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1167 (.I0(x195), .I1(x196), .I2(x197), .I3(n1161), .I4(n1162), .O(n1167));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1168 (.I0(x201), .I1(x202), .I2(x203), .I3(n1166), .I4(n1167), .O(n1168));
  LUT3 #(.INIT(8'hE8)) lut_n1169 (.I0(x210), .I1(x211), .I2(x212), .O(n1169));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1170 (.I0(x201), .I1(x202), .I2(x203), .I3(n1166), .I4(n1167), .O(n1170));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1171 (.I0(x207), .I1(x208), .I2(x209), .I3(n1169), .I4(n1170), .O(n1171));
  LUT3 #(.INIT(8'h96)) lut_n1172 (.I0(n1160), .I1(n1163), .I2(n1164), .O(n1172));
  LUT3 #(.INIT(8'hE8)) lut_n1173 (.I0(n1168), .I1(n1171), .I2(n1172), .O(n1173));
  LUT3 #(.INIT(8'h96)) lut_n1174 (.I0(n1144), .I1(n1152), .I2(n1153), .O(n1174));
  LUT3 #(.INIT(8'hE8)) lut_n1175 (.I0(n1165), .I1(n1173), .I2(n1174), .O(n1175));
  LUT3 #(.INIT(8'hE8)) lut_n1176 (.I0(x216), .I1(x217), .I2(x218), .O(n1176));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1177 (.I0(x207), .I1(x208), .I2(x209), .I3(n1169), .I4(n1170), .O(n1177));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1178 (.I0(x213), .I1(x214), .I2(x215), .I3(n1176), .I4(n1177), .O(n1178));
  LUT3 #(.INIT(8'hE8)) lut_n1179 (.I0(x222), .I1(x223), .I2(x224), .O(n1179));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1180 (.I0(x213), .I1(x214), .I2(x215), .I3(n1176), .I4(n1177), .O(n1180));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1181 (.I0(x219), .I1(x220), .I2(x221), .I3(n1179), .I4(n1180), .O(n1181));
  LUT3 #(.INIT(8'h96)) lut_n1182 (.I0(n1168), .I1(n1171), .I2(n1172), .O(n1182));
  LUT3 #(.INIT(8'hE8)) lut_n1183 (.I0(n1178), .I1(n1181), .I2(n1182), .O(n1183));
  LUT3 #(.INIT(8'hE8)) lut_n1184 (.I0(x228), .I1(x229), .I2(x230), .O(n1184));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1185 (.I0(x219), .I1(x220), .I2(x221), .I3(n1179), .I4(n1180), .O(n1185));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1186 (.I0(x225), .I1(x226), .I2(x227), .I3(n1184), .I4(n1185), .O(n1186));
  LUT3 #(.INIT(8'hE8)) lut_n1187 (.I0(x234), .I1(x235), .I2(x236), .O(n1187));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1188 (.I0(x225), .I1(x226), .I2(x227), .I3(n1184), .I4(n1185), .O(n1188));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1189 (.I0(x231), .I1(x232), .I2(x233), .I3(n1187), .I4(n1188), .O(n1189));
  LUT3 #(.INIT(8'h96)) lut_n1190 (.I0(n1178), .I1(n1181), .I2(n1182), .O(n1190));
  LUT3 #(.INIT(8'hE8)) lut_n1191 (.I0(n1186), .I1(n1189), .I2(n1190), .O(n1191));
  LUT3 #(.INIT(8'h96)) lut_n1192 (.I0(n1165), .I1(n1173), .I2(n1174), .O(n1192));
  LUT3 #(.INIT(8'hE8)) lut_n1193 (.I0(n1183), .I1(n1191), .I2(n1192), .O(n1193));
  LUT3 #(.INIT(8'h96)) lut_n1194 (.I0(n1136), .I1(n1154), .I2(n1155), .O(n1194));
  LUT3 #(.INIT(8'hE8)) lut_n1195 (.I0(n1175), .I1(n1193), .I2(n1194), .O(n1195));
  LUT3 #(.INIT(8'hE8)) lut_n1196 (.I0(x240), .I1(x241), .I2(x242), .O(n1196));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1197 (.I0(x231), .I1(x232), .I2(x233), .I3(n1187), .I4(n1188), .O(n1197));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1198 (.I0(x237), .I1(x238), .I2(x239), .I3(n1196), .I4(n1197), .O(n1198));
  LUT3 #(.INIT(8'hE8)) lut_n1199 (.I0(x246), .I1(x247), .I2(x248), .O(n1199));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1200 (.I0(x237), .I1(x238), .I2(x239), .I3(n1196), .I4(n1197), .O(n1200));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1201 (.I0(x243), .I1(x244), .I2(x245), .I3(n1199), .I4(n1200), .O(n1201));
  LUT3 #(.INIT(8'h96)) lut_n1202 (.I0(n1186), .I1(n1189), .I2(n1190), .O(n1202));
  LUT3 #(.INIT(8'hE8)) lut_n1203 (.I0(n1198), .I1(n1201), .I2(n1202), .O(n1203));
  LUT3 #(.INIT(8'hE8)) lut_n1204 (.I0(x252), .I1(x253), .I2(x254), .O(n1204));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1205 (.I0(x243), .I1(x244), .I2(x245), .I3(n1199), .I4(n1200), .O(n1205));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1206 (.I0(x249), .I1(x250), .I2(x251), .I3(n1204), .I4(n1205), .O(n1206));
  LUT3 #(.INIT(8'hE8)) lut_n1207 (.I0(x258), .I1(x259), .I2(x260), .O(n1207));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1208 (.I0(x249), .I1(x250), .I2(x251), .I3(n1204), .I4(n1205), .O(n1208));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1209 (.I0(x255), .I1(x256), .I2(x257), .I3(n1207), .I4(n1208), .O(n1209));
  LUT3 #(.INIT(8'h96)) lut_n1210 (.I0(n1198), .I1(n1201), .I2(n1202), .O(n1210));
  LUT3 #(.INIT(8'hE8)) lut_n1211 (.I0(n1206), .I1(n1209), .I2(n1210), .O(n1211));
  LUT3 #(.INIT(8'h96)) lut_n1212 (.I0(n1183), .I1(n1191), .I2(n1192), .O(n1212));
  LUT3 #(.INIT(8'hE8)) lut_n1213 (.I0(n1203), .I1(n1211), .I2(n1212), .O(n1213));
  LUT3 #(.INIT(8'hE8)) lut_n1214 (.I0(x264), .I1(x265), .I2(x266), .O(n1214));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1215 (.I0(x255), .I1(x256), .I2(x257), .I3(n1207), .I4(n1208), .O(n1215));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1216 (.I0(x261), .I1(x262), .I2(x263), .I3(n1214), .I4(n1215), .O(n1216));
  LUT3 #(.INIT(8'hE8)) lut_n1217 (.I0(x270), .I1(x271), .I2(x272), .O(n1217));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1218 (.I0(x261), .I1(x262), .I2(x263), .I3(n1214), .I4(n1215), .O(n1218));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1219 (.I0(x267), .I1(x268), .I2(x269), .I3(n1217), .I4(n1218), .O(n1219));
  LUT3 #(.INIT(8'h96)) lut_n1220 (.I0(n1206), .I1(n1209), .I2(n1210), .O(n1220));
  LUT3 #(.INIT(8'hE8)) lut_n1221 (.I0(n1216), .I1(n1219), .I2(n1220), .O(n1221));
  LUT3 #(.INIT(8'hE8)) lut_n1222 (.I0(x276), .I1(x277), .I2(x278), .O(n1222));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1223 (.I0(x267), .I1(x268), .I2(x269), .I3(n1217), .I4(n1218), .O(n1223));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1224 (.I0(x273), .I1(x274), .I2(x275), .I3(n1222), .I4(n1223), .O(n1224));
  LUT3 #(.INIT(8'hE8)) lut_n1225 (.I0(x282), .I1(x283), .I2(x284), .O(n1225));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1226 (.I0(x273), .I1(x274), .I2(x275), .I3(n1222), .I4(n1223), .O(n1226));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1227 (.I0(x279), .I1(x280), .I2(x281), .I3(n1225), .I4(n1226), .O(n1227));
  LUT3 #(.INIT(8'h96)) lut_n1228 (.I0(n1216), .I1(n1219), .I2(n1220), .O(n1228));
  LUT3 #(.INIT(8'hE8)) lut_n1229 (.I0(n1224), .I1(n1227), .I2(n1228), .O(n1229));
  LUT3 #(.INIT(8'h96)) lut_n1230 (.I0(n1203), .I1(n1211), .I2(n1212), .O(n1230));
  LUT3 #(.INIT(8'hE8)) lut_n1231 (.I0(n1221), .I1(n1229), .I2(n1230), .O(n1231));
  LUT3 #(.INIT(8'h96)) lut_n1232 (.I0(n1175), .I1(n1193), .I2(n1194), .O(n1232));
  LUT3 #(.INIT(8'hE8)) lut_n1233 (.I0(n1213), .I1(n1231), .I2(n1232), .O(n1233));
  LUT3 #(.INIT(8'h96)) lut_n1234 (.I0(n1080), .I1(n1118), .I2(n1156), .O(n1234));
  LUT3 #(.INIT(8'hE8)) lut_n1235 (.I0(n1195), .I1(n1233), .I2(n1234), .O(n1235));
  LUT3 #(.INIT(8'hE8)) lut_n1236 (.I0(x288), .I1(x289), .I2(x290), .O(n1236));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1237 (.I0(x279), .I1(x280), .I2(x281), .I3(n1225), .I4(n1226), .O(n1237));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1238 (.I0(x285), .I1(x286), .I2(x287), .I3(n1236), .I4(n1237), .O(n1238));
  LUT3 #(.INIT(8'hE8)) lut_n1239 (.I0(x294), .I1(x295), .I2(x296), .O(n1239));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1240 (.I0(x285), .I1(x286), .I2(x287), .I3(n1236), .I4(n1237), .O(n1240));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1241 (.I0(x291), .I1(x292), .I2(x293), .I3(n1239), .I4(n1240), .O(n1241));
  LUT3 #(.INIT(8'h96)) lut_n1242 (.I0(n1224), .I1(n1227), .I2(n1228), .O(n1242));
  LUT3 #(.INIT(8'hE8)) lut_n1243 (.I0(n1238), .I1(n1241), .I2(n1242), .O(n1243));
  LUT3 #(.INIT(8'hE8)) lut_n1244 (.I0(x297), .I1(x298), .I2(x299), .O(n1244));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1245 (.I0(x291), .I1(x292), .I2(x293), .I3(n1239), .I4(n1240), .O(n1245));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1246 (.I0(x300), .I1(x301), .I2(x302), .I3(n1244), .I4(n1245), .O(n1246));
  LUT3 #(.INIT(8'hE8)) lut_n1247 (.I0(x306), .I1(x307), .I2(x308), .O(n1247));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1248 (.I0(x300), .I1(x301), .I2(x302), .I3(n1244), .I4(n1245), .O(n1248));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1249 (.I0(x303), .I1(x304), .I2(x305), .I3(n1247), .I4(n1248), .O(n1249));
  LUT3 #(.INIT(8'h96)) lut_n1250 (.I0(n1238), .I1(n1241), .I2(n1242), .O(n1250));
  LUT3 #(.INIT(8'hE8)) lut_n1251 (.I0(n1246), .I1(n1249), .I2(n1250), .O(n1251));
  LUT3 #(.INIT(8'h96)) lut_n1252 (.I0(n1221), .I1(n1229), .I2(n1230), .O(n1252));
  LUT3 #(.INIT(8'hE8)) lut_n1253 (.I0(n1243), .I1(n1251), .I2(n1252), .O(n1253));
  LUT3 #(.INIT(8'hE8)) lut_n1254 (.I0(x312), .I1(x313), .I2(x314), .O(n1254));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1255 (.I0(x303), .I1(x304), .I2(x305), .I3(n1247), .I4(n1248), .O(n1255));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1256 (.I0(x309), .I1(x310), .I2(x311), .I3(n1254), .I4(n1255), .O(n1256));
  LUT3 #(.INIT(8'hE8)) lut_n1257 (.I0(x318), .I1(x319), .I2(x320), .O(n1257));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1258 (.I0(x309), .I1(x310), .I2(x311), .I3(n1254), .I4(n1255), .O(n1258));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1259 (.I0(x315), .I1(x316), .I2(x317), .I3(n1257), .I4(n1258), .O(n1259));
  LUT3 #(.INIT(8'h96)) lut_n1260 (.I0(n1246), .I1(n1249), .I2(n1250), .O(n1260));
  LUT3 #(.INIT(8'hE8)) lut_n1261 (.I0(n1256), .I1(n1259), .I2(n1260), .O(n1261));
  LUT3 #(.INIT(8'hE8)) lut_n1262 (.I0(x324), .I1(x325), .I2(x326), .O(n1262));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1263 (.I0(x315), .I1(x316), .I2(x317), .I3(n1257), .I4(n1258), .O(n1263));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1264 (.I0(x321), .I1(x322), .I2(x323), .I3(n1262), .I4(n1263), .O(n1264));
  LUT3 #(.INIT(8'hE8)) lut_n1265 (.I0(x330), .I1(x331), .I2(x332), .O(n1265));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1266 (.I0(x321), .I1(x322), .I2(x323), .I3(n1262), .I4(n1263), .O(n1266));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1267 (.I0(x327), .I1(x328), .I2(x329), .I3(n1265), .I4(n1266), .O(n1267));
  LUT3 #(.INIT(8'h96)) lut_n1268 (.I0(n1256), .I1(n1259), .I2(n1260), .O(n1268));
  LUT3 #(.INIT(8'hE8)) lut_n1269 (.I0(n1264), .I1(n1267), .I2(n1268), .O(n1269));
  LUT3 #(.INIT(8'h96)) lut_n1270 (.I0(n1243), .I1(n1251), .I2(n1252), .O(n1270));
  LUT3 #(.INIT(8'hE8)) lut_n1271 (.I0(n1261), .I1(n1269), .I2(n1270), .O(n1271));
  LUT3 #(.INIT(8'h96)) lut_n1272 (.I0(n1213), .I1(n1231), .I2(n1232), .O(n1272));
  LUT3 #(.INIT(8'hE8)) lut_n1273 (.I0(n1253), .I1(n1271), .I2(n1272), .O(n1273));
  LUT3 #(.INIT(8'hE8)) lut_n1274 (.I0(x336), .I1(x337), .I2(x338), .O(n1274));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1275 (.I0(x327), .I1(x328), .I2(x329), .I3(n1265), .I4(n1266), .O(n1275));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1276 (.I0(x333), .I1(x334), .I2(x335), .I3(n1274), .I4(n1275), .O(n1276));
  LUT3 #(.INIT(8'hE8)) lut_n1277 (.I0(x342), .I1(x343), .I2(x344), .O(n1277));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1278 (.I0(x333), .I1(x334), .I2(x335), .I3(n1274), .I4(n1275), .O(n1278));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1279 (.I0(x339), .I1(x340), .I2(x341), .I3(n1277), .I4(n1278), .O(n1279));
  LUT3 #(.INIT(8'h96)) lut_n1280 (.I0(n1264), .I1(n1267), .I2(n1268), .O(n1280));
  LUT3 #(.INIT(8'hE8)) lut_n1281 (.I0(n1276), .I1(n1279), .I2(n1280), .O(n1281));
  LUT3 #(.INIT(8'hE8)) lut_n1282 (.I0(x348), .I1(x349), .I2(x350), .O(n1282));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1283 (.I0(x339), .I1(x340), .I2(x341), .I3(n1277), .I4(n1278), .O(n1283));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1284 (.I0(x345), .I1(x346), .I2(x347), .I3(n1282), .I4(n1283), .O(n1284));
  LUT3 #(.INIT(8'hE8)) lut_n1285 (.I0(x354), .I1(x355), .I2(x356), .O(n1285));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1286 (.I0(x345), .I1(x346), .I2(x347), .I3(n1282), .I4(n1283), .O(n1286));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1287 (.I0(x351), .I1(x352), .I2(x353), .I3(n1285), .I4(n1286), .O(n1287));
  LUT3 #(.INIT(8'h96)) lut_n1288 (.I0(n1276), .I1(n1279), .I2(n1280), .O(n1288));
  LUT3 #(.INIT(8'hE8)) lut_n1289 (.I0(n1284), .I1(n1287), .I2(n1288), .O(n1289));
  LUT3 #(.INIT(8'h96)) lut_n1290 (.I0(n1261), .I1(n1269), .I2(n1270), .O(n1290));
  LUT3 #(.INIT(8'hE8)) lut_n1291 (.I0(n1281), .I1(n1289), .I2(n1290), .O(n1291));
  LUT3 #(.INIT(8'hE8)) lut_n1292 (.I0(x360), .I1(x361), .I2(x362), .O(n1292));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1293 (.I0(x351), .I1(x352), .I2(x353), .I3(n1285), .I4(n1286), .O(n1293));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1294 (.I0(x357), .I1(x358), .I2(x359), .I3(n1292), .I4(n1293), .O(n1294));
  LUT3 #(.INIT(8'hE8)) lut_n1295 (.I0(x366), .I1(x367), .I2(x368), .O(n1295));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1296 (.I0(x357), .I1(x358), .I2(x359), .I3(n1292), .I4(n1293), .O(n1296));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1297 (.I0(x363), .I1(x364), .I2(x365), .I3(n1295), .I4(n1296), .O(n1297));
  LUT3 #(.INIT(8'h96)) lut_n1298 (.I0(n1284), .I1(n1287), .I2(n1288), .O(n1298));
  LUT3 #(.INIT(8'hE8)) lut_n1299 (.I0(n1294), .I1(n1297), .I2(n1298), .O(n1299));
  LUT3 #(.INIT(8'hE8)) lut_n1300 (.I0(x372), .I1(x373), .I2(x374), .O(n1300));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1301 (.I0(x363), .I1(x364), .I2(x365), .I3(n1295), .I4(n1296), .O(n1301));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1302 (.I0(x369), .I1(x370), .I2(x371), .I3(n1300), .I4(n1301), .O(n1302));
  LUT3 #(.INIT(8'hE8)) lut_n1303 (.I0(x378), .I1(x379), .I2(x380), .O(n1303));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1304 (.I0(x369), .I1(x370), .I2(x371), .I3(n1300), .I4(n1301), .O(n1304));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1305 (.I0(x375), .I1(x376), .I2(x377), .I3(n1303), .I4(n1304), .O(n1305));
  LUT3 #(.INIT(8'h96)) lut_n1306 (.I0(n1294), .I1(n1297), .I2(n1298), .O(n1306));
  LUT3 #(.INIT(8'hE8)) lut_n1307 (.I0(n1302), .I1(n1305), .I2(n1306), .O(n1307));
  LUT3 #(.INIT(8'h96)) lut_n1308 (.I0(n1281), .I1(n1289), .I2(n1290), .O(n1308));
  LUT3 #(.INIT(8'hE8)) lut_n1309 (.I0(n1299), .I1(n1307), .I2(n1308), .O(n1309));
  LUT3 #(.INIT(8'h96)) lut_n1310 (.I0(n1253), .I1(n1271), .I2(n1272), .O(n1310));
  LUT3 #(.INIT(8'hE8)) lut_n1311 (.I0(n1291), .I1(n1309), .I2(n1310), .O(n1311));
  LUT3 #(.INIT(8'h96)) lut_n1312 (.I0(n1195), .I1(n1233), .I2(n1234), .O(n1312));
  LUT3 #(.INIT(8'hE8)) lut_n1313 (.I0(n1273), .I1(n1311), .I2(n1312), .O(n1313));
  LUT3 #(.INIT(8'hE8)) lut_n1314 (.I0(n1157), .I1(n1235), .I2(n1313), .O(n1314));
  LUT3 #(.INIT(8'hE8)) lut_n1315 (.I0(x384), .I1(x385), .I2(x386), .O(n1315));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1316 (.I0(x375), .I1(x376), .I2(x377), .I3(n1303), .I4(n1304), .O(n1316));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1317 (.I0(x381), .I1(x382), .I2(x383), .I3(n1315), .I4(n1316), .O(n1317));
  LUT3 #(.INIT(8'hE8)) lut_n1318 (.I0(x390), .I1(x391), .I2(x392), .O(n1318));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1319 (.I0(x381), .I1(x382), .I2(x383), .I3(n1315), .I4(n1316), .O(n1319));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1320 (.I0(x387), .I1(x388), .I2(x389), .I3(n1318), .I4(n1319), .O(n1320));
  LUT3 #(.INIT(8'h96)) lut_n1321 (.I0(n1302), .I1(n1305), .I2(n1306), .O(n1321));
  LUT3 #(.INIT(8'hE8)) lut_n1322 (.I0(n1317), .I1(n1320), .I2(n1321), .O(n1322));
  LUT3 #(.INIT(8'hE8)) lut_n1323 (.I0(x396), .I1(x397), .I2(x398), .O(n1323));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1324 (.I0(x387), .I1(x388), .I2(x389), .I3(n1318), .I4(n1319), .O(n1324));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1325 (.I0(x393), .I1(x394), .I2(x395), .I3(n1323), .I4(n1324), .O(n1325));
  LUT3 #(.INIT(8'hE8)) lut_n1326 (.I0(x402), .I1(x403), .I2(x404), .O(n1326));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1327 (.I0(x393), .I1(x394), .I2(x395), .I3(n1323), .I4(n1324), .O(n1327));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1328 (.I0(x399), .I1(x400), .I2(x401), .I3(n1326), .I4(n1327), .O(n1328));
  LUT3 #(.INIT(8'h96)) lut_n1329 (.I0(n1317), .I1(n1320), .I2(n1321), .O(n1329));
  LUT3 #(.INIT(8'hE8)) lut_n1330 (.I0(n1325), .I1(n1328), .I2(n1329), .O(n1330));
  LUT3 #(.INIT(8'h96)) lut_n1331 (.I0(n1299), .I1(n1307), .I2(n1308), .O(n1331));
  LUT3 #(.INIT(8'hE8)) lut_n1332 (.I0(n1322), .I1(n1330), .I2(n1331), .O(n1332));
  LUT3 #(.INIT(8'hE8)) lut_n1333 (.I0(x408), .I1(x409), .I2(x410), .O(n1333));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1334 (.I0(x399), .I1(x400), .I2(x401), .I3(n1326), .I4(n1327), .O(n1334));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1335 (.I0(x405), .I1(x406), .I2(x407), .I3(n1333), .I4(n1334), .O(n1335));
  LUT3 #(.INIT(8'hE8)) lut_n1336 (.I0(x414), .I1(x415), .I2(x416), .O(n1336));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1337 (.I0(x405), .I1(x406), .I2(x407), .I3(n1333), .I4(n1334), .O(n1337));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1338 (.I0(x411), .I1(x412), .I2(x413), .I3(n1336), .I4(n1337), .O(n1338));
  LUT3 #(.INIT(8'h96)) lut_n1339 (.I0(n1325), .I1(n1328), .I2(n1329), .O(n1339));
  LUT3 #(.INIT(8'hE8)) lut_n1340 (.I0(n1335), .I1(n1338), .I2(n1339), .O(n1340));
  LUT3 #(.INIT(8'hE8)) lut_n1341 (.I0(x420), .I1(x421), .I2(x422), .O(n1341));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1342 (.I0(x411), .I1(x412), .I2(x413), .I3(n1336), .I4(n1337), .O(n1342));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1343 (.I0(x417), .I1(x418), .I2(x419), .I3(n1341), .I4(n1342), .O(n1343));
  LUT3 #(.INIT(8'hE8)) lut_n1344 (.I0(x426), .I1(x427), .I2(x428), .O(n1344));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1345 (.I0(x417), .I1(x418), .I2(x419), .I3(n1341), .I4(n1342), .O(n1345));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1346 (.I0(x423), .I1(x424), .I2(x425), .I3(n1344), .I4(n1345), .O(n1346));
  LUT3 #(.INIT(8'h96)) lut_n1347 (.I0(n1335), .I1(n1338), .I2(n1339), .O(n1347));
  LUT3 #(.INIT(8'hE8)) lut_n1348 (.I0(n1343), .I1(n1346), .I2(n1347), .O(n1348));
  LUT3 #(.INIT(8'h96)) lut_n1349 (.I0(n1322), .I1(n1330), .I2(n1331), .O(n1349));
  LUT3 #(.INIT(8'hE8)) lut_n1350 (.I0(n1340), .I1(n1348), .I2(n1349), .O(n1350));
  LUT3 #(.INIT(8'h96)) lut_n1351 (.I0(n1291), .I1(n1309), .I2(n1310), .O(n1351));
  LUT3 #(.INIT(8'hE8)) lut_n1352 (.I0(n1332), .I1(n1350), .I2(n1351), .O(n1352));
  LUT3 #(.INIT(8'hE8)) lut_n1353 (.I0(x432), .I1(x433), .I2(x434), .O(n1353));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1354 (.I0(x423), .I1(x424), .I2(x425), .I3(n1344), .I4(n1345), .O(n1354));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1355 (.I0(x429), .I1(x430), .I2(x431), .I3(n1353), .I4(n1354), .O(n1355));
  LUT3 #(.INIT(8'hE8)) lut_n1356 (.I0(x438), .I1(x439), .I2(x440), .O(n1356));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1357 (.I0(x429), .I1(x430), .I2(x431), .I3(n1353), .I4(n1354), .O(n1357));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1358 (.I0(x435), .I1(x436), .I2(x437), .I3(n1356), .I4(n1357), .O(n1358));
  LUT3 #(.INIT(8'h96)) lut_n1359 (.I0(n1343), .I1(n1346), .I2(n1347), .O(n1359));
  LUT3 #(.INIT(8'hE8)) lut_n1360 (.I0(n1355), .I1(n1358), .I2(n1359), .O(n1360));
  LUT3 #(.INIT(8'hE8)) lut_n1361 (.I0(x444), .I1(x445), .I2(x446), .O(n1361));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1362 (.I0(x435), .I1(x436), .I2(x437), .I3(n1356), .I4(n1357), .O(n1362));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1363 (.I0(x441), .I1(x442), .I2(x443), .I3(n1361), .I4(n1362), .O(n1363));
  LUT3 #(.INIT(8'hE8)) lut_n1364 (.I0(x450), .I1(x451), .I2(x452), .O(n1364));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1365 (.I0(x441), .I1(x442), .I2(x443), .I3(n1361), .I4(n1362), .O(n1365));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1366 (.I0(x447), .I1(x448), .I2(x449), .I3(n1364), .I4(n1365), .O(n1366));
  LUT3 #(.INIT(8'h96)) lut_n1367 (.I0(n1355), .I1(n1358), .I2(n1359), .O(n1367));
  LUT3 #(.INIT(8'hE8)) lut_n1368 (.I0(n1363), .I1(n1366), .I2(n1367), .O(n1368));
  LUT3 #(.INIT(8'h96)) lut_n1369 (.I0(n1340), .I1(n1348), .I2(n1349), .O(n1369));
  LUT3 #(.INIT(8'hE8)) lut_n1370 (.I0(n1360), .I1(n1368), .I2(n1369), .O(n1370));
  LUT3 #(.INIT(8'hE8)) lut_n1371 (.I0(x456), .I1(x457), .I2(x458), .O(n1371));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1372 (.I0(x447), .I1(x448), .I2(x449), .I3(n1364), .I4(n1365), .O(n1372));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1373 (.I0(x453), .I1(x454), .I2(x455), .I3(n1371), .I4(n1372), .O(n1373));
  LUT3 #(.INIT(8'hE8)) lut_n1374 (.I0(x462), .I1(x463), .I2(x464), .O(n1374));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1375 (.I0(x453), .I1(x454), .I2(x455), .I3(n1371), .I4(n1372), .O(n1375));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1376 (.I0(x459), .I1(x460), .I2(x461), .I3(n1374), .I4(n1375), .O(n1376));
  LUT3 #(.INIT(8'h96)) lut_n1377 (.I0(n1363), .I1(n1366), .I2(n1367), .O(n1377));
  LUT3 #(.INIT(8'hE8)) lut_n1378 (.I0(n1373), .I1(n1376), .I2(n1377), .O(n1378));
  LUT3 #(.INIT(8'hE8)) lut_n1379 (.I0(x468), .I1(x469), .I2(x470), .O(n1379));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1380 (.I0(x459), .I1(x460), .I2(x461), .I3(n1374), .I4(n1375), .O(n1380));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1381 (.I0(x465), .I1(x466), .I2(x467), .I3(n1379), .I4(n1380), .O(n1381));
  LUT3 #(.INIT(8'hE8)) lut_n1382 (.I0(x474), .I1(x475), .I2(x476), .O(n1382));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1383 (.I0(x465), .I1(x466), .I2(x467), .I3(n1379), .I4(n1380), .O(n1383));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1384 (.I0(x471), .I1(x472), .I2(x473), .I3(n1382), .I4(n1383), .O(n1384));
  LUT3 #(.INIT(8'h96)) lut_n1385 (.I0(n1373), .I1(n1376), .I2(n1377), .O(n1385));
  LUT3 #(.INIT(8'hE8)) lut_n1386 (.I0(n1381), .I1(n1384), .I2(n1385), .O(n1386));
  LUT3 #(.INIT(8'h96)) lut_n1387 (.I0(n1360), .I1(n1368), .I2(n1369), .O(n1387));
  LUT3 #(.INIT(8'hE8)) lut_n1388 (.I0(n1378), .I1(n1386), .I2(n1387), .O(n1388));
  LUT3 #(.INIT(8'h96)) lut_n1389 (.I0(n1332), .I1(n1350), .I2(n1351), .O(n1389));
  LUT3 #(.INIT(8'hE8)) lut_n1390 (.I0(n1370), .I1(n1388), .I2(n1389), .O(n1390));
  LUT3 #(.INIT(8'h96)) lut_n1391 (.I0(n1273), .I1(n1311), .I2(n1312), .O(n1391));
  LUT3 #(.INIT(8'hE8)) lut_n1392 (.I0(n1352), .I1(n1390), .I2(n1391), .O(n1392));
  LUT3 #(.INIT(8'hE8)) lut_n1393 (.I0(x480), .I1(x481), .I2(x482), .O(n1393));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1394 (.I0(x471), .I1(x472), .I2(x473), .I3(n1382), .I4(n1383), .O(n1394));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1395 (.I0(x477), .I1(x478), .I2(x479), .I3(n1393), .I4(n1394), .O(n1395));
  LUT3 #(.INIT(8'hE8)) lut_n1396 (.I0(x486), .I1(x487), .I2(x488), .O(n1396));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1397 (.I0(x477), .I1(x478), .I2(x479), .I3(n1393), .I4(n1394), .O(n1397));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1398 (.I0(x483), .I1(x484), .I2(x485), .I3(n1396), .I4(n1397), .O(n1398));
  LUT3 #(.INIT(8'h96)) lut_n1399 (.I0(n1381), .I1(n1384), .I2(n1385), .O(n1399));
  LUT3 #(.INIT(8'hE8)) lut_n1400 (.I0(n1395), .I1(n1398), .I2(n1399), .O(n1400));
  LUT3 #(.INIT(8'hE8)) lut_n1401 (.I0(x492), .I1(x493), .I2(x494), .O(n1401));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1402 (.I0(x483), .I1(x484), .I2(x485), .I3(n1396), .I4(n1397), .O(n1402));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1403 (.I0(x489), .I1(x490), .I2(x491), .I3(n1401), .I4(n1402), .O(n1403));
  LUT3 #(.INIT(8'hE8)) lut_n1404 (.I0(x498), .I1(x499), .I2(x500), .O(n1404));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1405 (.I0(x489), .I1(x490), .I2(x491), .I3(n1401), .I4(n1402), .O(n1405));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1406 (.I0(x495), .I1(x496), .I2(x497), .I3(n1404), .I4(n1405), .O(n1406));
  LUT3 #(.INIT(8'h96)) lut_n1407 (.I0(n1395), .I1(n1398), .I2(n1399), .O(n1407));
  LUT3 #(.INIT(8'hE8)) lut_n1408 (.I0(n1403), .I1(n1406), .I2(n1407), .O(n1408));
  LUT3 #(.INIT(8'h96)) lut_n1409 (.I0(n1378), .I1(n1386), .I2(n1387), .O(n1409));
  LUT3 #(.INIT(8'hE8)) lut_n1410 (.I0(n1400), .I1(n1408), .I2(n1409), .O(n1410));
  LUT3 #(.INIT(8'hE8)) lut_n1411 (.I0(x504), .I1(x505), .I2(x506), .O(n1411));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1412 (.I0(x495), .I1(x496), .I2(x497), .I3(n1404), .I4(n1405), .O(n1412));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1413 (.I0(x501), .I1(x502), .I2(x503), .I3(n1411), .I4(n1412), .O(n1413));
  LUT3 #(.INIT(8'hE8)) lut_n1414 (.I0(x510), .I1(x511), .I2(x512), .O(n1414));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1415 (.I0(x501), .I1(x502), .I2(x503), .I3(n1411), .I4(n1412), .O(n1415));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1416 (.I0(x507), .I1(x508), .I2(x509), .I3(n1414), .I4(n1415), .O(n1416));
  LUT3 #(.INIT(8'h96)) lut_n1417 (.I0(n1403), .I1(n1406), .I2(n1407), .O(n1417));
  LUT3 #(.INIT(8'hE8)) lut_n1418 (.I0(n1413), .I1(n1416), .I2(n1417), .O(n1418));
  LUT3 #(.INIT(8'hE8)) lut_n1419 (.I0(x516), .I1(x517), .I2(x518), .O(n1419));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1420 (.I0(x507), .I1(x508), .I2(x509), .I3(n1414), .I4(n1415), .O(n1420));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1421 (.I0(x513), .I1(x514), .I2(x515), .I3(n1419), .I4(n1420), .O(n1421));
  LUT3 #(.INIT(8'hE8)) lut_n1422 (.I0(x522), .I1(x523), .I2(x524), .O(n1422));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1423 (.I0(x513), .I1(x514), .I2(x515), .I3(n1419), .I4(n1420), .O(n1423));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1424 (.I0(x519), .I1(x520), .I2(x521), .I3(n1422), .I4(n1423), .O(n1424));
  LUT3 #(.INIT(8'h96)) lut_n1425 (.I0(n1413), .I1(n1416), .I2(n1417), .O(n1425));
  LUT3 #(.INIT(8'hE8)) lut_n1426 (.I0(n1421), .I1(n1424), .I2(n1425), .O(n1426));
  LUT3 #(.INIT(8'h96)) lut_n1427 (.I0(n1400), .I1(n1408), .I2(n1409), .O(n1427));
  LUT3 #(.INIT(8'hE8)) lut_n1428 (.I0(n1418), .I1(n1426), .I2(n1427), .O(n1428));
  LUT3 #(.INIT(8'h96)) lut_n1429 (.I0(n1370), .I1(n1388), .I2(n1389), .O(n1429));
  LUT3 #(.INIT(8'hE8)) lut_n1430 (.I0(n1410), .I1(n1428), .I2(n1429), .O(n1430));
  LUT3 #(.INIT(8'hE8)) lut_n1431 (.I0(x528), .I1(x529), .I2(x530), .O(n1431));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1432 (.I0(x519), .I1(x520), .I2(x521), .I3(n1422), .I4(n1423), .O(n1432));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1433 (.I0(x525), .I1(x526), .I2(x527), .I3(n1431), .I4(n1432), .O(n1433));
  LUT3 #(.INIT(8'hE8)) lut_n1434 (.I0(x534), .I1(x535), .I2(x536), .O(n1434));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1435 (.I0(x525), .I1(x526), .I2(x527), .I3(n1431), .I4(n1432), .O(n1435));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1436 (.I0(x531), .I1(x532), .I2(x533), .I3(n1434), .I4(n1435), .O(n1436));
  LUT3 #(.INIT(8'h96)) lut_n1437 (.I0(n1421), .I1(n1424), .I2(n1425), .O(n1437));
  LUT3 #(.INIT(8'hE8)) lut_n1438 (.I0(n1433), .I1(n1436), .I2(n1437), .O(n1438));
  LUT3 #(.INIT(8'hE8)) lut_n1439 (.I0(x540), .I1(x541), .I2(x542), .O(n1439));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1440 (.I0(x531), .I1(x532), .I2(x533), .I3(n1434), .I4(n1435), .O(n1440));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1441 (.I0(x537), .I1(x538), .I2(x539), .I3(n1439), .I4(n1440), .O(n1441));
  LUT3 #(.INIT(8'hE8)) lut_n1442 (.I0(x546), .I1(x547), .I2(x548), .O(n1442));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1443 (.I0(x537), .I1(x538), .I2(x539), .I3(n1439), .I4(n1440), .O(n1443));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1444 (.I0(x543), .I1(x544), .I2(x545), .I3(n1442), .I4(n1443), .O(n1444));
  LUT3 #(.INIT(8'h96)) lut_n1445 (.I0(n1433), .I1(n1436), .I2(n1437), .O(n1445));
  LUT3 #(.INIT(8'hE8)) lut_n1446 (.I0(n1441), .I1(n1444), .I2(n1445), .O(n1446));
  LUT3 #(.INIT(8'h96)) lut_n1447 (.I0(n1418), .I1(n1426), .I2(n1427), .O(n1447));
  LUT3 #(.INIT(8'hE8)) lut_n1448 (.I0(n1438), .I1(n1446), .I2(n1447), .O(n1448));
  LUT3 #(.INIT(8'hE8)) lut_n1449 (.I0(x552), .I1(x553), .I2(x554), .O(n1449));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1450 (.I0(x543), .I1(x544), .I2(x545), .I3(n1442), .I4(n1443), .O(n1450));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1451 (.I0(x549), .I1(x550), .I2(x551), .I3(n1449), .I4(n1450), .O(n1451));
  LUT3 #(.INIT(8'hE8)) lut_n1452 (.I0(x558), .I1(x559), .I2(x560), .O(n1452));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1453 (.I0(x549), .I1(x550), .I2(x551), .I3(n1449), .I4(n1450), .O(n1453));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1454 (.I0(x555), .I1(x556), .I2(x557), .I3(n1452), .I4(n1453), .O(n1454));
  LUT3 #(.INIT(8'h96)) lut_n1455 (.I0(n1441), .I1(n1444), .I2(n1445), .O(n1455));
  LUT3 #(.INIT(8'hE8)) lut_n1456 (.I0(n1451), .I1(n1454), .I2(n1455), .O(n1456));
  LUT3 #(.INIT(8'hE8)) lut_n1457 (.I0(x564), .I1(x565), .I2(x566), .O(n1457));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1458 (.I0(x555), .I1(x556), .I2(x557), .I3(n1452), .I4(n1453), .O(n1458));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1459 (.I0(x561), .I1(x562), .I2(x563), .I3(n1457), .I4(n1458), .O(n1459));
  LUT3 #(.INIT(8'hE8)) lut_n1460 (.I0(x570), .I1(x571), .I2(x572), .O(n1460));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1461 (.I0(x561), .I1(x562), .I2(x563), .I3(n1457), .I4(n1458), .O(n1461));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1462 (.I0(x567), .I1(x568), .I2(x569), .I3(n1460), .I4(n1461), .O(n1462));
  LUT3 #(.INIT(8'h96)) lut_n1463 (.I0(n1451), .I1(n1454), .I2(n1455), .O(n1463));
  LUT3 #(.INIT(8'hE8)) lut_n1464 (.I0(n1459), .I1(n1462), .I2(n1463), .O(n1464));
  LUT3 #(.INIT(8'h96)) lut_n1465 (.I0(n1438), .I1(n1446), .I2(n1447), .O(n1465));
  LUT3 #(.INIT(8'hE8)) lut_n1466 (.I0(n1456), .I1(n1464), .I2(n1465), .O(n1466));
  LUT3 #(.INIT(8'h96)) lut_n1467 (.I0(n1410), .I1(n1428), .I2(n1429), .O(n1467));
  LUT3 #(.INIT(8'hE8)) lut_n1468 (.I0(n1448), .I1(n1466), .I2(n1467), .O(n1468));
  LUT3 #(.INIT(8'h96)) lut_n1469 (.I0(n1352), .I1(n1390), .I2(n1391), .O(n1469));
  LUT3 #(.INIT(8'hE8)) lut_n1470 (.I0(n1430), .I1(n1468), .I2(n1469), .O(n1470));
  LUT3 #(.INIT(8'h96)) lut_n1471 (.I0(n1157), .I1(n1235), .I2(n1313), .O(n1471));
  LUT3 #(.INIT(8'hE8)) lut_n1472 (.I0(n1392), .I1(n1470), .I2(n1471), .O(n1472));
  LUT3 #(.INIT(8'hE8)) lut_n1473 (.I0(x576), .I1(x577), .I2(x578), .O(n1473));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1474 (.I0(x567), .I1(x568), .I2(x569), .I3(n1460), .I4(n1461), .O(n1474));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1475 (.I0(x573), .I1(x574), .I2(x575), .I3(n1473), .I4(n1474), .O(n1475));
  LUT3 #(.INIT(8'hE8)) lut_n1476 (.I0(x582), .I1(x583), .I2(x584), .O(n1476));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1477 (.I0(x573), .I1(x574), .I2(x575), .I3(n1473), .I4(n1474), .O(n1477));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1478 (.I0(x579), .I1(x580), .I2(x581), .I3(n1476), .I4(n1477), .O(n1478));
  LUT3 #(.INIT(8'h96)) lut_n1479 (.I0(n1459), .I1(n1462), .I2(n1463), .O(n1479));
  LUT3 #(.INIT(8'hE8)) lut_n1480 (.I0(n1475), .I1(n1478), .I2(n1479), .O(n1480));
  LUT3 #(.INIT(8'hE8)) lut_n1481 (.I0(x588), .I1(x589), .I2(x590), .O(n1481));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1482 (.I0(x579), .I1(x580), .I2(x581), .I3(n1476), .I4(n1477), .O(n1482));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1483 (.I0(x585), .I1(x586), .I2(x587), .I3(n1481), .I4(n1482), .O(n1483));
  LUT3 #(.INIT(8'hE8)) lut_n1484 (.I0(x594), .I1(x595), .I2(x596), .O(n1484));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1485 (.I0(x585), .I1(x586), .I2(x587), .I3(n1481), .I4(n1482), .O(n1485));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1486 (.I0(x591), .I1(x592), .I2(x593), .I3(n1484), .I4(n1485), .O(n1486));
  LUT3 #(.INIT(8'h96)) lut_n1487 (.I0(n1475), .I1(n1478), .I2(n1479), .O(n1487));
  LUT3 #(.INIT(8'hE8)) lut_n1488 (.I0(n1483), .I1(n1486), .I2(n1487), .O(n1488));
  LUT3 #(.INIT(8'h96)) lut_n1489 (.I0(n1456), .I1(n1464), .I2(n1465), .O(n1489));
  LUT3 #(.INIT(8'hE8)) lut_n1490 (.I0(n1480), .I1(n1488), .I2(n1489), .O(n1490));
  LUT3 #(.INIT(8'hE8)) lut_n1491 (.I0(x600), .I1(x601), .I2(x602), .O(n1491));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1492 (.I0(x591), .I1(x592), .I2(x593), .I3(n1484), .I4(n1485), .O(n1492));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1493 (.I0(x597), .I1(x598), .I2(x599), .I3(n1491), .I4(n1492), .O(n1493));
  LUT3 #(.INIT(8'hE8)) lut_n1494 (.I0(x606), .I1(x607), .I2(x608), .O(n1494));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1495 (.I0(x597), .I1(x598), .I2(x599), .I3(n1491), .I4(n1492), .O(n1495));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1496 (.I0(x603), .I1(x604), .I2(x605), .I3(n1494), .I4(n1495), .O(n1496));
  LUT3 #(.INIT(8'h96)) lut_n1497 (.I0(n1483), .I1(n1486), .I2(n1487), .O(n1497));
  LUT3 #(.INIT(8'hE8)) lut_n1498 (.I0(n1493), .I1(n1496), .I2(n1497), .O(n1498));
  LUT3 #(.INIT(8'hE8)) lut_n1499 (.I0(x612), .I1(x613), .I2(x614), .O(n1499));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1500 (.I0(x603), .I1(x604), .I2(x605), .I3(n1494), .I4(n1495), .O(n1500));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1501 (.I0(x609), .I1(x610), .I2(x611), .I3(n1499), .I4(n1500), .O(n1501));
  LUT3 #(.INIT(8'hE8)) lut_n1502 (.I0(x618), .I1(x619), .I2(x620), .O(n1502));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1503 (.I0(x609), .I1(x610), .I2(x611), .I3(n1499), .I4(n1500), .O(n1503));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1504 (.I0(x615), .I1(x616), .I2(x617), .I3(n1502), .I4(n1503), .O(n1504));
  LUT3 #(.INIT(8'h96)) lut_n1505 (.I0(n1493), .I1(n1496), .I2(n1497), .O(n1505));
  LUT3 #(.INIT(8'hE8)) lut_n1506 (.I0(n1501), .I1(n1504), .I2(n1505), .O(n1506));
  LUT3 #(.INIT(8'h96)) lut_n1507 (.I0(n1480), .I1(n1488), .I2(n1489), .O(n1507));
  LUT3 #(.INIT(8'hE8)) lut_n1508 (.I0(n1498), .I1(n1506), .I2(n1507), .O(n1508));
  LUT3 #(.INIT(8'h96)) lut_n1509 (.I0(n1448), .I1(n1466), .I2(n1467), .O(n1509));
  LUT3 #(.INIT(8'hE8)) lut_n1510 (.I0(n1490), .I1(n1508), .I2(n1509), .O(n1510));
  LUT3 #(.INIT(8'hE8)) lut_n1511 (.I0(x624), .I1(x625), .I2(x626), .O(n1511));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1512 (.I0(x615), .I1(x616), .I2(x617), .I3(n1502), .I4(n1503), .O(n1512));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1513 (.I0(x621), .I1(x622), .I2(x623), .I3(n1511), .I4(n1512), .O(n1513));
  LUT3 #(.INIT(8'hE8)) lut_n1514 (.I0(x630), .I1(x631), .I2(x632), .O(n1514));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1515 (.I0(x621), .I1(x622), .I2(x623), .I3(n1511), .I4(n1512), .O(n1515));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1516 (.I0(x627), .I1(x628), .I2(x629), .I3(n1514), .I4(n1515), .O(n1516));
  LUT3 #(.INIT(8'h96)) lut_n1517 (.I0(n1501), .I1(n1504), .I2(n1505), .O(n1517));
  LUT3 #(.INIT(8'hE8)) lut_n1518 (.I0(n1513), .I1(n1516), .I2(n1517), .O(n1518));
  LUT3 #(.INIT(8'hE8)) lut_n1519 (.I0(x636), .I1(x637), .I2(x638), .O(n1519));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1520 (.I0(x627), .I1(x628), .I2(x629), .I3(n1514), .I4(n1515), .O(n1520));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1521 (.I0(x633), .I1(x634), .I2(x635), .I3(n1519), .I4(n1520), .O(n1521));
  LUT3 #(.INIT(8'hE8)) lut_n1522 (.I0(x642), .I1(x643), .I2(x644), .O(n1522));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1523 (.I0(x633), .I1(x634), .I2(x635), .I3(n1519), .I4(n1520), .O(n1523));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1524 (.I0(x639), .I1(x640), .I2(x641), .I3(n1522), .I4(n1523), .O(n1524));
  LUT3 #(.INIT(8'h96)) lut_n1525 (.I0(n1513), .I1(n1516), .I2(n1517), .O(n1525));
  LUT3 #(.INIT(8'hE8)) lut_n1526 (.I0(n1521), .I1(n1524), .I2(n1525), .O(n1526));
  LUT3 #(.INIT(8'h96)) lut_n1527 (.I0(n1498), .I1(n1506), .I2(n1507), .O(n1527));
  LUT3 #(.INIT(8'hE8)) lut_n1528 (.I0(n1518), .I1(n1526), .I2(n1527), .O(n1528));
  LUT3 #(.INIT(8'hE8)) lut_n1529 (.I0(x648), .I1(x649), .I2(x650), .O(n1529));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1530 (.I0(x639), .I1(x640), .I2(x641), .I3(n1522), .I4(n1523), .O(n1530));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1531 (.I0(x645), .I1(x646), .I2(x647), .I3(n1529), .I4(n1530), .O(n1531));
  LUT3 #(.INIT(8'hE8)) lut_n1532 (.I0(x654), .I1(x655), .I2(x656), .O(n1532));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1533 (.I0(x645), .I1(x646), .I2(x647), .I3(n1529), .I4(n1530), .O(n1533));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1534 (.I0(x651), .I1(x652), .I2(x653), .I3(n1532), .I4(n1533), .O(n1534));
  LUT3 #(.INIT(8'h96)) lut_n1535 (.I0(n1521), .I1(n1524), .I2(n1525), .O(n1535));
  LUT3 #(.INIT(8'hE8)) lut_n1536 (.I0(n1531), .I1(n1534), .I2(n1535), .O(n1536));
  LUT3 #(.INIT(8'hE8)) lut_n1537 (.I0(x660), .I1(x661), .I2(x662), .O(n1537));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1538 (.I0(x651), .I1(x652), .I2(x653), .I3(n1532), .I4(n1533), .O(n1538));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1539 (.I0(x657), .I1(x658), .I2(x659), .I3(n1537), .I4(n1538), .O(n1539));
  LUT3 #(.INIT(8'hE8)) lut_n1540 (.I0(x666), .I1(x667), .I2(x668), .O(n1540));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1541 (.I0(x657), .I1(x658), .I2(x659), .I3(n1537), .I4(n1538), .O(n1541));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1542 (.I0(x663), .I1(x664), .I2(x665), .I3(n1540), .I4(n1541), .O(n1542));
  LUT3 #(.INIT(8'h96)) lut_n1543 (.I0(n1531), .I1(n1534), .I2(n1535), .O(n1543));
  LUT3 #(.INIT(8'hE8)) lut_n1544 (.I0(n1539), .I1(n1542), .I2(n1543), .O(n1544));
  LUT3 #(.INIT(8'h96)) lut_n1545 (.I0(n1518), .I1(n1526), .I2(n1527), .O(n1545));
  LUT3 #(.INIT(8'hE8)) lut_n1546 (.I0(n1536), .I1(n1544), .I2(n1545), .O(n1546));
  LUT3 #(.INIT(8'h96)) lut_n1547 (.I0(n1490), .I1(n1508), .I2(n1509), .O(n1547));
  LUT3 #(.INIT(8'hE8)) lut_n1548 (.I0(n1528), .I1(n1546), .I2(n1547), .O(n1548));
  LUT3 #(.INIT(8'h96)) lut_n1549 (.I0(n1430), .I1(n1468), .I2(n1469), .O(n1549));
  LUT3 #(.INIT(8'hE8)) lut_n1550 (.I0(n1510), .I1(n1548), .I2(n1549), .O(n1550));
  LUT3 #(.INIT(8'hE8)) lut_n1551 (.I0(x672), .I1(x673), .I2(x674), .O(n1551));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1552 (.I0(x663), .I1(x664), .I2(x665), .I3(n1540), .I4(n1541), .O(n1552));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1553 (.I0(x669), .I1(x670), .I2(x671), .I3(n1551), .I4(n1552), .O(n1553));
  LUT3 #(.INIT(8'hE8)) lut_n1554 (.I0(x678), .I1(x679), .I2(x680), .O(n1554));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1555 (.I0(x669), .I1(x670), .I2(x671), .I3(n1551), .I4(n1552), .O(n1555));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1556 (.I0(x675), .I1(x676), .I2(x677), .I3(n1554), .I4(n1555), .O(n1556));
  LUT3 #(.INIT(8'h96)) lut_n1557 (.I0(n1539), .I1(n1542), .I2(n1543), .O(n1557));
  LUT3 #(.INIT(8'hE8)) lut_n1558 (.I0(n1553), .I1(n1556), .I2(n1557), .O(n1558));
  LUT3 #(.INIT(8'hE8)) lut_n1559 (.I0(x684), .I1(x685), .I2(x686), .O(n1559));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1560 (.I0(x675), .I1(x676), .I2(x677), .I3(n1554), .I4(n1555), .O(n1560));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1561 (.I0(x681), .I1(x682), .I2(x683), .I3(n1559), .I4(n1560), .O(n1561));
  LUT3 #(.INIT(8'hE8)) lut_n1562 (.I0(x690), .I1(x691), .I2(x692), .O(n1562));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1563 (.I0(x681), .I1(x682), .I2(x683), .I3(n1559), .I4(n1560), .O(n1563));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1564 (.I0(x687), .I1(x688), .I2(x689), .I3(n1562), .I4(n1563), .O(n1564));
  LUT3 #(.INIT(8'h96)) lut_n1565 (.I0(n1553), .I1(n1556), .I2(n1557), .O(n1565));
  LUT3 #(.INIT(8'hE8)) lut_n1566 (.I0(n1561), .I1(n1564), .I2(n1565), .O(n1566));
  LUT3 #(.INIT(8'h96)) lut_n1567 (.I0(n1536), .I1(n1544), .I2(n1545), .O(n1567));
  LUT3 #(.INIT(8'hE8)) lut_n1568 (.I0(n1558), .I1(n1566), .I2(n1567), .O(n1568));
  LUT3 #(.INIT(8'hE8)) lut_n1569 (.I0(x696), .I1(x697), .I2(x698), .O(n1569));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1570 (.I0(x687), .I1(x688), .I2(x689), .I3(n1562), .I4(n1563), .O(n1570));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1571 (.I0(x693), .I1(x694), .I2(x695), .I3(n1569), .I4(n1570), .O(n1571));
  LUT3 #(.INIT(8'hE8)) lut_n1572 (.I0(x702), .I1(x703), .I2(x704), .O(n1572));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1573 (.I0(x693), .I1(x694), .I2(x695), .I3(n1569), .I4(n1570), .O(n1573));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1574 (.I0(x699), .I1(x700), .I2(x701), .I3(n1572), .I4(n1573), .O(n1574));
  LUT3 #(.INIT(8'h96)) lut_n1575 (.I0(n1561), .I1(n1564), .I2(n1565), .O(n1575));
  LUT3 #(.INIT(8'hE8)) lut_n1576 (.I0(n1571), .I1(n1574), .I2(n1575), .O(n1576));
  LUT3 #(.INIT(8'hE8)) lut_n1577 (.I0(x708), .I1(x709), .I2(x710), .O(n1577));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1578 (.I0(x699), .I1(x700), .I2(x701), .I3(n1572), .I4(n1573), .O(n1578));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1579 (.I0(x705), .I1(x706), .I2(x707), .I3(n1577), .I4(n1578), .O(n1579));
  LUT3 #(.INIT(8'hE8)) lut_n1580 (.I0(x714), .I1(x715), .I2(x716), .O(n1580));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1581 (.I0(x705), .I1(x706), .I2(x707), .I3(n1577), .I4(n1578), .O(n1581));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1582 (.I0(x711), .I1(x712), .I2(x713), .I3(n1580), .I4(n1581), .O(n1582));
  LUT3 #(.INIT(8'h96)) lut_n1583 (.I0(n1571), .I1(n1574), .I2(n1575), .O(n1583));
  LUT3 #(.INIT(8'hE8)) lut_n1584 (.I0(n1579), .I1(n1582), .I2(n1583), .O(n1584));
  LUT3 #(.INIT(8'h96)) lut_n1585 (.I0(n1558), .I1(n1566), .I2(n1567), .O(n1585));
  LUT3 #(.INIT(8'hE8)) lut_n1586 (.I0(n1576), .I1(n1584), .I2(n1585), .O(n1586));
  LUT3 #(.INIT(8'h96)) lut_n1587 (.I0(n1528), .I1(n1546), .I2(n1547), .O(n1587));
  LUT3 #(.INIT(8'hE8)) lut_n1588 (.I0(n1568), .I1(n1586), .I2(n1587), .O(n1588));
  LUT3 #(.INIT(8'hE8)) lut_n1589 (.I0(x720), .I1(x721), .I2(x722), .O(n1589));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1590 (.I0(x711), .I1(x712), .I2(x713), .I3(n1580), .I4(n1581), .O(n1590));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1591 (.I0(x717), .I1(x718), .I2(x719), .I3(n1589), .I4(n1590), .O(n1591));
  LUT3 #(.INIT(8'hE8)) lut_n1592 (.I0(x726), .I1(x727), .I2(x728), .O(n1592));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1593 (.I0(x717), .I1(x718), .I2(x719), .I3(n1589), .I4(n1590), .O(n1593));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1594 (.I0(x723), .I1(x724), .I2(x725), .I3(n1592), .I4(n1593), .O(n1594));
  LUT3 #(.INIT(8'h96)) lut_n1595 (.I0(n1579), .I1(n1582), .I2(n1583), .O(n1595));
  LUT3 #(.INIT(8'hE8)) lut_n1596 (.I0(n1591), .I1(n1594), .I2(n1595), .O(n1596));
  LUT3 #(.INIT(8'hE8)) lut_n1597 (.I0(x732), .I1(x733), .I2(x734), .O(n1597));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1598 (.I0(x723), .I1(x724), .I2(x725), .I3(n1592), .I4(n1593), .O(n1598));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1599 (.I0(x729), .I1(x730), .I2(x731), .I3(n1597), .I4(n1598), .O(n1599));
  LUT3 #(.INIT(8'hE8)) lut_n1600 (.I0(x738), .I1(x739), .I2(x740), .O(n1600));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1601 (.I0(x729), .I1(x730), .I2(x731), .I3(n1597), .I4(n1598), .O(n1601));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1602 (.I0(x735), .I1(x736), .I2(x737), .I3(n1600), .I4(n1601), .O(n1602));
  LUT3 #(.INIT(8'h96)) lut_n1603 (.I0(n1591), .I1(n1594), .I2(n1595), .O(n1603));
  LUT3 #(.INIT(8'hE8)) lut_n1604 (.I0(n1599), .I1(n1602), .I2(n1603), .O(n1604));
  LUT3 #(.INIT(8'h96)) lut_n1605 (.I0(n1576), .I1(n1584), .I2(n1585), .O(n1605));
  LUT3 #(.INIT(8'hE8)) lut_n1606 (.I0(n1596), .I1(n1604), .I2(n1605), .O(n1606));
  LUT3 #(.INIT(8'hE8)) lut_n1607 (.I0(x744), .I1(x745), .I2(x746), .O(n1607));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1608 (.I0(x735), .I1(x736), .I2(x737), .I3(n1600), .I4(n1601), .O(n1608));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1609 (.I0(x741), .I1(x742), .I2(x743), .I3(n1607), .I4(n1608), .O(n1609));
  LUT3 #(.INIT(8'hE8)) lut_n1610 (.I0(x750), .I1(x751), .I2(x752), .O(n1610));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1611 (.I0(x741), .I1(x742), .I2(x743), .I3(n1607), .I4(n1608), .O(n1611));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1612 (.I0(x747), .I1(x748), .I2(x749), .I3(n1610), .I4(n1611), .O(n1612));
  LUT3 #(.INIT(8'h96)) lut_n1613 (.I0(n1599), .I1(n1602), .I2(n1603), .O(n1613));
  LUT3 #(.INIT(8'hE8)) lut_n1614 (.I0(n1609), .I1(n1612), .I2(n1613), .O(n1614));
  LUT3 #(.INIT(8'hE8)) lut_n1615 (.I0(x756), .I1(x757), .I2(x758), .O(n1615));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1616 (.I0(x747), .I1(x748), .I2(x749), .I3(n1610), .I4(n1611), .O(n1616));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1617 (.I0(x753), .I1(x754), .I2(x755), .I3(n1615), .I4(n1616), .O(n1617));
  LUT3 #(.INIT(8'hE8)) lut_n1618 (.I0(x762), .I1(x763), .I2(x764), .O(n1618));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1619 (.I0(x753), .I1(x754), .I2(x755), .I3(n1615), .I4(n1616), .O(n1619));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1620 (.I0(x759), .I1(x760), .I2(x761), .I3(n1618), .I4(n1619), .O(n1620));
  LUT3 #(.INIT(8'h96)) lut_n1621 (.I0(n1609), .I1(n1612), .I2(n1613), .O(n1621));
  LUT3 #(.INIT(8'hE8)) lut_n1622 (.I0(n1617), .I1(n1620), .I2(n1621), .O(n1622));
  LUT3 #(.INIT(8'h96)) lut_n1623 (.I0(n1596), .I1(n1604), .I2(n1605), .O(n1623));
  LUT3 #(.INIT(8'hE8)) lut_n1624 (.I0(n1614), .I1(n1622), .I2(n1623), .O(n1624));
  LUT3 #(.INIT(8'h96)) lut_n1625 (.I0(n1568), .I1(n1586), .I2(n1587), .O(n1625));
  LUT3 #(.INIT(8'hE8)) lut_n1626 (.I0(n1606), .I1(n1624), .I2(n1625), .O(n1626));
  LUT3 #(.INIT(8'h96)) lut_n1627 (.I0(n1510), .I1(n1548), .I2(n1549), .O(n1627));
  LUT3 #(.INIT(8'hE8)) lut_n1628 (.I0(n1588), .I1(n1626), .I2(n1627), .O(n1628));
  LUT3 #(.INIT(8'h96)) lut_n1629 (.I0(n1392), .I1(n1470), .I2(n1471), .O(n1629));
  LUT3 #(.INIT(8'hE8)) lut_n1630 (.I0(n1550), .I1(n1628), .I2(n1629), .O(n1630));
  LUT3 #(.INIT(8'hE8)) lut_n1631 (.I0(x768), .I1(x769), .I2(x770), .O(n1631));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1632 (.I0(x759), .I1(x760), .I2(x761), .I3(n1618), .I4(n1619), .O(n1632));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1633 (.I0(x765), .I1(x766), .I2(x767), .I3(n1631), .I4(n1632), .O(n1633));
  LUT3 #(.INIT(8'hE8)) lut_n1634 (.I0(x774), .I1(x775), .I2(x776), .O(n1634));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1635 (.I0(x765), .I1(x766), .I2(x767), .I3(n1631), .I4(n1632), .O(n1635));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1636 (.I0(x771), .I1(x772), .I2(x773), .I3(n1634), .I4(n1635), .O(n1636));
  LUT3 #(.INIT(8'h96)) lut_n1637 (.I0(n1617), .I1(n1620), .I2(n1621), .O(n1637));
  LUT3 #(.INIT(8'hE8)) lut_n1638 (.I0(n1633), .I1(n1636), .I2(n1637), .O(n1638));
  LUT3 #(.INIT(8'hE8)) lut_n1639 (.I0(x780), .I1(x781), .I2(x782), .O(n1639));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1640 (.I0(x771), .I1(x772), .I2(x773), .I3(n1634), .I4(n1635), .O(n1640));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1641 (.I0(x777), .I1(x778), .I2(x779), .I3(n1639), .I4(n1640), .O(n1641));
  LUT3 #(.INIT(8'hE8)) lut_n1642 (.I0(x786), .I1(x787), .I2(x788), .O(n1642));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1643 (.I0(x777), .I1(x778), .I2(x779), .I3(n1639), .I4(n1640), .O(n1643));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1644 (.I0(x783), .I1(x784), .I2(x785), .I3(n1642), .I4(n1643), .O(n1644));
  LUT3 #(.INIT(8'h96)) lut_n1645 (.I0(n1633), .I1(n1636), .I2(n1637), .O(n1645));
  LUT3 #(.INIT(8'hE8)) lut_n1646 (.I0(n1641), .I1(n1644), .I2(n1645), .O(n1646));
  LUT3 #(.INIT(8'h96)) lut_n1647 (.I0(n1614), .I1(n1622), .I2(n1623), .O(n1647));
  LUT3 #(.INIT(8'hE8)) lut_n1648 (.I0(n1638), .I1(n1646), .I2(n1647), .O(n1648));
  LUT3 #(.INIT(8'hE8)) lut_n1649 (.I0(x792), .I1(x793), .I2(x794), .O(n1649));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1650 (.I0(x783), .I1(x784), .I2(x785), .I3(n1642), .I4(n1643), .O(n1650));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1651 (.I0(x789), .I1(x790), .I2(x791), .I3(n1649), .I4(n1650), .O(n1651));
  LUT3 #(.INIT(8'hE8)) lut_n1652 (.I0(x798), .I1(x799), .I2(x800), .O(n1652));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1653 (.I0(x789), .I1(x790), .I2(x791), .I3(n1649), .I4(n1650), .O(n1653));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1654 (.I0(x795), .I1(x796), .I2(x797), .I3(n1652), .I4(n1653), .O(n1654));
  LUT3 #(.INIT(8'h96)) lut_n1655 (.I0(n1641), .I1(n1644), .I2(n1645), .O(n1655));
  LUT3 #(.INIT(8'hE8)) lut_n1656 (.I0(n1651), .I1(n1654), .I2(n1655), .O(n1656));
  LUT3 #(.INIT(8'hE8)) lut_n1657 (.I0(x804), .I1(x805), .I2(x806), .O(n1657));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1658 (.I0(x795), .I1(x796), .I2(x797), .I3(n1652), .I4(n1653), .O(n1658));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1659 (.I0(x801), .I1(x802), .I2(x803), .I3(n1657), .I4(n1658), .O(n1659));
  LUT3 #(.INIT(8'hE8)) lut_n1660 (.I0(x810), .I1(x811), .I2(x812), .O(n1660));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1661 (.I0(x801), .I1(x802), .I2(x803), .I3(n1657), .I4(n1658), .O(n1661));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1662 (.I0(x807), .I1(x808), .I2(x809), .I3(n1660), .I4(n1661), .O(n1662));
  LUT3 #(.INIT(8'h96)) lut_n1663 (.I0(n1651), .I1(n1654), .I2(n1655), .O(n1663));
  LUT3 #(.INIT(8'hE8)) lut_n1664 (.I0(n1659), .I1(n1662), .I2(n1663), .O(n1664));
  LUT3 #(.INIT(8'h96)) lut_n1665 (.I0(n1638), .I1(n1646), .I2(n1647), .O(n1665));
  LUT3 #(.INIT(8'hE8)) lut_n1666 (.I0(n1656), .I1(n1664), .I2(n1665), .O(n1666));
  LUT3 #(.INIT(8'h96)) lut_n1667 (.I0(n1606), .I1(n1624), .I2(n1625), .O(n1667));
  LUT3 #(.INIT(8'hE8)) lut_n1668 (.I0(n1648), .I1(n1666), .I2(n1667), .O(n1668));
  LUT3 #(.INIT(8'hE8)) lut_n1669 (.I0(x816), .I1(x817), .I2(x818), .O(n1669));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1670 (.I0(x807), .I1(x808), .I2(x809), .I3(n1660), .I4(n1661), .O(n1670));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1671 (.I0(x813), .I1(x814), .I2(x815), .I3(n1669), .I4(n1670), .O(n1671));
  LUT3 #(.INIT(8'hE8)) lut_n1672 (.I0(x822), .I1(x823), .I2(x824), .O(n1672));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1673 (.I0(x813), .I1(x814), .I2(x815), .I3(n1669), .I4(n1670), .O(n1673));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1674 (.I0(x819), .I1(x820), .I2(x821), .I3(n1672), .I4(n1673), .O(n1674));
  LUT3 #(.INIT(8'h96)) lut_n1675 (.I0(n1659), .I1(n1662), .I2(n1663), .O(n1675));
  LUT3 #(.INIT(8'hE8)) lut_n1676 (.I0(n1671), .I1(n1674), .I2(n1675), .O(n1676));
  LUT3 #(.INIT(8'hE8)) lut_n1677 (.I0(x828), .I1(x829), .I2(x830), .O(n1677));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1678 (.I0(x819), .I1(x820), .I2(x821), .I3(n1672), .I4(n1673), .O(n1678));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1679 (.I0(x825), .I1(x826), .I2(x827), .I3(n1677), .I4(n1678), .O(n1679));
  LUT3 #(.INIT(8'hE8)) lut_n1680 (.I0(x834), .I1(x835), .I2(x836), .O(n1680));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1681 (.I0(x825), .I1(x826), .I2(x827), .I3(n1677), .I4(n1678), .O(n1681));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1682 (.I0(x831), .I1(x832), .I2(x833), .I3(n1680), .I4(n1681), .O(n1682));
  LUT3 #(.INIT(8'h96)) lut_n1683 (.I0(n1671), .I1(n1674), .I2(n1675), .O(n1683));
  LUT3 #(.INIT(8'hE8)) lut_n1684 (.I0(n1679), .I1(n1682), .I2(n1683), .O(n1684));
  LUT3 #(.INIT(8'h96)) lut_n1685 (.I0(n1656), .I1(n1664), .I2(n1665), .O(n1685));
  LUT3 #(.INIT(8'hE8)) lut_n1686 (.I0(n1676), .I1(n1684), .I2(n1685), .O(n1686));
  LUT3 #(.INIT(8'hE8)) lut_n1687 (.I0(x840), .I1(x841), .I2(x842), .O(n1687));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1688 (.I0(x831), .I1(x832), .I2(x833), .I3(n1680), .I4(n1681), .O(n1688));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1689 (.I0(x837), .I1(x838), .I2(x839), .I3(n1687), .I4(n1688), .O(n1689));
  LUT3 #(.INIT(8'hE8)) lut_n1690 (.I0(x846), .I1(x847), .I2(x848), .O(n1690));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1691 (.I0(x837), .I1(x838), .I2(x839), .I3(n1687), .I4(n1688), .O(n1691));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1692 (.I0(x843), .I1(x844), .I2(x845), .I3(n1690), .I4(n1691), .O(n1692));
  LUT3 #(.INIT(8'h96)) lut_n1693 (.I0(n1679), .I1(n1682), .I2(n1683), .O(n1693));
  LUT3 #(.INIT(8'hE8)) lut_n1694 (.I0(n1689), .I1(n1692), .I2(n1693), .O(n1694));
  LUT3 #(.INIT(8'hE8)) lut_n1695 (.I0(x852), .I1(x853), .I2(x854), .O(n1695));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1696 (.I0(x843), .I1(x844), .I2(x845), .I3(n1690), .I4(n1691), .O(n1696));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1697 (.I0(x849), .I1(x850), .I2(x851), .I3(n1695), .I4(n1696), .O(n1697));
  LUT3 #(.INIT(8'hE8)) lut_n1698 (.I0(x858), .I1(x859), .I2(x860), .O(n1698));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1699 (.I0(x849), .I1(x850), .I2(x851), .I3(n1695), .I4(n1696), .O(n1699));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1700 (.I0(x855), .I1(x856), .I2(x857), .I3(n1698), .I4(n1699), .O(n1700));
  LUT3 #(.INIT(8'h96)) lut_n1701 (.I0(n1689), .I1(n1692), .I2(n1693), .O(n1701));
  LUT3 #(.INIT(8'hE8)) lut_n1702 (.I0(n1697), .I1(n1700), .I2(n1701), .O(n1702));
  LUT3 #(.INIT(8'h96)) lut_n1703 (.I0(n1676), .I1(n1684), .I2(n1685), .O(n1703));
  LUT3 #(.INIT(8'hE8)) lut_n1704 (.I0(n1694), .I1(n1702), .I2(n1703), .O(n1704));
  LUT3 #(.INIT(8'h96)) lut_n1705 (.I0(n1648), .I1(n1666), .I2(n1667), .O(n1705));
  LUT3 #(.INIT(8'hE8)) lut_n1706 (.I0(n1686), .I1(n1704), .I2(n1705), .O(n1706));
  LUT3 #(.INIT(8'h96)) lut_n1707 (.I0(n1588), .I1(n1626), .I2(n1627), .O(n1707));
  LUT3 #(.INIT(8'hE8)) lut_n1708 (.I0(n1668), .I1(n1706), .I2(n1707), .O(n1708));
  LUT3 #(.INIT(8'hE8)) lut_n1709 (.I0(x864), .I1(x865), .I2(x866), .O(n1709));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1710 (.I0(x855), .I1(x856), .I2(x857), .I3(n1698), .I4(n1699), .O(n1710));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1711 (.I0(x861), .I1(x862), .I2(x863), .I3(n1709), .I4(n1710), .O(n1711));
  LUT3 #(.INIT(8'hE8)) lut_n1712 (.I0(x870), .I1(x871), .I2(x872), .O(n1712));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1713 (.I0(x861), .I1(x862), .I2(x863), .I3(n1709), .I4(n1710), .O(n1713));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1714 (.I0(x867), .I1(x868), .I2(x869), .I3(n1712), .I4(n1713), .O(n1714));
  LUT3 #(.INIT(8'h96)) lut_n1715 (.I0(n1697), .I1(n1700), .I2(n1701), .O(n1715));
  LUT3 #(.INIT(8'hE8)) lut_n1716 (.I0(n1711), .I1(n1714), .I2(n1715), .O(n1716));
  LUT3 #(.INIT(8'hE8)) lut_n1717 (.I0(x876), .I1(x877), .I2(x878), .O(n1717));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1718 (.I0(x867), .I1(x868), .I2(x869), .I3(n1712), .I4(n1713), .O(n1718));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1719 (.I0(x873), .I1(x874), .I2(x875), .I3(n1717), .I4(n1718), .O(n1719));
  LUT3 #(.INIT(8'hE8)) lut_n1720 (.I0(x882), .I1(x883), .I2(x884), .O(n1720));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1721 (.I0(x873), .I1(x874), .I2(x875), .I3(n1717), .I4(n1718), .O(n1721));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1722 (.I0(x879), .I1(x880), .I2(x881), .I3(n1720), .I4(n1721), .O(n1722));
  LUT3 #(.INIT(8'h96)) lut_n1723 (.I0(n1711), .I1(n1714), .I2(n1715), .O(n1723));
  LUT3 #(.INIT(8'hE8)) lut_n1724 (.I0(n1719), .I1(n1722), .I2(n1723), .O(n1724));
  LUT3 #(.INIT(8'h96)) lut_n1725 (.I0(n1694), .I1(n1702), .I2(n1703), .O(n1725));
  LUT3 #(.INIT(8'hE8)) lut_n1726 (.I0(n1716), .I1(n1724), .I2(n1725), .O(n1726));
  LUT3 #(.INIT(8'hE8)) lut_n1727 (.I0(x888), .I1(x889), .I2(x890), .O(n1727));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1728 (.I0(x879), .I1(x880), .I2(x881), .I3(n1720), .I4(n1721), .O(n1728));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1729 (.I0(x885), .I1(x886), .I2(x887), .I3(n1727), .I4(n1728), .O(n1729));
  LUT3 #(.INIT(8'hE8)) lut_n1730 (.I0(x894), .I1(x895), .I2(x896), .O(n1730));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1731 (.I0(x885), .I1(x886), .I2(x887), .I3(n1727), .I4(n1728), .O(n1731));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1732 (.I0(x891), .I1(x892), .I2(x893), .I3(n1730), .I4(n1731), .O(n1732));
  LUT3 #(.INIT(8'h96)) lut_n1733 (.I0(n1719), .I1(n1722), .I2(n1723), .O(n1733));
  LUT3 #(.INIT(8'hE8)) lut_n1734 (.I0(n1729), .I1(n1732), .I2(n1733), .O(n1734));
  LUT3 #(.INIT(8'hE8)) lut_n1735 (.I0(x900), .I1(x901), .I2(x902), .O(n1735));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1736 (.I0(x891), .I1(x892), .I2(x893), .I3(n1730), .I4(n1731), .O(n1736));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1737 (.I0(x897), .I1(x898), .I2(x899), .I3(n1735), .I4(n1736), .O(n1737));
  LUT3 #(.INIT(8'hE8)) lut_n1738 (.I0(x906), .I1(x907), .I2(x908), .O(n1738));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1739 (.I0(x897), .I1(x898), .I2(x899), .I3(n1735), .I4(n1736), .O(n1739));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1740 (.I0(x903), .I1(x904), .I2(x905), .I3(n1738), .I4(n1739), .O(n1740));
  LUT3 #(.INIT(8'h96)) lut_n1741 (.I0(n1729), .I1(n1732), .I2(n1733), .O(n1741));
  LUT3 #(.INIT(8'hE8)) lut_n1742 (.I0(n1737), .I1(n1740), .I2(n1741), .O(n1742));
  LUT3 #(.INIT(8'h96)) lut_n1743 (.I0(n1716), .I1(n1724), .I2(n1725), .O(n1743));
  LUT3 #(.INIT(8'hE8)) lut_n1744 (.I0(n1734), .I1(n1742), .I2(n1743), .O(n1744));
  LUT3 #(.INIT(8'h96)) lut_n1745 (.I0(n1686), .I1(n1704), .I2(n1705), .O(n1745));
  LUT3 #(.INIT(8'hE8)) lut_n1746 (.I0(n1726), .I1(n1744), .I2(n1745), .O(n1746));
  LUT3 #(.INIT(8'hE8)) lut_n1747 (.I0(x912), .I1(x913), .I2(x914), .O(n1747));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1748 (.I0(x903), .I1(x904), .I2(x905), .I3(n1738), .I4(n1739), .O(n1748));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1749 (.I0(x909), .I1(x910), .I2(x911), .I3(n1747), .I4(n1748), .O(n1749));
  LUT3 #(.INIT(8'hE8)) lut_n1750 (.I0(x918), .I1(x919), .I2(x920), .O(n1750));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1751 (.I0(x909), .I1(x910), .I2(x911), .I3(n1747), .I4(n1748), .O(n1751));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1752 (.I0(x915), .I1(x916), .I2(x917), .I3(n1750), .I4(n1751), .O(n1752));
  LUT3 #(.INIT(8'h96)) lut_n1753 (.I0(n1737), .I1(n1740), .I2(n1741), .O(n1753));
  LUT3 #(.INIT(8'hE8)) lut_n1754 (.I0(n1749), .I1(n1752), .I2(n1753), .O(n1754));
  LUT3 #(.INIT(8'hE8)) lut_n1755 (.I0(x924), .I1(x925), .I2(x926), .O(n1755));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1756 (.I0(x915), .I1(x916), .I2(x917), .I3(n1750), .I4(n1751), .O(n1756));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1757 (.I0(x921), .I1(x922), .I2(x923), .I3(n1755), .I4(n1756), .O(n1757));
  LUT3 #(.INIT(8'hE8)) lut_n1758 (.I0(x930), .I1(x931), .I2(x932), .O(n1758));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1759 (.I0(x921), .I1(x922), .I2(x923), .I3(n1755), .I4(n1756), .O(n1759));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1760 (.I0(x927), .I1(x928), .I2(x929), .I3(n1758), .I4(n1759), .O(n1760));
  LUT3 #(.INIT(8'h96)) lut_n1761 (.I0(n1749), .I1(n1752), .I2(n1753), .O(n1761));
  LUT3 #(.INIT(8'hE8)) lut_n1762 (.I0(n1757), .I1(n1760), .I2(n1761), .O(n1762));
  LUT3 #(.INIT(8'h96)) lut_n1763 (.I0(n1734), .I1(n1742), .I2(n1743), .O(n1763));
  LUT3 #(.INIT(8'hE8)) lut_n1764 (.I0(n1754), .I1(n1762), .I2(n1763), .O(n1764));
  LUT3 #(.INIT(8'hE8)) lut_n1765 (.I0(x936), .I1(x937), .I2(x938), .O(n1765));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1766 (.I0(x927), .I1(x928), .I2(x929), .I3(n1758), .I4(n1759), .O(n1766));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1767 (.I0(x933), .I1(x934), .I2(x935), .I3(n1765), .I4(n1766), .O(n1767));
  LUT3 #(.INIT(8'hE8)) lut_n1768 (.I0(x942), .I1(x943), .I2(x944), .O(n1768));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1769 (.I0(x933), .I1(x934), .I2(x935), .I3(n1765), .I4(n1766), .O(n1769));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1770 (.I0(x939), .I1(x940), .I2(x941), .I3(n1768), .I4(n1769), .O(n1770));
  LUT3 #(.INIT(8'h96)) lut_n1771 (.I0(n1757), .I1(n1760), .I2(n1761), .O(n1771));
  LUT3 #(.INIT(8'hE8)) lut_n1772 (.I0(n1767), .I1(n1770), .I2(n1771), .O(n1772));
  LUT3 #(.INIT(8'hE8)) lut_n1773 (.I0(x948), .I1(x949), .I2(x950), .O(n1773));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1774 (.I0(x939), .I1(x940), .I2(x941), .I3(n1768), .I4(n1769), .O(n1774));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1775 (.I0(x945), .I1(x946), .I2(x947), .I3(n1773), .I4(n1774), .O(n1775));
  LUT3 #(.INIT(8'hE8)) lut_n1776 (.I0(x954), .I1(x955), .I2(x956), .O(n1776));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1777 (.I0(x945), .I1(x946), .I2(x947), .I3(n1773), .I4(n1774), .O(n1777));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1778 (.I0(x951), .I1(x952), .I2(x953), .I3(n1776), .I4(n1777), .O(n1778));
  LUT3 #(.INIT(8'h96)) lut_n1779 (.I0(n1767), .I1(n1770), .I2(n1771), .O(n1779));
  LUT3 #(.INIT(8'hE8)) lut_n1780 (.I0(n1775), .I1(n1778), .I2(n1779), .O(n1780));
  LUT3 #(.INIT(8'h96)) lut_n1781 (.I0(n1754), .I1(n1762), .I2(n1763), .O(n1781));
  LUT3 #(.INIT(8'hE8)) lut_n1782 (.I0(n1772), .I1(n1780), .I2(n1781), .O(n1782));
  LUT3 #(.INIT(8'h96)) lut_n1783 (.I0(n1726), .I1(n1744), .I2(n1745), .O(n1783));
  LUT3 #(.INIT(8'hE8)) lut_n1784 (.I0(n1764), .I1(n1782), .I2(n1783), .O(n1784));
  LUT3 #(.INIT(8'h96)) lut_n1785 (.I0(n1668), .I1(n1706), .I2(n1707), .O(n1785));
  LUT3 #(.INIT(8'hE8)) lut_n1786 (.I0(n1746), .I1(n1784), .I2(n1785), .O(n1786));
  LUT3 #(.INIT(8'h96)) lut_n1787 (.I0(n1550), .I1(n1628), .I2(n1629), .O(n1787));
  LUT3 #(.INIT(8'hE8)) lut_n1788 (.I0(n1708), .I1(n1786), .I2(n1787), .O(n1788));
  LUT3 #(.INIT(8'hE8)) lut_n1789 (.I0(x960), .I1(x961), .I2(x962), .O(n1789));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1790 (.I0(x951), .I1(x952), .I2(x953), .I3(n1776), .I4(n1777), .O(n1790));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1791 (.I0(x957), .I1(x958), .I2(x959), .I3(n1789), .I4(n1790), .O(n1791));
  LUT3 #(.INIT(8'hE8)) lut_n1792 (.I0(x966), .I1(x967), .I2(x968), .O(n1792));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1793 (.I0(x957), .I1(x958), .I2(x959), .I3(n1789), .I4(n1790), .O(n1793));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1794 (.I0(x963), .I1(x964), .I2(x965), .I3(n1792), .I4(n1793), .O(n1794));
  LUT3 #(.INIT(8'h96)) lut_n1795 (.I0(n1775), .I1(n1778), .I2(n1779), .O(n1795));
  LUT3 #(.INIT(8'hE8)) lut_n1796 (.I0(n1791), .I1(n1794), .I2(n1795), .O(n1796));
  LUT3 #(.INIT(8'hE8)) lut_n1797 (.I0(x972), .I1(x973), .I2(x974), .O(n1797));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1798 (.I0(x963), .I1(x964), .I2(x965), .I3(n1792), .I4(n1793), .O(n1798));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1799 (.I0(x969), .I1(x970), .I2(x971), .I3(n1797), .I4(n1798), .O(n1799));
  LUT3 #(.INIT(8'hE8)) lut_n1800 (.I0(x978), .I1(x979), .I2(x980), .O(n1800));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1801 (.I0(x969), .I1(x970), .I2(x971), .I3(n1797), .I4(n1798), .O(n1801));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1802 (.I0(x975), .I1(x976), .I2(x977), .I3(n1800), .I4(n1801), .O(n1802));
  LUT3 #(.INIT(8'h96)) lut_n1803 (.I0(n1791), .I1(n1794), .I2(n1795), .O(n1803));
  LUT3 #(.INIT(8'hE8)) lut_n1804 (.I0(n1799), .I1(n1802), .I2(n1803), .O(n1804));
  LUT3 #(.INIT(8'h96)) lut_n1805 (.I0(n1772), .I1(n1780), .I2(n1781), .O(n1805));
  LUT3 #(.INIT(8'hE8)) lut_n1806 (.I0(n1796), .I1(n1804), .I2(n1805), .O(n1806));
  LUT3 #(.INIT(8'hE8)) lut_n1807 (.I0(x984), .I1(x985), .I2(x986), .O(n1807));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1808 (.I0(x975), .I1(x976), .I2(x977), .I3(n1800), .I4(n1801), .O(n1808));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1809 (.I0(x981), .I1(x982), .I2(x983), .I3(n1807), .I4(n1808), .O(n1809));
  LUT3 #(.INIT(8'hE8)) lut_n1810 (.I0(x990), .I1(x991), .I2(x992), .O(n1810));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1811 (.I0(x981), .I1(x982), .I2(x983), .I3(n1807), .I4(n1808), .O(n1811));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1812 (.I0(x987), .I1(x988), .I2(x989), .I3(n1810), .I4(n1811), .O(n1812));
  LUT3 #(.INIT(8'h96)) lut_n1813 (.I0(n1799), .I1(n1802), .I2(n1803), .O(n1813));
  LUT3 #(.INIT(8'hE8)) lut_n1814 (.I0(n1809), .I1(n1812), .I2(n1813), .O(n1814));
  LUT3 #(.INIT(8'hE8)) lut_n1815 (.I0(x996), .I1(x997), .I2(x998), .O(n1815));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1816 (.I0(x987), .I1(x988), .I2(x989), .I3(n1810), .I4(n1811), .O(n1816));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1817 (.I0(x993), .I1(x994), .I2(x995), .I3(n1815), .I4(n1816), .O(n1817));
  LUT3 #(.INIT(8'hE8)) lut_n1818 (.I0(x1002), .I1(x1003), .I2(x1004), .O(n1818));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1819 (.I0(x993), .I1(x994), .I2(x995), .I3(n1815), .I4(n1816), .O(n1819));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1820 (.I0(x999), .I1(x1000), .I2(x1001), .I3(n1818), .I4(n1819), .O(n1820));
  LUT3 #(.INIT(8'h96)) lut_n1821 (.I0(n1809), .I1(n1812), .I2(n1813), .O(n1821));
  LUT3 #(.INIT(8'hE8)) lut_n1822 (.I0(n1817), .I1(n1820), .I2(n1821), .O(n1822));
  LUT3 #(.INIT(8'h96)) lut_n1823 (.I0(n1796), .I1(n1804), .I2(n1805), .O(n1823));
  LUT3 #(.INIT(8'hE8)) lut_n1824 (.I0(n1814), .I1(n1822), .I2(n1823), .O(n1824));
  LUT3 #(.INIT(8'h96)) lut_n1825 (.I0(n1764), .I1(n1782), .I2(n1783), .O(n1825));
  LUT3 #(.INIT(8'hE8)) lut_n1826 (.I0(n1806), .I1(n1824), .I2(n1825), .O(n1826));
  LUT3 #(.INIT(8'hE8)) lut_n1827 (.I0(x1008), .I1(x1009), .I2(x1010), .O(n1827));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1828 (.I0(x999), .I1(x1000), .I2(x1001), .I3(n1818), .I4(n1819), .O(n1828));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n1829 (.I0(x1005), .I1(x1006), .I2(x1007), .I3(n1827), .I4(n1828), .O(n1829));
  LUT5 #(.INIT(32'hE81717E8)) lut_n1830 (.I0(x1005), .I1(x1006), .I2(x1007), .I3(n1827), .I4(n1828), .O(n1830));
  LUT4 #(.INIT(16'hFFE8)) lut_n1831 (.I0(x1011), .I1(x1012), .I2(x1013), .I3(n1830), .O(n1831));
  LUT3 #(.INIT(8'h96)) lut_n1832 (.I0(n1817), .I1(n1820), .I2(n1821), .O(n1832));
  LUT3 #(.INIT(8'hE8)) lut_n1833 (.I0(n1829), .I1(n1831), .I2(n1832), .O(n1833));
  LUT4 #(.INIT(16'h17E8)) lut_n1834 (.I0(x1011), .I1(x1012), .I2(x1013), .I3(n1830), .O(n1834));
  LUT3 #(.INIT(8'h96)) lut_n1835 (.I0(x0), .I1(x1), .I2(x2), .O(n1835));
  LUT3 #(.INIT(8'h96)) lut_n1836 (.I0(x6), .I1(x7), .I2(x8), .O(n1836));
  LUT5 #(.INIT(32'hFF969600)) lut_n1837 (.I0(x3), .I1(x4), .I2(x5), .I3(n1835), .I4(n1836), .O(n1837));
  LUT3 #(.INIT(8'h96)) lut_n1838 (.I0(x12), .I1(x13), .I2(x14), .O(n1838));
  LUT5 #(.INIT(32'h96696996)) lut_n1839 (.I0(x3), .I1(x4), .I2(x5), .I3(n1835), .I4(n1836), .O(n1839));
  LUT5 #(.INIT(32'hFF969600)) lut_n1840 (.I0(x9), .I1(x10), .I2(x11), .I3(n1838), .I4(n1839), .O(n1840));
  LUT3 #(.INIT(8'hE8)) lut_n1841 (.I0(n1834), .I1(n1837), .I2(n1840), .O(n1841));
  LUT3 #(.INIT(8'h96)) lut_n1842 (.I0(n1829), .I1(n1831), .I2(n1832), .O(n1842));
  LUT3 #(.INIT(8'hD4)) lut_n1843 (.I0(n1834), .I1(n1841), .I2(n1842), .O(n1843));
  LUT3 #(.INIT(8'h96)) lut_n1844 (.I0(n1814), .I1(n1822), .I2(n1823), .O(n1844));
  LUT3 #(.INIT(8'hE8)) lut_n1845 (.I0(n1833), .I1(n1843), .I2(n1844), .O(n1845));
  LUT3 #(.INIT(8'h96)) lut_n1846 (.I0(x18), .I1(x19), .I2(x20), .O(n1846));
  LUT5 #(.INIT(32'h96696996)) lut_n1847 (.I0(x9), .I1(x10), .I2(x11), .I3(n1838), .I4(n1839), .O(n1847));
  LUT5 #(.INIT(32'hFF969600)) lut_n1848 (.I0(x15), .I1(x16), .I2(x17), .I3(n1846), .I4(n1847), .O(n1848));
  LUT3 #(.INIT(8'h96)) lut_n1849 (.I0(x24), .I1(x25), .I2(x26), .O(n1849));
  LUT5 #(.INIT(32'h96696996)) lut_n1850 (.I0(x15), .I1(x16), .I2(x17), .I3(n1846), .I4(n1847), .O(n1850));
  LUT5 #(.INIT(32'hFF969600)) lut_n1851 (.I0(x21), .I1(x22), .I2(x23), .I3(n1849), .I4(n1850), .O(n1851));
  LUT3 #(.INIT(8'h96)) lut_n1852 (.I0(n1834), .I1(n1837), .I2(n1840), .O(n1852));
  LUT3 #(.INIT(8'hE8)) lut_n1853 (.I0(n1848), .I1(n1851), .I2(n1852), .O(n1853));
  LUT3 #(.INIT(8'h96)) lut_n1854 (.I0(x27), .I1(x28), .I2(x29), .O(n1854));
  LUT5 #(.INIT(32'h96696996)) lut_n1855 (.I0(x21), .I1(x22), .I2(x23), .I3(n1849), .I4(n1850), .O(n1855));
  LUT5 #(.INIT(32'hFF969600)) lut_n1856 (.I0(x30), .I1(x31), .I2(x32), .I3(n1854), .I4(n1855), .O(n1856));
  LUT3 #(.INIT(8'h96)) lut_n1857 (.I0(x36), .I1(x37), .I2(x38), .O(n1857));
  LUT5 #(.INIT(32'h96696996)) lut_n1858 (.I0(x30), .I1(x31), .I2(x32), .I3(n1854), .I4(n1855), .O(n1858));
  LUT5 #(.INIT(32'hFF969600)) lut_n1859 (.I0(x33), .I1(x34), .I2(x35), .I3(n1857), .I4(n1858), .O(n1859));
  LUT3 #(.INIT(8'h96)) lut_n1860 (.I0(n1848), .I1(n1851), .I2(n1852), .O(n1860));
  LUT3 #(.INIT(8'hE8)) lut_n1861 (.I0(n1856), .I1(n1859), .I2(n1860), .O(n1861));
  LUT3 #(.INIT(8'h96)) lut_n1862 (.I0(n1834), .I1(n1841), .I2(n1842), .O(n1862));
  LUT3 #(.INIT(8'h8E)) lut_n1863 (.I0(n1853), .I1(n1861), .I2(n1862), .O(n1863));
  LUT3 #(.INIT(8'h96)) lut_n1864 (.I0(x42), .I1(x43), .I2(x44), .O(n1864));
  LUT5 #(.INIT(32'h96696996)) lut_n1865 (.I0(x33), .I1(x34), .I2(x35), .I3(n1857), .I4(n1858), .O(n1865));
  LUT5 #(.INIT(32'hFF969600)) lut_n1866 (.I0(x39), .I1(x40), .I2(x41), .I3(n1864), .I4(n1865), .O(n1866));
  LUT3 #(.INIT(8'h96)) lut_n1867 (.I0(x48), .I1(x49), .I2(x50), .O(n1867));
  LUT5 #(.INIT(32'h96696996)) lut_n1868 (.I0(x39), .I1(x40), .I2(x41), .I3(n1864), .I4(n1865), .O(n1868));
  LUT5 #(.INIT(32'hFF969600)) lut_n1869 (.I0(x45), .I1(x46), .I2(x47), .I3(n1867), .I4(n1868), .O(n1869));
  LUT3 #(.INIT(8'h96)) lut_n1870 (.I0(n1856), .I1(n1859), .I2(n1860), .O(n1870));
  LUT3 #(.INIT(8'hE8)) lut_n1871 (.I0(n1866), .I1(n1869), .I2(n1870), .O(n1871));
  LUT3 #(.INIT(8'h96)) lut_n1872 (.I0(x54), .I1(x55), .I2(x56), .O(n1872));
  LUT5 #(.INIT(32'h96696996)) lut_n1873 (.I0(x45), .I1(x46), .I2(x47), .I3(n1867), .I4(n1868), .O(n1873));
  LUT5 #(.INIT(32'hFF969600)) lut_n1874 (.I0(x51), .I1(x52), .I2(x53), .I3(n1872), .I4(n1873), .O(n1874));
  LUT3 #(.INIT(8'h96)) lut_n1875 (.I0(x60), .I1(x61), .I2(x62), .O(n1875));
  LUT5 #(.INIT(32'h96696996)) lut_n1876 (.I0(x51), .I1(x52), .I2(x53), .I3(n1872), .I4(n1873), .O(n1876));
  LUT5 #(.INIT(32'hFF969600)) lut_n1877 (.I0(x57), .I1(x58), .I2(x59), .I3(n1875), .I4(n1876), .O(n1877));
  LUT3 #(.INIT(8'h96)) lut_n1878 (.I0(n1866), .I1(n1869), .I2(n1870), .O(n1878));
  LUT3 #(.INIT(8'hE8)) lut_n1879 (.I0(n1874), .I1(n1877), .I2(n1878), .O(n1879));
  LUT3 #(.INIT(8'h96)) lut_n1880 (.I0(n1853), .I1(n1861), .I2(n1862), .O(n1880));
  LUT3 #(.INIT(8'h8E)) lut_n1881 (.I0(n1871), .I1(n1879), .I2(n1880), .O(n1881));
  LUT3 #(.INIT(8'h96)) lut_n1882 (.I0(n1833), .I1(n1843), .I2(n1844), .O(n1882));
  LUT3 #(.INIT(8'hE8)) lut_n1883 (.I0(n1863), .I1(n1881), .I2(n1882), .O(n1883));
  LUT3 #(.INIT(8'h96)) lut_n1884 (.I0(n1806), .I1(n1824), .I2(n1825), .O(n1884));
  LUT3 #(.INIT(8'hE8)) lut_n1885 (.I0(n1845), .I1(n1883), .I2(n1884), .O(n1885));
  LUT3 #(.INIT(8'h96)) lut_n1886 (.I0(n1746), .I1(n1784), .I2(n1785), .O(n1886));
  LUT3 #(.INIT(8'hE8)) lut_n1887 (.I0(n1826), .I1(n1885), .I2(n1886), .O(n1887));
  LUT3 #(.INIT(8'h96)) lut_n1888 (.I0(x66), .I1(x67), .I2(x68), .O(n1888));
  LUT5 #(.INIT(32'h96696996)) lut_n1889 (.I0(x57), .I1(x58), .I2(x59), .I3(n1875), .I4(n1876), .O(n1889));
  LUT5 #(.INIT(32'hFF969600)) lut_n1890 (.I0(x63), .I1(x64), .I2(x65), .I3(n1888), .I4(n1889), .O(n1890));
  LUT3 #(.INIT(8'h96)) lut_n1891 (.I0(x72), .I1(x73), .I2(x74), .O(n1891));
  LUT5 #(.INIT(32'h96696996)) lut_n1892 (.I0(x63), .I1(x64), .I2(x65), .I3(n1888), .I4(n1889), .O(n1892));
  LUT5 #(.INIT(32'hFF969600)) lut_n1893 (.I0(x69), .I1(x70), .I2(x71), .I3(n1891), .I4(n1892), .O(n1893));
  LUT3 #(.INIT(8'h96)) lut_n1894 (.I0(n1874), .I1(n1877), .I2(n1878), .O(n1894));
  LUT3 #(.INIT(8'hE8)) lut_n1895 (.I0(n1890), .I1(n1893), .I2(n1894), .O(n1895));
  LUT3 #(.INIT(8'h96)) lut_n1896 (.I0(x78), .I1(x79), .I2(x80), .O(n1896));
  LUT5 #(.INIT(32'h96696996)) lut_n1897 (.I0(x69), .I1(x70), .I2(x71), .I3(n1891), .I4(n1892), .O(n1897));
  LUT5 #(.INIT(32'hFF969600)) lut_n1898 (.I0(x75), .I1(x76), .I2(x77), .I3(n1896), .I4(n1897), .O(n1898));
  LUT3 #(.INIT(8'h96)) lut_n1899 (.I0(x84), .I1(x85), .I2(x86), .O(n1899));
  LUT5 #(.INIT(32'h96696996)) lut_n1900 (.I0(x75), .I1(x76), .I2(x77), .I3(n1896), .I4(n1897), .O(n1900));
  LUT5 #(.INIT(32'hFF969600)) lut_n1901 (.I0(x81), .I1(x82), .I2(x83), .I3(n1899), .I4(n1900), .O(n1901));
  LUT3 #(.INIT(8'h96)) lut_n1902 (.I0(n1890), .I1(n1893), .I2(n1894), .O(n1902));
  LUT3 #(.INIT(8'hE8)) lut_n1903 (.I0(n1898), .I1(n1901), .I2(n1902), .O(n1903));
  LUT3 #(.INIT(8'h96)) lut_n1904 (.I0(n1871), .I1(n1879), .I2(n1880), .O(n1904));
  LUT3 #(.INIT(8'h8E)) lut_n1905 (.I0(n1895), .I1(n1903), .I2(n1904), .O(n1905));
  LUT3 #(.INIT(8'h96)) lut_n1906 (.I0(x90), .I1(x91), .I2(x92), .O(n1906));
  LUT5 #(.INIT(32'h96696996)) lut_n1907 (.I0(x81), .I1(x82), .I2(x83), .I3(n1899), .I4(n1900), .O(n1907));
  LUT5 #(.INIT(32'hFF969600)) lut_n1908 (.I0(x87), .I1(x88), .I2(x89), .I3(n1906), .I4(n1907), .O(n1908));
  LUT3 #(.INIT(8'h96)) lut_n1909 (.I0(x96), .I1(x97), .I2(x98), .O(n1909));
  LUT5 #(.INIT(32'h96696996)) lut_n1910 (.I0(x87), .I1(x88), .I2(x89), .I3(n1906), .I4(n1907), .O(n1910));
  LUT5 #(.INIT(32'hFF969600)) lut_n1911 (.I0(x93), .I1(x94), .I2(x95), .I3(n1909), .I4(n1910), .O(n1911));
  LUT3 #(.INIT(8'h96)) lut_n1912 (.I0(n1898), .I1(n1901), .I2(n1902), .O(n1912));
  LUT3 #(.INIT(8'hE8)) lut_n1913 (.I0(n1908), .I1(n1911), .I2(n1912), .O(n1913));
  LUT3 #(.INIT(8'h96)) lut_n1914 (.I0(x102), .I1(x103), .I2(x104), .O(n1914));
  LUT5 #(.INIT(32'h96696996)) lut_n1915 (.I0(x93), .I1(x94), .I2(x95), .I3(n1909), .I4(n1910), .O(n1915));
  LUT5 #(.INIT(32'hFF969600)) lut_n1916 (.I0(x99), .I1(x100), .I2(x101), .I3(n1914), .I4(n1915), .O(n1916));
  LUT3 #(.INIT(8'h96)) lut_n1917 (.I0(x108), .I1(x109), .I2(x110), .O(n1917));
  LUT5 #(.INIT(32'h96696996)) lut_n1918 (.I0(x99), .I1(x100), .I2(x101), .I3(n1914), .I4(n1915), .O(n1918));
  LUT5 #(.INIT(32'hFF969600)) lut_n1919 (.I0(x105), .I1(x106), .I2(x107), .I3(n1917), .I4(n1918), .O(n1919));
  LUT3 #(.INIT(8'h96)) lut_n1920 (.I0(n1908), .I1(n1911), .I2(n1912), .O(n1920));
  LUT3 #(.INIT(8'hE8)) lut_n1921 (.I0(n1916), .I1(n1919), .I2(n1920), .O(n1921));
  LUT3 #(.INIT(8'h96)) lut_n1922 (.I0(n1895), .I1(n1903), .I2(n1904), .O(n1922));
  LUT3 #(.INIT(8'h8E)) lut_n1923 (.I0(n1913), .I1(n1921), .I2(n1922), .O(n1923));
  LUT3 #(.INIT(8'h96)) lut_n1924 (.I0(n1863), .I1(n1881), .I2(n1882), .O(n1924));
  LUT3 #(.INIT(8'hE8)) lut_n1925 (.I0(n1905), .I1(n1923), .I2(n1924), .O(n1925));
  LUT3 #(.INIT(8'h96)) lut_n1926 (.I0(x114), .I1(x115), .I2(x116), .O(n1926));
  LUT5 #(.INIT(32'h96696996)) lut_n1927 (.I0(x105), .I1(x106), .I2(x107), .I3(n1917), .I4(n1918), .O(n1927));
  LUT5 #(.INIT(32'hFF969600)) lut_n1928 (.I0(x111), .I1(x112), .I2(x113), .I3(n1926), .I4(n1927), .O(n1928));
  LUT3 #(.INIT(8'h96)) lut_n1929 (.I0(x120), .I1(x121), .I2(x122), .O(n1929));
  LUT5 #(.INIT(32'h96696996)) lut_n1930 (.I0(x111), .I1(x112), .I2(x113), .I3(n1926), .I4(n1927), .O(n1930));
  LUT5 #(.INIT(32'hFF969600)) lut_n1931 (.I0(x117), .I1(x118), .I2(x119), .I3(n1929), .I4(n1930), .O(n1931));
  LUT3 #(.INIT(8'h96)) lut_n1932 (.I0(n1916), .I1(n1919), .I2(n1920), .O(n1932));
  LUT3 #(.INIT(8'hE8)) lut_n1933 (.I0(n1928), .I1(n1931), .I2(n1932), .O(n1933));
  LUT3 #(.INIT(8'h96)) lut_n1934 (.I0(x126), .I1(x127), .I2(x128), .O(n1934));
  LUT5 #(.INIT(32'h96696996)) lut_n1935 (.I0(x117), .I1(x118), .I2(x119), .I3(n1929), .I4(n1930), .O(n1935));
  LUT5 #(.INIT(32'hFF969600)) lut_n1936 (.I0(x123), .I1(x124), .I2(x125), .I3(n1934), .I4(n1935), .O(n1936));
  LUT3 #(.INIT(8'h96)) lut_n1937 (.I0(x132), .I1(x133), .I2(x134), .O(n1937));
  LUT5 #(.INIT(32'h96696996)) lut_n1938 (.I0(x123), .I1(x124), .I2(x125), .I3(n1934), .I4(n1935), .O(n1938));
  LUT5 #(.INIT(32'hFF969600)) lut_n1939 (.I0(x129), .I1(x130), .I2(x131), .I3(n1937), .I4(n1938), .O(n1939));
  LUT3 #(.INIT(8'h96)) lut_n1940 (.I0(n1928), .I1(n1931), .I2(n1932), .O(n1940));
  LUT3 #(.INIT(8'hE8)) lut_n1941 (.I0(n1936), .I1(n1939), .I2(n1940), .O(n1941));
  LUT3 #(.INIT(8'h96)) lut_n1942 (.I0(n1913), .I1(n1921), .I2(n1922), .O(n1942));
  LUT3 #(.INIT(8'h8E)) lut_n1943 (.I0(n1933), .I1(n1941), .I2(n1942), .O(n1943));
  LUT3 #(.INIT(8'h96)) lut_n1944 (.I0(x138), .I1(x139), .I2(x140), .O(n1944));
  LUT5 #(.INIT(32'h96696996)) lut_n1945 (.I0(x129), .I1(x130), .I2(x131), .I3(n1937), .I4(n1938), .O(n1945));
  LUT5 #(.INIT(32'hFF969600)) lut_n1946 (.I0(x135), .I1(x136), .I2(x137), .I3(n1944), .I4(n1945), .O(n1946));
  LUT3 #(.INIT(8'h96)) lut_n1947 (.I0(x144), .I1(x145), .I2(x146), .O(n1947));
  LUT5 #(.INIT(32'h96696996)) lut_n1948 (.I0(x135), .I1(x136), .I2(x137), .I3(n1944), .I4(n1945), .O(n1948));
  LUT5 #(.INIT(32'hFF969600)) lut_n1949 (.I0(x141), .I1(x142), .I2(x143), .I3(n1947), .I4(n1948), .O(n1949));
  LUT3 #(.INIT(8'h96)) lut_n1950 (.I0(n1936), .I1(n1939), .I2(n1940), .O(n1950));
  LUT3 #(.INIT(8'hE8)) lut_n1951 (.I0(n1946), .I1(n1949), .I2(n1950), .O(n1951));
  LUT3 #(.INIT(8'h96)) lut_n1952 (.I0(x150), .I1(x151), .I2(x152), .O(n1952));
  LUT5 #(.INIT(32'h96696996)) lut_n1953 (.I0(x141), .I1(x142), .I2(x143), .I3(n1947), .I4(n1948), .O(n1953));
  LUT5 #(.INIT(32'hFF969600)) lut_n1954 (.I0(x147), .I1(x148), .I2(x149), .I3(n1952), .I4(n1953), .O(n1954));
  LUT3 #(.INIT(8'h96)) lut_n1955 (.I0(x156), .I1(x157), .I2(x158), .O(n1955));
  LUT5 #(.INIT(32'h96696996)) lut_n1956 (.I0(x147), .I1(x148), .I2(x149), .I3(n1952), .I4(n1953), .O(n1956));
  LUT5 #(.INIT(32'hFF969600)) lut_n1957 (.I0(x153), .I1(x154), .I2(x155), .I3(n1955), .I4(n1956), .O(n1957));
  LUT3 #(.INIT(8'h96)) lut_n1958 (.I0(n1946), .I1(n1949), .I2(n1950), .O(n1958));
  LUT3 #(.INIT(8'hE8)) lut_n1959 (.I0(n1954), .I1(n1957), .I2(n1958), .O(n1959));
  LUT3 #(.INIT(8'h96)) lut_n1960 (.I0(n1933), .I1(n1941), .I2(n1942), .O(n1960));
  LUT3 #(.INIT(8'h8E)) lut_n1961 (.I0(n1951), .I1(n1959), .I2(n1960), .O(n1961));
  LUT3 #(.INIT(8'h96)) lut_n1962 (.I0(n1905), .I1(n1923), .I2(n1924), .O(n1962));
  LUT3 #(.INIT(8'hE8)) lut_n1963 (.I0(n1943), .I1(n1961), .I2(n1962), .O(n1963));
  LUT3 #(.INIT(8'h96)) lut_n1964 (.I0(n1845), .I1(n1883), .I2(n1884), .O(n1964));
  LUT3 #(.INIT(8'hE8)) lut_n1965 (.I0(n1925), .I1(n1963), .I2(n1964), .O(n1965));
  LUT3 #(.INIT(8'h96)) lut_n1966 (.I0(x162), .I1(x163), .I2(x164), .O(n1966));
  LUT5 #(.INIT(32'h96696996)) lut_n1967 (.I0(x153), .I1(x154), .I2(x155), .I3(n1955), .I4(n1956), .O(n1967));
  LUT5 #(.INIT(32'hFF969600)) lut_n1968 (.I0(x159), .I1(x160), .I2(x161), .I3(n1966), .I4(n1967), .O(n1968));
  LUT3 #(.INIT(8'h96)) lut_n1969 (.I0(x168), .I1(x169), .I2(x170), .O(n1969));
  LUT5 #(.INIT(32'h96696996)) lut_n1970 (.I0(x159), .I1(x160), .I2(x161), .I3(n1966), .I4(n1967), .O(n1970));
  LUT5 #(.INIT(32'hFF969600)) lut_n1971 (.I0(x165), .I1(x166), .I2(x167), .I3(n1969), .I4(n1970), .O(n1971));
  LUT3 #(.INIT(8'h96)) lut_n1972 (.I0(n1954), .I1(n1957), .I2(n1958), .O(n1972));
  LUT3 #(.INIT(8'hE8)) lut_n1973 (.I0(n1968), .I1(n1971), .I2(n1972), .O(n1973));
  LUT3 #(.INIT(8'h96)) lut_n1974 (.I0(x174), .I1(x175), .I2(x176), .O(n1974));
  LUT5 #(.INIT(32'h96696996)) lut_n1975 (.I0(x165), .I1(x166), .I2(x167), .I3(n1969), .I4(n1970), .O(n1975));
  LUT5 #(.INIT(32'hFF969600)) lut_n1976 (.I0(x171), .I1(x172), .I2(x173), .I3(n1974), .I4(n1975), .O(n1976));
  LUT3 #(.INIT(8'h96)) lut_n1977 (.I0(x180), .I1(x181), .I2(x182), .O(n1977));
  LUT5 #(.INIT(32'h96696996)) lut_n1978 (.I0(x171), .I1(x172), .I2(x173), .I3(n1974), .I4(n1975), .O(n1978));
  LUT5 #(.INIT(32'hFF969600)) lut_n1979 (.I0(x177), .I1(x178), .I2(x179), .I3(n1977), .I4(n1978), .O(n1979));
  LUT3 #(.INIT(8'h96)) lut_n1980 (.I0(n1968), .I1(n1971), .I2(n1972), .O(n1980));
  LUT3 #(.INIT(8'hE8)) lut_n1981 (.I0(n1976), .I1(n1979), .I2(n1980), .O(n1981));
  LUT3 #(.INIT(8'h96)) lut_n1982 (.I0(n1951), .I1(n1959), .I2(n1960), .O(n1982));
  LUT3 #(.INIT(8'h8E)) lut_n1983 (.I0(n1973), .I1(n1981), .I2(n1982), .O(n1983));
  LUT3 #(.INIT(8'h96)) lut_n1984 (.I0(x186), .I1(x187), .I2(x188), .O(n1984));
  LUT5 #(.INIT(32'h96696996)) lut_n1985 (.I0(x177), .I1(x178), .I2(x179), .I3(n1977), .I4(n1978), .O(n1985));
  LUT5 #(.INIT(32'hFF969600)) lut_n1986 (.I0(x183), .I1(x184), .I2(x185), .I3(n1984), .I4(n1985), .O(n1986));
  LUT3 #(.INIT(8'h96)) lut_n1987 (.I0(x192), .I1(x193), .I2(x194), .O(n1987));
  LUT5 #(.INIT(32'h96696996)) lut_n1988 (.I0(x183), .I1(x184), .I2(x185), .I3(n1984), .I4(n1985), .O(n1988));
  LUT5 #(.INIT(32'hFF969600)) lut_n1989 (.I0(x189), .I1(x190), .I2(x191), .I3(n1987), .I4(n1988), .O(n1989));
  LUT3 #(.INIT(8'h96)) lut_n1990 (.I0(n1976), .I1(n1979), .I2(n1980), .O(n1990));
  LUT3 #(.INIT(8'hE8)) lut_n1991 (.I0(n1986), .I1(n1989), .I2(n1990), .O(n1991));
  LUT3 #(.INIT(8'h96)) lut_n1992 (.I0(x198), .I1(x199), .I2(x200), .O(n1992));
  LUT5 #(.INIT(32'h96696996)) lut_n1993 (.I0(x189), .I1(x190), .I2(x191), .I3(n1987), .I4(n1988), .O(n1993));
  LUT5 #(.INIT(32'hFF969600)) lut_n1994 (.I0(x195), .I1(x196), .I2(x197), .I3(n1992), .I4(n1993), .O(n1994));
  LUT3 #(.INIT(8'h96)) lut_n1995 (.I0(x204), .I1(x205), .I2(x206), .O(n1995));
  LUT5 #(.INIT(32'h96696996)) lut_n1996 (.I0(x195), .I1(x196), .I2(x197), .I3(n1992), .I4(n1993), .O(n1996));
  LUT5 #(.INIT(32'hFF969600)) lut_n1997 (.I0(x201), .I1(x202), .I2(x203), .I3(n1995), .I4(n1996), .O(n1997));
  LUT3 #(.INIT(8'h96)) lut_n1998 (.I0(n1986), .I1(n1989), .I2(n1990), .O(n1998));
  LUT3 #(.INIT(8'hE8)) lut_n1999 (.I0(n1994), .I1(n1997), .I2(n1998), .O(n1999));
  LUT3 #(.INIT(8'h96)) lut_n2000 (.I0(n1973), .I1(n1981), .I2(n1982), .O(n2000));
  LUT3 #(.INIT(8'h8E)) lut_n2001 (.I0(n1991), .I1(n1999), .I2(n2000), .O(n2001));
  LUT3 #(.INIT(8'h96)) lut_n2002 (.I0(n1943), .I1(n1961), .I2(n1962), .O(n2002));
  LUT3 #(.INIT(8'hE8)) lut_n2003 (.I0(n1983), .I1(n2001), .I2(n2002), .O(n2003));
  LUT3 #(.INIT(8'h96)) lut_n2004 (.I0(x210), .I1(x211), .I2(x212), .O(n2004));
  LUT5 #(.INIT(32'h96696996)) lut_n2005 (.I0(x201), .I1(x202), .I2(x203), .I3(n1995), .I4(n1996), .O(n2005));
  LUT5 #(.INIT(32'hFF969600)) lut_n2006 (.I0(x207), .I1(x208), .I2(x209), .I3(n2004), .I4(n2005), .O(n2006));
  LUT3 #(.INIT(8'h96)) lut_n2007 (.I0(x216), .I1(x217), .I2(x218), .O(n2007));
  LUT5 #(.INIT(32'h96696996)) lut_n2008 (.I0(x207), .I1(x208), .I2(x209), .I3(n2004), .I4(n2005), .O(n2008));
  LUT5 #(.INIT(32'hFF969600)) lut_n2009 (.I0(x213), .I1(x214), .I2(x215), .I3(n2007), .I4(n2008), .O(n2009));
  LUT3 #(.INIT(8'h96)) lut_n2010 (.I0(n1994), .I1(n1997), .I2(n1998), .O(n2010));
  LUT3 #(.INIT(8'hE8)) lut_n2011 (.I0(n2006), .I1(n2009), .I2(n2010), .O(n2011));
  LUT3 #(.INIT(8'h96)) lut_n2012 (.I0(x222), .I1(x223), .I2(x224), .O(n2012));
  LUT5 #(.INIT(32'h96696996)) lut_n2013 (.I0(x213), .I1(x214), .I2(x215), .I3(n2007), .I4(n2008), .O(n2013));
  LUT5 #(.INIT(32'hFF969600)) lut_n2014 (.I0(x219), .I1(x220), .I2(x221), .I3(n2012), .I4(n2013), .O(n2014));
  LUT3 #(.INIT(8'h96)) lut_n2015 (.I0(x228), .I1(x229), .I2(x230), .O(n2015));
  LUT5 #(.INIT(32'h96696996)) lut_n2016 (.I0(x219), .I1(x220), .I2(x221), .I3(n2012), .I4(n2013), .O(n2016));
  LUT5 #(.INIT(32'hFF969600)) lut_n2017 (.I0(x225), .I1(x226), .I2(x227), .I3(n2015), .I4(n2016), .O(n2017));
  LUT3 #(.INIT(8'h96)) lut_n2018 (.I0(n2006), .I1(n2009), .I2(n2010), .O(n2018));
  LUT3 #(.INIT(8'hE8)) lut_n2019 (.I0(n2014), .I1(n2017), .I2(n2018), .O(n2019));
  LUT3 #(.INIT(8'h96)) lut_n2020 (.I0(n1991), .I1(n1999), .I2(n2000), .O(n2020));
  LUT3 #(.INIT(8'h8E)) lut_n2021 (.I0(n2011), .I1(n2019), .I2(n2020), .O(n2021));
  LUT3 #(.INIT(8'h96)) lut_n2022 (.I0(x234), .I1(x235), .I2(x236), .O(n2022));
  LUT5 #(.INIT(32'h96696996)) lut_n2023 (.I0(x225), .I1(x226), .I2(x227), .I3(n2015), .I4(n2016), .O(n2023));
  LUT5 #(.INIT(32'hFF969600)) lut_n2024 (.I0(x231), .I1(x232), .I2(x233), .I3(n2022), .I4(n2023), .O(n2024));
  LUT3 #(.INIT(8'h96)) lut_n2025 (.I0(x240), .I1(x241), .I2(x242), .O(n2025));
  LUT5 #(.INIT(32'h96696996)) lut_n2026 (.I0(x231), .I1(x232), .I2(x233), .I3(n2022), .I4(n2023), .O(n2026));
  LUT5 #(.INIT(32'hFF969600)) lut_n2027 (.I0(x237), .I1(x238), .I2(x239), .I3(n2025), .I4(n2026), .O(n2027));
  LUT3 #(.INIT(8'h96)) lut_n2028 (.I0(n2014), .I1(n2017), .I2(n2018), .O(n2028));
  LUT3 #(.INIT(8'hE8)) lut_n2029 (.I0(n2024), .I1(n2027), .I2(n2028), .O(n2029));
  LUT3 #(.INIT(8'h96)) lut_n2030 (.I0(x246), .I1(x247), .I2(x248), .O(n2030));
  LUT5 #(.INIT(32'h96696996)) lut_n2031 (.I0(x237), .I1(x238), .I2(x239), .I3(n2025), .I4(n2026), .O(n2031));
  LUT5 #(.INIT(32'hFF969600)) lut_n2032 (.I0(x243), .I1(x244), .I2(x245), .I3(n2030), .I4(n2031), .O(n2032));
  LUT3 #(.INIT(8'h96)) lut_n2033 (.I0(x252), .I1(x253), .I2(x254), .O(n2033));
  LUT5 #(.INIT(32'h96696996)) lut_n2034 (.I0(x243), .I1(x244), .I2(x245), .I3(n2030), .I4(n2031), .O(n2034));
  LUT5 #(.INIT(32'hFF969600)) lut_n2035 (.I0(x249), .I1(x250), .I2(x251), .I3(n2033), .I4(n2034), .O(n2035));
  LUT3 #(.INIT(8'h96)) lut_n2036 (.I0(n2024), .I1(n2027), .I2(n2028), .O(n2036));
  LUT3 #(.INIT(8'hE8)) lut_n2037 (.I0(n2032), .I1(n2035), .I2(n2036), .O(n2037));
  LUT3 #(.INIT(8'h96)) lut_n2038 (.I0(n2011), .I1(n2019), .I2(n2020), .O(n2038));
  LUT3 #(.INIT(8'h8E)) lut_n2039 (.I0(n2029), .I1(n2037), .I2(n2038), .O(n2039));
  LUT3 #(.INIT(8'h96)) lut_n2040 (.I0(n1983), .I1(n2001), .I2(n2002), .O(n2040));
  LUT3 #(.INIT(8'hE8)) lut_n2041 (.I0(n2021), .I1(n2039), .I2(n2040), .O(n2041));
  LUT3 #(.INIT(8'h96)) lut_n2042 (.I0(n1925), .I1(n1963), .I2(n1964), .O(n2042));
  LUT3 #(.INIT(8'hE8)) lut_n2043 (.I0(n2003), .I1(n2041), .I2(n2042), .O(n2043));
  LUT3 #(.INIT(8'h96)) lut_n2044 (.I0(n1826), .I1(n1885), .I2(n1886), .O(n2044));
  LUT3 #(.INIT(8'hE8)) lut_n2045 (.I0(n1965), .I1(n2043), .I2(n2044), .O(n2045));
  LUT3 #(.INIT(8'h96)) lut_n2046 (.I0(n1708), .I1(n1786), .I2(n1787), .O(n2046));
  LUT3 #(.INIT(8'hE8)) lut_n2047 (.I0(n1887), .I1(n2045), .I2(n2046), .O(n2047));
  LUT3 #(.INIT(8'h96)) lut_n2048 (.I0(n1314), .I1(n1472), .I2(n1630), .O(n2048));
  LUT3 #(.INIT(8'hE8)) lut_n2049 (.I0(n1788), .I1(n2047), .I2(n2048), .O(n2049));
  LUT3 #(.INIT(8'h96)) lut_n2050 (.I0(x258), .I1(x259), .I2(x260), .O(n2050));
  LUT5 #(.INIT(32'h96696996)) lut_n2051 (.I0(x249), .I1(x250), .I2(x251), .I3(n2033), .I4(n2034), .O(n2051));
  LUT5 #(.INIT(32'hFF969600)) lut_n2052 (.I0(x255), .I1(x256), .I2(x257), .I3(n2050), .I4(n2051), .O(n2052));
  LUT3 #(.INIT(8'h96)) lut_n2053 (.I0(x264), .I1(x265), .I2(x266), .O(n2053));
  LUT5 #(.INIT(32'h96696996)) lut_n2054 (.I0(x255), .I1(x256), .I2(x257), .I3(n2050), .I4(n2051), .O(n2054));
  LUT5 #(.INIT(32'hFF969600)) lut_n2055 (.I0(x261), .I1(x262), .I2(x263), .I3(n2053), .I4(n2054), .O(n2055));
  LUT3 #(.INIT(8'h96)) lut_n2056 (.I0(n2032), .I1(n2035), .I2(n2036), .O(n2056));
  LUT3 #(.INIT(8'hE8)) lut_n2057 (.I0(n2052), .I1(n2055), .I2(n2056), .O(n2057));
  LUT3 #(.INIT(8'h96)) lut_n2058 (.I0(x270), .I1(x271), .I2(x272), .O(n2058));
  LUT5 #(.INIT(32'h96696996)) lut_n2059 (.I0(x261), .I1(x262), .I2(x263), .I3(n2053), .I4(n2054), .O(n2059));
  LUT5 #(.INIT(32'hFF969600)) lut_n2060 (.I0(x267), .I1(x268), .I2(x269), .I3(n2058), .I4(n2059), .O(n2060));
  LUT3 #(.INIT(8'h96)) lut_n2061 (.I0(x276), .I1(x277), .I2(x278), .O(n2061));
  LUT5 #(.INIT(32'h96696996)) lut_n2062 (.I0(x267), .I1(x268), .I2(x269), .I3(n2058), .I4(n2059), .O(n2062));
  LUT5 #(.INIT(32'hFF969600)) lut_n2063 (.I0(x273), .I1(x274), .I2(x275), .I3(n2061), .I4(n2062), .O(n2063));
  LUT3 #(.INIT(8'h96)) lut_n2064 (.I0(n2052), .I1(n2055), .I2(n2056), .O(n2064));
  LUT3 #(.INIT(8'hE8)) lut_n2065 (.I0(n2060), .I1(n2063), .I2(n2064), .O(n2065));
  LUT3 #(.INIT(8'h96)) lut_n2066 (.I0(n2029), .I1(n2037), .I2(n2038), .O(n2066));
  LUT3 #(.INIT(8'h8E)) lut_n2067 (.I0(n2057), .I1(n2065), .I2(n2066), .O(n2067));
  LUT3 #(.INIT(8'h96)) lut_n2068 (.I0(x282), .I1(x283), .I2(x284), .O(n2068));
  LUT5 #(.INIT(32'h96696996)) lut_n2069 (.I0(x273), .I1(x274), .I2(x275), .I3(n2061), .I4(n2062), .O(n2069));
  LUT5 #(.INIT(32'hFF969600)) lut_n2070 (.I0(x279), .I1(x280), .I2(x281), .I3(n2068), .I4(n2069), .O(n2070));
  LUT3 #(.INIT(8'h96)) lut_n2071 (.I0(x288), .I1(x289), .I2(x290), .O(n2071));
  LUT5 #(.INIT(32'h96696996)) lut_n2072 (.I0(x279), .I1(x280), .I2(x281), .I3(n2068), .I4(n2069), .O(n2072));
  LUT5 #(.INIT(32'hFF969600)) lut_n2073 (.I0(x285), .I1(x286), .I2(x287), .I3(n2071), .I4(n2072), .O(n2073));
  LUT3 #(.INIT(8'h96)) lut_n2074 (.I0(n2060), .I1(n2063), .I2(n2064), .O(n2074));
  LUT3 #(.INIT(8'hE8)) lut_n2075 (.I0(n2070), .I1(n2073), .I2(n2074), .O(n2075));
  LUT3 #(.INIT(8'h96)) lut_n2076 (.I0(x294), .I1(x295), .I2(x296), .O(n2076));
  LUT5 #(.INIT(32'h96696996)) lut_n2077 (.I0(x285), .I1(x286), .I2(x287), .I3(n2071), .I4(n2072), .O(n2077));
  LUT5 #(.INIT(32'hFF969600)) lut_n2078 (.I0(x291), .I1(x292), .I2(x293), .I3(n2076), .I4(n2077), .O(n2078));
  LUT3 #(.INIT(8'h96)) lut_n2079 (.I0(x297), .I1(x298), .I2(x299), .O(n2079));
  LUT5 #(.INIT(32'h96696996)) lut_n2080 (.I0(x291), .I1(x292), .I2(x293), .I3(n2076), .I4(n2077), .O(n2080));
  LUT5 #(.INIT(32'hFF969600)) lut_n2081 (.I0(x300), .I1(x301), .I2(x302), .I3(n2079), .I4(n2080), .O(n2081));
  LUT3 #(.INIT(8'h96)) lut_n2082 (.I0(n2070), .I1(n2073), .I2(n2074), .O(n2082));
  LUT3 #(.INIT(8'hE8)) lut_n2083 (.I0(n2078), .I1(n2081), .I2(n2082), .O(n2083));
  LUT3 #(.INIT(8'h96)) lut_n2084 (.I0(n2057), .I1(n2065), .I2(n2066), .O(n2084));
  LUT3 #(.INIT(8'h8E)) lut_n2085 (.I0(n2075), .I1(n2083), .I2(n2084), .O(n2085));
  LUT3 #(.INIT(8'h96)) lut_n2086 (.I0(n2021), .I1(n2039), .I2(n2040), .O(n2086));
  LUT3 #(.INIT(8'hE8)) lut_n2087 (.I0(n2067), .I1(n2085), .I2(n2086), .O(n2087));
  LUT3 #(.INIT(8'h96)) lut_n2088 (.I0(x306), .I1(x307), .I2(x308), .O(n2088));
  LUT5 #(.INIT(32'h96696996)) lut_n2089 (.I0(x300), .I1(x301), .I2(x302), .I3(n2079), .I4(n2080), .O(n2089));
  LUT5 #(.INIT(32'hFF969600)) lut_n2090 (.I0(x303), .I1(x304), .I2(x305), .I3(n2088), .I4(n2089), .O(n2090));
  LUT3 #(.INIT(8'h96)) lut_n2091 (.I0(x312), .I1(x313), .I2(x314), .O(n2091));
  LUT5 #(.INIT(32'h96696996)) lut_n2092 (.I0(x303), .I1(x304), .I2(x305), .I3(n2088), .I4(n2089), .O(n2092));
  LUT5 #(.INIT(32'hFF969600)) lut_n2093 (.I0(x309), .I1(x310), .I2(x311), .I3(n2091), .I4(n2092), .O(n2093));
  LUT3 #(.INIT(8'h96)) lut_n2094 (.I0(n2078), .I1(n2081), .I2(n2082), .O(n2094));
  LUT3 #(.INIT(8'hE8)) lut_n2095 (.I0(n2090), .I1(n2093), .I2(n2094), .O(n2095));
  LUT3 #(.INIT(8'h96)) lut_n2096 (.I0(x318), .I1(x319), .I2(x320), .O(n2096));
  LUT5 #(.INIT(32'h96696996)) lut_n2097 (.I0(x309), .I1(x310), .I2(x311), .I3(n2091), .I4(n2092), .O(n2097));
  LUT5 #(.INIT(32'hFF969600)) lut_n2098 (.I0(x315), .I1(x316), .I2(x317), .I3(n2096), .I4(n2097), .O(n2098));
  LUT3 #(.INIT(8'h96)) lut_n2099 (.I0(x324), .I1(x325), .I2(x326), .O(n2099));
  LUT5 #(.INIT(32'h96696996)) lut_n2100 (.I0(x315), .I1(x316), .I2(x317), .I3(n2096), .I4(n2097), .O(n2100));
  LUT5 #(.INIT(32'hFF969600)) lut_n2101 (.I0(x321), .I1(x322), .I2(x323), .I3(n2099), .I4(n2100), .O(n2101));
  LUT3 #(.INIT(8'h96)) lut_n2102 (.I0(n2090), .I1(n2093), .I2(n2094), .O(n2102));
  LUT3 #(.INIT(8'hE8)) lut_n2103 (.I0(n2098), .I1(n2101), .I2(n2102), .O(n2103));
  LUT3 #(.INIT(8'h96)) lut_n2104 (.I0(n2075), .I1(n2083), .I2(n2084), .O(n2104));
  LUT3 #(.INIT(8'h8E)) lut_n2105 (.I0(n2095), .I1(n2103), .I2(n2104), .O(n2105));
  LUT3 #(.INIT(8'h96)) lut_n2106 (.I0(x330), .I1(x331), .I2(x332), .O(n2106));
  LUT5 #(.INIT(32'h96696996)) lut_n2107 (.I0(x321), .I1(x322), .I2(x323), .I3(n2099), .I4(n2100), .O(n2107));
  LUT5 #(.INIT(32'hFF969600)) lut_n2108 (.I0(x327), .I1(x328), .I2(x329), .I3(n2106), .I4(n2107), .O(n2108));
  LUT3 #(.INIT(8'h96)) lut_n2109 (.I0(x336), .I1(x337), .I2(x338), .O(n2109));
  LUT5 #(.INIT(32'h96696996)) lut_n2110 (.I0(x327), .I1(x328), .I2(x329), .I3(n2106), .I4(n2107), .O(n2110));
  LUT5 #(.INIT(32'hFF969600)) lut_n2111 (.I0(x333), .I1(x334), .I2(x335), .I3(n2109), .I4(n2110), .O(n2111));
  LUT3 #(.INIT(8'h96)) lut_n2112 (.I0(n2098), .I1(n2101), .I2(n2102), .O(n2112));
  LUT3 #(.INIT(8'hE8)) lut_n2113 (.I0(n2108), .I1(n2111), .I2(n2112), .O(n2113));
  LUT3 #(.INIT(8'h96)) lut_n2114 (.I0(x342), .I1(x343), .I2(x344), .O(n2114));
  LUT5 #(.INIT(32'h96696996)) lut_n2115 (.I0(x333), .I1(x334), .I2(x335), .I3(n2109), .I4(n2110), .O(n2115));
  LUT5 #(.INIT(32'hFF969600)) lut_n2116 (.I0(x339), .I1(x340), .I2(x341), .I3(n2114), .I4(n2115), .O(n2116));
  LUT3 #(.INIT(8'h96)) lut_n2117 (.I0(x348), .I1(x349), .I2(x350), .O(n2117));
  LUT5 #(.INIT(32'h96696996)) lut_n2118 (.I0(x339), .I1(x340), .I2(x341), .I3(n2114), .I4(n2115), .O(n2118));
  LUT5 #(.INIT(32'hFF969600)) lut_n2119 (.I0(x345), .I1(x346), .I2(x347), .I3(n2117), .I4(n2118), .O(n2119));
  LUT3 #(.INIT(8'h96)) lut_n2120 (.I0(n2108), .I1(n2111), .I2(n2112), .O(n2120));
  LUT3 #(.INIT(8'hE8)) lut_n2121 (.I0(n2116), .I1(n2119), .I2(n2120), .O(n2121));
  LUT3 #(.INIT(8'h96)) lut_n2122 (.I0(n2095), .I1(n2103), .I2(n2104), .O(n2122));
  LUT3 #(.INIT(8'h8E)) lut_n2123 (.I0(n2113), .I1(n2121), .I2(n2122), .O(n2123));
  LUT3 #(.INIT(8'h96)) lut_n2124 (.I0(n2067), .I1(n2085), .I2(n2086), .O(n2124));
  LUT3 #(.INIT(8'hE8)) lut_n2125 (.I0(n2105), .I1(n2123), .I2(n2124), .O(n2125));
  LUT3 #(.INIT(8'h96)) lut_n2126 (.I0(n2003), .I1(n2041), .I2(n2042), .O(n2126));
  LUT3 #(.INIT(8'hE8)) lut_n2127 (.I0(n2087), .I1(n2125), .I2(n2126), .O(n2127));
  LUT3 #(.INIT(8'h96)) lut_n2128 (.I0(x354), .I1(x355), .I2(x356), .O(n2128));
  LUT5 #(.INIT(32'h96696996)) lut_n2129 (.I0(x345), .I1(x346), .I2(x347), .I3(n2117), .I4(n2118), .O(n2129));
  LUT5 #(.INIT(32'hFF969600)) lut_n2130 (.I0(x351), .I1(x352), .I2(x353), .I3(n2128), .I4(n2129), .O(n2130));
  LUT3 #(.INIT(8'h96)) lut_n2131 (.I0(x360), .I1(x361), .I2(x362), .O(n2131));
  LUT5 #(.INIT(32'h96696996)) lut_n2132 (.I0(x351), .I1(x352), .I2(x353), .I3(n2128), .I4(n2129), .O(n2132));
  LUT5 #(.INIT(32'hFF969600)) lut_n2133 (.I0(x357), .I1(x358), .I2(x359), .I3(n2131), .I4(n2132), .O(n2133));
  LUT3 #(.INIT(8'h96)) lut_n2134 (.I0(n2116), .I1(n2119), .I2(n2120), .O(n2134));
  LUT3 #(.INIT(8'hE8)) lut_n2135 (.I0(n2130), .I1(n2133), .I2(n2134), .O(n2135));
  LUT3 #(.INIT(8'h96)) lut_n2136 (.I0(x366), .I1(x367), .I2(x368), .O(n2136));
  LUT5 #(.INIT(32'h96696996)) lut_n2137 (.I0(x357), .I1(x358), .I2(x359), .I3(n2131), .I4(n2132), .O(n2137));
  LUT5 #(.INIT(32'hFF969600)) lut_n2138 (.I0(x363), .I1(x364), .I2(x365), .I3(n2136), .I4(n2137), .O(n2138));
  LUT3 #(.INIT(8'h96)) lut_n2139 (.I0(x372), .I1(x373), .I2(x374), .O(n2139));
  LUT5 #(.INIT(32'h96696996)) lut_n2140 (.I0(x363), .I1(x364), .I2(x365), .I3(n2136), .I4(n2137), .O(n2140));
  LUT5 #(.INIT(32'hFF969600)) lut_n2141 (.I0(x369), .I1(x370), .I2(x371), .I3(n2139), .I4(n2140), .O(n2141));
  LUT3 #(.INIT(8'h96)) lut_n2142 (.I0(n2130), .I1(n2133), .I2(n2134), .O(n2142));
  LUT3 #(.INIT(8'hE8)) lut_n2143 (.I0(n2138), .I1(n2141), .I2(n2142), .O(n2143));
  LUT3 #(.INIT(8'h96)) lut_n2144 (.I0(n2113), .I1(n2121), .I2(n2122), .O(n2144));
  LUT3 #(.INIT(8'h8E)) lut_n2145 (.I0(n2135), .I1(n2143), .I2(n2144), .O(n2145));
  LUT3 #(.INIT(8'h96)) lut_n2146 (.I0(x378), .I1(x379), .I2(x380), .O(n2146));
  LUT5 #(.INIT(32'h96696996)) lut_n2147 (.I0(x369), .I1(x370), .I2(x371), .I3(n2139), .I4(n2140), .O(n2147));
  LUT5 #(.INIT(32'hFF969600)) lut_n2148 (.I0(x375), .I1(x376), .I2(x377), .I3(n2146), .I4(n2147), .O(n2148));
  LUT3 #(.INIT(8'h96)) lut_n2149 (.I0(x384), .I1(x385), .I2(x386), .O(n2149));
  LUT5 #(.INIT(32'h96696996)) lut_n2150 (.I0(x375), .I1(x376), .I2(x377), .I3(n2146), .I4(n2147), .O(n2150));
  LUT5 #(.INIT(32'hFF969600)) lut_n2151 (.I0(x381), .I1(x382), .I2(x383), .I3(n2149), .I4(n2150), .O(n2151));
  LUT3 #(.INIT(8'h96)) lut_n2152 (.I0(n2138), .I1(n2141), .I2(n2142), .O(n2152));
  LUT3 #(.INIT(8'hE8)) lut_n2153 (.I0(n2148), .I1(n2151), .I2(n2152), .O(n2153));
  LUT3 #(.INIT(8'h96)) lut_n2154 (.I0(x390), .I1(x391), .I2(x392), .O(n2154));
  LUT5 #(.INIT(32'h96696996)) lut_n2155 (.I0(x381), .I1(x382), .I2(x383), .I3(n2149), .I4(n2150), .O(n2155));
  LUT5 #(.INIT(32'hFF969600)) lut_n2156 (.I0(x387), .I1(x388), .I2(x389), .I3(n2154), .I4(n2155), .O(n2156));
  LUT3 #(.INIT(8'h96)) lut_n2157 (.I0(x396), .I1(x397), .I2(x398), .O(n2157));
  LUT5 #(.INIT(32'h96696996)) lut_n2158 (.I0(x387), .I1(x388), .I2(x389), .I3(n2154), .I4(n2155), .O(n2158));
  LUT5 #(.INIT(32'hFF969600)) lut_n2159 (.I0(x393), .I1(x394), .I2(x395), .I3(n2157), .I4(n2158), .O(n2159));
  LUT3 #(.INIT(8'h96)) lut_n2160 (.I0(n2148), .I1(n2151), .I2(n2152), .O(n2160));
  LUT3 #(.INIT(8'hE8)) lut_n2161 (.I0(n2156), .I1(n2159), .I2(n2160), .O(n2161));
  LUT3 #(.INIT(8'h96)) lut_n2162 (.I0(n2135), .I1(n2143), .I2(n2144), .O(n2162));
  LUT3 #(.INIT(8'h8E)) lut_n2163 (.I0(n2153), .I1(n2161), .I2(n2162), .O(n2163));
  LUT3 #(.INIT(8'h96)) lut_n2164 (.I0(n2105), .I1(n2123), .I2(n2124), .O(n2164));
  LUT3 #(.INIT(8'hE8)) lut_n2165 (.I0(n2145), .I1(n2163), .I2(n2164), .O(n2165));
  LUT3 #(.INIT(8'h96)) lut_n2166 (.I0(x402), .I1(x403), .I2(x404), .O(n2166));
  LUT5 #(.INIT(32'h96696996)) lut_n2167 (.I0(x393), .I1(x394), .I2(x395), .I3(n2157), .I4(n2158), .O(n2167));
  LUT5 #(.INIT(32'hFF969600)) lut_n2168 (.I0(x399), .I1(x400), .I2(x401), .I3(n2166), .I4(n2167), .O(n2168));
  LUT3 #(.INIT(8'h96)) lut_n2169 (.I0(x408), .I1(x409), .I2(x410), .O(n2169));
  LUT5 #(.INIT(32'h96696996)) lut_n2170 (.I0(x399), .I1(x400), .I2(x401), .I3(n2166), .I4(n2167), .O(n2170));
  LUT5 #(.INIT(32'hFF969600)) lut_n2171 (.I0(x405), .I1(x406), .I2(x407), .I3(n2169), .I4(n2170), .O(n2171));
  LUT3 #(.INIT(8'h96)) lut_n2172 (.I0(n2156), .I1(n2159), .I2(n2160), .O(n2172));
  LUT3 #(.INIT(8'hE8)) lut_n2173 (.I0(n2168), .I1(n2171), .I2(n2172), .O(n2173));
  LUT3 #(.INIT(8'h96)) lut_n2174 (.I0(x414), .I1(x415), .I2(x416), .O(n2174));
  LUT5 #(.INIT(32'h96696996)) lut_n2175 (.I0(x405), .I1(x406), .I2(x407), .I3(n2169), .I4(n2170), .O(n2175));
  LUT5 #(.INIT(32'hFF969600)) lut_n2176 (.I0(x411), .I1(x412), .I2(x413), .I3(n2174), .I4(n2175), .O(n2176));
  LUT3 #(.INIT(8'h96)) lut_n2177 (.I0(x420), .I1(x421), .I2(x422), .O(n2177));
  LUT5 #(.INIT(32'h96696996)) lut_n2178 (.I0(x411), .I1(x412), .I2(x413), .I3(n2174), .I4(n2175), .O(n2178));
  LUT5 #(.INIT(32'hFF969600)) lut_n2179 (.I0(x417), .I1(x418), .I2(x419), .I3(n2177), .I4(n2178), .O(n2179));
  LUT3 #(.INIT(8'h96)) lut_n2180 (.I0(n2168), .I1(n2171), .I2(n2172), .O(n2180));
  LUT3 #(.INIT(8'hE8)) lut_n2181 (.I0(n2176), .I1(n2179), .I2(n2180), .O(n2181));
  LUT3 #(.INIT(8'h96)) lut_n2182 (.I0(n2153), .I1(n2161), .I2(n2162), .O(n2182));
  LUT3 #(.INIT(8'h8E)) lut_n2183 (.I0(n2173), .I1(n2181), .I2(n2182), .O(n2183));
  LUT3 #(.INIT(8'h96)) lut_n2184 (.I0(x426), .I1(x427), .I2(x428), .O(n2184));
  LUT5 #(.INIT(32'h96696996)) lut_n2185 (.I0(x417), .I1(x418), .I2(x419), .I3(n2177), .I4(n2178), .O(n2185));
  LUT5 #(.INIT(32'hFF969600)) lut_n2186 (.I0(x423), .I1(x424), .I2(x425), .I3(n2184), .I4(n2185), .O(n2186));
  LUT3 #(.INIT(8'h96)) lut_n2187 (.I0(x432), .I1(x433), .I2(x434), .O(n2187));
  LUT5 #(.INIT(32'h96696996)) lut_n2188 (.I0(x423), .I1(x424), .I2(x425), .I3(n2184), .I4(n2185), .O(n2188));
  LUT5 #(.INIT(32'hFF969600)) lut_n2189 (.I0(x429), .I1(x430), .I2(x431), .I3(n2187), .I4(n2188), .O(n2189));
  LUT3 #(.INIT(8'h96)) lut_n2190 (.I0(n2176), .I1(n2179), .I2(n2180), .O(n2190));
  LUT3 #(.INIT(8'hE8)) lut_n2191 (.I0(n2186), .I1(n2189), .I2(n2190), .O(n2191));
  LUT3 #(.INIT(8'h96)) lut_n2192 (.I0(x438), .I1(x439), .I2(x440), .O(n2192));
  LUT5 #(.INIT(32'h96696996)) lut_n2193 (.I0(x429), .I1(x430), .I2(x431), .I3(n2187), .I4(n2188), .O(n2193));
  LUT5 #(.INIT(32'hFF969600)) lut_n2194 (.I0(x435), .I1(x436), .I2(x437), .I3(n2192), .I4(n2193), .O(n2194));
  LUT3 #(.INIT(8'h96)) lut_n2195 (.I0(x444), .I1(x445), .I2(x446), .O(n2195));
  LUT5 #(.INIT(32'h96696996)) lut_n2196 (.I0(x435), .I1(x436), .I2(x437), .I3(n2192), .I4(n2193), .O(n2196));
  LUT5 #(.INIT(32'hFF969600)) lut_n2197 (.I0(x441), .I1(x442), .I2(x443), .I3(n2195), .I4(n2196), .O(n2197));
  LUT3 #(.INIT(8'h96)) lut_n2198 (.I0(n2186), .I1(n2189), .I2(n2190), .O(n2198));
  LUT3 #(.INIT(8'hE8)) lut_n2199 (.I0(n2194), .I1(n2197), .I2(n2198), .O(n2199));
  LUT3 #(.INIT(8'h96)) lut_n2200 (.I0(n2173), .I1(n2181), .I2(n2182), .O(n2200));
  LUT3 #(.INIT(8'h8E)) lut_n2201 (.I0(n2191), .I1(n2199), .I2(n2200), .O(n2201));
  LUT3 #(.INIT(8'h96)) lut_n2202 (.I0(n2145), .I1(n2163), .I2(n2164), .O(n2202));
  LUT3 #(.INIT(8'hE8)) lut_n2203 (.I0(n2183), .I1(n2201), .I2(n2202), .O(n2203));
  LUT3 #(.INIT(8'h96)) lut_n2204 (.I0(n2087), .I1(n2125), .I2(n2126), .O(n2204));
  LUT3 #(.INIT(8'hE8)) lut_n2205 (.I0(n2165), .I1(n2203), .I2(n2204), .O(n2205));
  LUT3 #(.INIT(8'h96)) lut_n2206 (.I0(n1965), .I1(n2043), .I2(n2044), .O(n2206));
  LUT3 #(.INIT(8'hE8)) lut_n2207 (.I0(n2127), .I1(n2205), .I2(n2206), .O(n2207));
  LUT3 #(.INIT(8'h96)) lut_n2208 (.I0(x450), .I1(x451), .I2(x452), .O(n2208));
  LUT5 #(.INIT(32'h96696996)) lut_n2209 (.I0(x441), .I1(x442), .I2(x443), .I3(n2195), .I4(n2196), .O(n2209));
  LUT5 #(.INIT(32'hFF969600)) lut_n2210 (.I0(x447), .I1(x448), .I2(x449), .I3(n2208), .I4(n2209), .O(n2210));
  LUT3 #(.INIT(8'h96)) lut_n2211 (.I0(x456), .I1(x457), .I2(x458), .O(n2211));
  LUT5 #(.INIT(32'h96696996)) lut_n2212 (.I0(x447), .I1(x448), .I2(x449), .I3(n2208), .I4(n2209), .O(n2212));
  LUT5 #(.INIT(32'hFF969600)) lut_n2213 (.I0(x453), .I1(x454), .I2(x455), .I3(n2211), .I4(n2212), .O(n2213));
  LUT3 #(.INIT(8'h96)) lut_n2214 (.I0(n2194), .I1(n2197), .I2(n2198), .O(n2214));
  LUT3 #(.INIT(8'hE8)) lut_n2215 (.I0(n2210), .I1(n2213), .I2(n2214), .O(n2215));
  LUT3 #(.INIT(8'h96)) lut_n2216 (.I0(x462), .I1(x463), .I2(x464), .O(n2216));
  LUT5 #(.INIT(32'h96696996)) lut_n2217 (.I0(x453), .I1(x454), .I2(x455), .I3(n2211), .I4(n2212), .O(n2217));
  LUT5 #(.INIT(32'hFF969600)) lut_n2218 (.I0(x459), .I1(x460), .I2(x461), .I3(n2216), .I4(n2217), .O(n2218));
  LUT3 #(.INIT(8'h96)) lut_n2219 (.I0(x468), .I1(x469), .I2(x470), .O(n2219));
  LUT5 #(.INIT(32'h96696996)) lut_n2220 (.I0(x459), .I1(x460), .I2(x461), .I3(n2216), .I4(n2217), .O(n2220));
  LUT5 #(.INIT(32'hFF969600)) lut_n2221 (.I0(x465), .I1(x466), .I2(x467), .I3(n2219), .I4(n2220), .O(n2221));
  LUT3 #(.INIT(8'h96)) lut_n2222 (.I0(n2210), .I1(n2213), .I2(n2214), .O(n2222));
  LUT3 #(.INIT(8'hE8)) lut_n2223 (.I0(n2218), .I1(n2221), .I2(n2222), .O(n2223));
  LUT3 #(.INIT(8'h96)) lut_n2224 (.I0(n2191), .I1(n2199), .I2(n2200), .O(n2224));
  LUT3 #(.INIT(8'h8E)) lut_n2225 (.I0(n2215), .I1(n2223), .I2(n2224), .O(n2225));
  LUT3 #(.INIT(8'h96)) lut_n2226 (.I0(x474), .I1(x475), .I2(x476), .O(n2226));
  LUT5 #(.INIT(32'h96696996)) lut_n2227 (.I0(x465), .I1(x466), .I2(x467), .I3(n2219), .I4(n2220), .O(n2227));
  LUT5 #(.INIT(32'hFF969600)) lut_n2228 (.I0(x471), .I1(x472), .I2(x473), .I3(n2226), .I4(n2227), .O(n2228));
  LUT3 #(.INIT(8'h96)) lut_n2229 (.I0(x480), .I1(x481), .I2(x482), .O(n2229));
  LUT5 #(.INIT(32'h96696996)) lut_n2230 (.I0(x471), .I1(x472), .I2(x473), .I3(n2226), .I4(n2227), .O(n2230));
  LUT5 #(.INIT(32'hFF969600)) lut_n2231 (.I0(x477), .I1(x478), .I2(x479), .I3(n2229), .I4(n2230), .O(n2231));
  LUT3 #(.INIT(8'h96)) lut_n2232 (.I0(n2218), .I1(n2221), .I2(n2222), .O(n2232));
  LUT3 #(.INIT(8'hE8)) lut_n2233 (.I0(n2228), .I1(n2231), .I2(n2232), .O(n2233));
  LUT3 #(.INIT(8'h96)) lut_n2234 (.I0(x486), .I1(x487), .I2(x488), .O(n2234));
  LUT5 #(.INIT(32'h96696996)) lut_n2235 (.I0(x477), .I1(x478), .I2(x479), .I3(n2229), .I4(n2230), .O(n2235));
  LUT5 #(.INIT(32'hFF969600)) lut_n2236 (.I0(x483), .I1(x484), .I2(x485), .I3(n2234), .I4(n2235), .O(n2236));
  LUT3 #(.INIT(8'h96)) lut_n2237 (.I0(x492), .I1(x493), .I2(x494), .O(n2237));
  LUT5 #(.INIT(32'h96696996)) lut_n2238 (.I0(x483), .I1(x484), .I2(x485), .I3(n2234), .I4(n2235), .O(n2238));
  LUT5 #(.INIT(32'hFF969600)) lut_n2239 (.I0(x489), .I1(x490), .I2(x491), .I3(n2237), .I4(n2238), .O(n2239));
  LUT3 #(.INIT(8'h96)) lut_n2240 (.I0(n2228), .I1(n2231), .I2(n2232), .O(n2240));
  LUT3 #(.INIT(8'hE8)) lut_n2241 (.I0(n2236), .I1(n2239), .I2(n2240), .O(n2241));
  LUT3 #(.INIT(8'h96)) lut_n2242 (.I0(n2215), .I1(n2223), .I2(n2224), .O(n2242));
  LUT3 #(.INIT(8'h8E)) lut_n2243 (.I0(n2233), .I1(n2241), .I2(n2242), .O(n2243));
  LUT3 #(.INIT(8'h96)) lut_n2244 (.I0(n2183), .I1(n2201), .I2(n2202), .O(n2244));
  LUT3 #(.INIT(8'hE8)) lut_n2245 (.I0(n2225), .I1(n2243), .I2(n2244), .O(n2245));
  LUT3 #(.INIT(8'h96)) lut_n2246 (.I0(x498), .I1(x499), .I2(x500), .O(n2246));
  LUT5 #(.INIT(32'h96696996)) lut_n2247 (.I0(x489), .I1(x490), .I2(x491), .I3(n2237), .I4(n2238), .O(n2247));
  LUT5 #(.INIT(32'hFF969600)) lut_n2248 (.I0(x495), .I1(x496), .I2(x497), .I3(n2246), .I4(n2247), .O(n2248));
  LUT3 #(.INIT(8'h96)) lut_n2249 (.I0(x504), .I1(x505), .I2(x506), .O(n2249));
  LUT5 #(.INIT(32'h96696996)) lut_n2250 (.I0(x495), .I1(x496), .I2(x497), .I3(n2246), .I4(n2247), .O(n2250));
  LUT5 #(.INIT(32'hFF969600)) lut_n2251 (.I0(x501), .I1(x502), .I2(x503), .I3(n2249), .I4(n2250), .O(n2251));
  LUT3 #(.INIT(8'h96)) lut_n2252 (.I0(n2236), .I1(n2239), .I2(n2240), .O(n2252));
  LUT3 #(.INIT(8'hE8)) lut_n2253 (.I0(n2248), .I1(n2251), .I2(n2252), .O(n2253));
  LUT3 #(.INIT(8'h96)) lut_n2254 (.I0(x510), .I1(x511), .I2(x512), .O(n2254));
  LUT5 #(.INIT(32'h96696996)) lut_n2255 (.I0(x501), .I1(x502), .I2(x503), .I3(n2249), .I4(n2250), .O(n2255));
  LUT5 #(.INIT(32'hFF969600)) lut_n2256 (.I0(x507), .I1(x508), .I2(x509), .I3(n2254), .I4(n2255), .O(n2256));
  LUT3 #(.INIT(8'h96)) lut_n2257 (.I0(x516), .I1(x517), .I2(x518), .O(n2257));
  LUT5 #(.INIT(32'h96696996)) lut_n2258 (.I0(x507), .I1(x508), .I2(x509), .I3(n2254), .I4(n2255), .O(n2258));
  LUT5 #(.INIT(32'hFF969600)) lut_n2259 (.I0(x513), .I1(x514), .I2(x515), .I3(n2257), .I4(n2258), .O(n2259));
  LUT3 #(.INIT(8'h96)) lut_n2260 (.I0(n2248), .I1(n2251), .I2(n2252), .O(n2260));
  LUT3 #(.INIT(8'hE8)) lut_n2261 (.I0(n2256), .I1(n2259), .I2(n2260), .O(n2261));
  LUT3 #(.INIT(8'h96)) lut_n2262 (.I0(n2233), .I1(n2241), .I2(n2242), .O(n2262));
  LUT3 #(.INIT(8'h8E)) lut_n2263 (.I0(n2253), .I1(n2261), .I2(n2262), .O(n2263));
  LUT3 #(.INIT(8'h96)) lut_n2264 (.I0(x522), .I1(x523), .I2(x524), .O(n2264));
  LUT5 #(.INIT(32'h96696996)) lut_n2265 (.I0(x513), .I1(x514), .I2(x515), .I3(n2257), .I4(n2258), .O(n2265));
  LUT5 #(.INIT(32'hFF969600)) lut_n2266 (.I0(x519), .I1(x520), .I2(x521), .I3(n2264), .I4(n2265), .O(n2266));
  LUT3 #(.INIT(8'h96)) lut_n2267 (.I0(x528), .I1(x529), .I2(x530), .O(n2267));
  LUT5 #(.INIT(32'h96696996)) lut_n2268 (.I0(x519), .I1(x520), .I2(x521), .I3(n2264), .I4(n2265), .O(n2268));
  LUT5 #(.INIT(32'hFF969600)) lut_n2269 (.I0(x525), .I1(x526), .I2(x527), .I3(n2267), .I4(n2268), .O(n2269));
  LUT3 #(.INIT(8'h96)) lut_n2270 (.I0(n2256), .I1(n2259), .I2(n2260), .O(n2270));
  LUT3 #(.INIT(8'hE8)) lut_n2271 (.I0(n2266), .I1(n2269), .I2(n2270), .O(n2271));
  LUT3 #(.INIT(8'h96)) lut_n2272 (.I0(x534), .I1(x535), .I2(x536), .O(n2272));
  LUT5 #(.INIT(32'h96696996)) lut_n2273 (.I0(x525), .I1(x526), .I2(x527), .I3(n2267), .I4(n2268), .O(n2273));
  LUT5 #(.INIT(32'hFF969600)) lut_n2274 (.I0(x531), .I1(x532), .I2(x533), .I3(n2272), .I4(n2273), .O(n2274));
  LUT3 #(.INIT(8'h96)) lut_n2275 (.I0(x540), .I1(x541), .I2(x542), .O(n2275));
  LUT5 #(.INIT(32'h96696996)) lut_n2276 (.I0(x531), .I1(x532), .I2(x533), .I3(n2272), .I4(n2273), .O(n2276));
  LUT5 #(.INIT(32'hFF969600)) lut_n2277 (.I0(x537), .I1(x538), .I2(x539), .I3(n2275), .I4(n2276), .O(n2277));
  LUT3 #(.INIT(8'h96)) lut_n2278 (.I0(n2266), .I1(n2269), .I2(n2270), .O(n2278));
  LUT3 #(.INIT(8'hE8)) lut_n2279 (.I0(n2274), .I1(n2277), .I2(n2278), .O(n2279));
  LUT3 #(.INIT(8'h96)) lut_n2280 (.I0(n2253), .I1(n2261), .I2(n2262), .O(n2280));
  LUT3 #(.INIT(8'h8E)) lut_n2281 (.I0(n2271), .I1(n2279), .I2(n2280), .O(n2281));
  LUT3 #(.INIT(8'h96)) lut_n2282 (.I0(n2225), .I1(n2243), .I2(n2244), .O(n2282));
  LUT3 #(.INIT(8'hE8)) lut_n2283 (.I0(n2263), .I1(n2281), .I2(n2282), .O(n2283));
  LUT3 #(.INIT(8'h96)) lut_n2284 (.I0(n2165), .I1(n2203), .I2(n2204), .O(n2284));
  LUT3 #(.INIT(8'hE8)) lut_n2285 (.I0(n2245), .I1(n2283), .I2(n2284), .O(n2285));
  LUT3 #(.INIT(8'h96)) lut_n2286 (.I0(x546), .I1(x547), .I2(x548), .O(n2286));
  LUT5 #(.INIT(32'h96696996)) lut_n2287 (.I0(x537), .I1(x538), .I2(x539), .I3(n2275), .I4(n2276), .O(n2287));
  LUT5 #(.INIT(32'hFF969600)) lut_n2288 (.I0(x543), .I1(x544), .I2(x545), .I3(n2286), .I4(n2287), .O(n2288));
  LUT3 #(.INIT(8'h96)) lut_n2289 (.I0(x552), .I1(x553), .I2(x554), .O(n2289));
  LUT5 #(.INIT(32'h96696996)) lut_n2290 (.I0(x543), .I1(x544), .I2(x545), .I3(n2286), .I4(n2287), .O(n2290));
  LUT5 #(.INIT(32'hFF969600)) lut_n2291 (.I0(x549), .I1(x550), .I2(x551), .I3(n2289), .I4(n2290), .O(n2291));
  LUT3 #(.INIT(8'h96)) lut_n2292 (.I0(n2274), .I1(n2277), .I2(n2278), .O(n2292));
  LUT3 #(.INIT(8'hE8)) lut_n2293 (.I0(n2288), .I1(n2291), .I2(n2292), .O(n2293));
  LUT3 #(.INIT(8'h96)) lut_n2294 (.I0(x558), .I1(x559), .I2(x560), .O(n2294));
  LUT5 #(.INIT(32'h96696996)) lut_n2295 (.I0(x549), .I1(x550), .I2(x551), .I3(n2289), .I4(n2290), .O(n2295));
  LUT5 #(.INIT(32'hFF969600)) lut_n2296 (.I0(x555), .I1(x556), .I2(x557), .I3(n2294), .I4(n2295), .O(n2296));
  LUT3 #(.INIT(8'h96)) lut_n2297 (.I0(x564), .I1(x565), .I2(x566), .O(n2297));
  LUT5 #(.INIT(32'h96696996)) lut_n2298 (.I0(x555), .I1(x556), .I2(x557), .I3(n2294), .I4(n2295), .O(n2298));
  LUT5 #(.INIT(32'hFF969600)) lut_n2299 (.I0(x561), .I1(x562), .I2(x563), .I3(n2297), .I4(n2298), .O(n2299));
  LUT3 #(.INIT(8'h96)) lut_n2300 (.I0(n2288), .I1(n2291), .I2(n2292), .O(n2300));
  LUT3 #(.INIT(8'hE8)) lut_n2301 (.I0(n2296), .I1(n2299), .I2(n2300), .O(n2301));
  LUT3 #(.INIT(8'h96)) lut_n2302 (.I0(n2271), .I1(n2279), .I2(n2280), .O(n2302));
  LUT3 #(.INIT(8'h8E)) lut_n2303 (.I0(n2293), .I1(n2301), .I2(n2302), .O(n2303));
  LUT3 #(.INIT(8'h96)) lut_n2304 (.I0(x570), .I1(x571), .I2(x572), .O(n2304));
  LUT5 #(.INIT(32'h96696996)) lut_n2305 (.I0(x561), .I1(x562), .I2(x563), .I3(n2297), .I4(n2298), .O(n2305));
  LUT5 #(.INIT(32'hFF969600)) lut_n2306 (.I0(x567), .I1(x568), .I2(x569), .I3(n2304), .I4(n2305), .O(n2306));
  LUT3 #(.INIT(8'h96)) lut_n2307 (.I0(x576), .I1(x577), .I2(x578), .O(n2307));
  LUT5 #(.INIT(32'h96696996)) lut_n2308 (.I0(x567), .I1(x568), .I2(x569), .I3(n2304), .I4(n2305), .O(n2308));
  LUT5 #(.INIT(32'hFF969600)) lut_n2309 (.I0(x573), .I1(x574), .I2(x575), .I3(n2307), .I4(n2308), .O(n2309));
  LUT3 #(.INIT(8'h96)) lut_n2310 (.I0(n2296), .I1(n2299), .I2(n2300), .O(n2310));
  LUT3 #(.INIT(8'hE8)) lut_n2311 (.I0(n2306), .I1(n2309), .I2(n2310), .O(n2311));
  LUT3 #(.INIT(8'h96)) lut_n2312 (.I0(x582), .I1(x583), .I2(x584), .O(n2312));
  LUT5 #(.INIT(32'h96696996)) lut_n2313 (.I0(x573), .I1(x574), .I2(x575), .I3(n2307), .I4(n2308), .O(n2313));
  LUT5 #(.INIT(32'hFF969600)) lut_n2314 (.I0(x579), .I1(x580), .I2(x581), .I3(n2312), .I4(n2313), .O(n2314));
  LUT3 #(.INIT(8'h96)) lut_n2315 (.I0(x588), .I1(x589), .I2(x590), .O(n2315));
  LUT5 #(.INIT(32'h96696996)) lut_n2316 (.I0(x579), .I1(x580), .I2(x581), .I3(n2312), .I4(n2313), .O(n2316));
  LUT5 #(.INIT(32'hFF969600)) lut_n2317 (.I0(x585), .I1(x586), .I2(x587), .I3(n2315), .I4(n2316), .O(n2317));
  LUT3 #(.INIT(8'h96)) lut_n2318 (.I0(n2306), .I1(n2309), .I2(n2310), .O(n2318));
  LUT3 #(.INIT(8'hE8)) lut_n2319 (.I0(n2314), .I1(n2317), .I2(n2318), .O(n2319));
  LUT3 #(.INIT(8'h96)) lut_n2320 (.I0(n2293), .I1(n2301), .I2(n2302), .O(n2320));
  LUT3 #(.INIT(8'h8E)) lut_n2321 (.I0(n2311), .I1(n2319), .I2(n2320), .O(n2321));
  LUT3 #(.INIT(8'h96)) lut_n2322 (.I0(n2263), .I1(n2281), .I2(n2282), .O(n2322));
  LUT3 #(.INIT(8'hE8)) lut_n2323 (.I0(n2303), .I1(n2321), .I2(n2322), .O(n2323));
  LUT3 #(.INIT(8'h96)) lut_n2324 (.I0(x594), .I1(x595), .I2(x596), .O(n2324));
  LUT5 #(.INIT(32'h96696996)) lut_n2325 (.I0(x585), .I1(x586), .I2(x587), .I3(n2315), .I4(n2316), .O(n2325));
  LUT5 #(.INIT(32'hFF969600)) lut_n2326 (.I0(x591), .I1(x592), .I2(x593), .I3(n2324), .I4(n2325), .O(n2326));
  LUT3 #(.INIT(8'h96)) lut_n2327 (.I0(x600), .I1(x601), .I2(x602), .O(n2327));
  LUT5 #(.INIT(32'h96696996)) lut_n2328 (.I0(x591), .I1(x592), .I2(x593), .I3(n2324), .I4(n2325), .O(n2328));
  LUT5 #(.INIT(32'hFF969600)) lut_n2329 (.I0(x597), .I1(x598), .I2(x599), .I3(n2327), .I4(n2328), .O(n2329));
  LUT3 #(.INIT(8'h96)) lut_n2330 (.I0(n2314), .I1(n2317), .I2(n2318), .O(n2330));
  LUT3 #(.INIT(8'hE8)) lut_n2331 (.I0(n2326), .I1(n2329), .I2(n2330), .O(n2331));
  LUT3 #(.INIT(8'h96)) lut_n2332 (.I0(x606), .I1(x607), .I2(x608), .O(n2332));
  LUT5 #(.INIT(32'h96696996)) lut_n2333 (.I0(x597), .I1(x598), .I2(x599), .I3(n2327), .I4(n2328), .O(n2333));
  LUT5 #(.INIT(32'hFF969600)) lut_n2334 (.I0(x603), .I1(x604), .I2(x605), .I3(n2332), .I4(n2333), .O(n2334));
  LUT3 #(.INIT(8'h96)) lut_n2335 (.I0(x612), .I1(x613), .I2(x614), .O(n2335));
  LUT5 #(.INIT(32'h96696996)) lut_n2336 (.I0(x603), .I1(x604), .I2(x605), .I3(n2332), .I4(n2333), .O(n2336));
  LUT5 #(.INIT(32'hFF969600)) lut_n2337 (.I0(x609), .I1(x610), .I2(x611), .I3(n2335), .I4(n2336), .O(n2337));
  LUT3 #(.INIT(8'h96)) lut_n2338 (.I0(n2326), .I1(n2329), .I2(n2330), .O(n2338));
  LUT3 #(.INIT(8'hE8)) lut_n2339 (.I0(n2334), .I1(n2337), .I2(n2338), .O(n2339));
  LUT3 #(.INIT(8'h96)) lut_n2340 (.I0(n2311), .I1(n2319), .I2(n2320), .O(n2340));
  LUT3 #(.INIT(8'h8E)) lut_n2341 (.I0(n2331), .I1(n2339), .I2(n2340), .O(n2341));
  LUT3 #(.INIT(8'h96)) lut_n2342 (.I0(x618), .I1(x619), .I2(x620), .O(n2342));
  LUT5 #(.INIT(32'h96696996)) lut_n2343 (.I0(x609), .I1(x610), .I2(x611), .I3(n2335), .I4(n2336), .O(n2343));
  LUT5 #(.INIT(32'hFF969600)) lut_n2344 (.I0(x615), .I1(x616), .I2(x617), .I3(n2342), .I4(n2343), .O(n2344));
  LUT3 #(.INIT(8'h96)) lut_n2345 (.I0(x624), .I1(x625), .I2(x626), .O(n2345));
  LUT5 #(.INIT(32'h96696996)) lut_n2346 (.I0(x615), .I1(x616), .I2(x617), .I3(n2342), .I4(n2343), .O(n2346));
  LUT5 #(.INIT(32'hFF969600)) lut_n2347 (.I0(x621), .I1(x622), .I2(x623), .I3(n2345), .I4(n2346), .O(n2347));
  LUT3 #(.INIT(8'h96)) lut_n2348 (.I0(n2334), .I1(n2337), .I2(n2338), .O(n2348));
  LUT3 #(.INIT(8'hE8)) lut_n2349 (.I0(n2344), .I1(n2347), .I2(n2348), .O(n2349));
  LUT3 #(.INIT(8'h96)) lut_n2350 (.I0(x630), .I1(x631), .I2(x632), .O(n2350));
  LUT5 #(.INIT(32'h96696996)) lut_n2351 (.I0(x621), .I1(x622), .I2(x623), .I3(n2345), .I4(n2346), .O(n2351));
  LUT5 #(.INIT(32'hFF969600)) lut_n2352 (.I0(x627), .I1(x628), .I2(x629), .I3(n2350), .I4(n2351), .O(n2352));
  LUT3 #(.INIT(8'h96)) lut_n2353 (.I0(x636), .I1(x637), .I2(x638), .O(n2353));
  LUT5 #(.INIT(32'h96696996)) lut_n2354 (.I0(x627), .I1(x628), .I2(x629), .I3(n2350), .I4(n2351), .O(n2354));
  LUT5 #(.INIT(32'hFF969600)) lut_n2355 (.I0(x633), .I1(x634), .I2(x635), .I3(n2353), .I4(n2354), .O(n2355));
  LUT3 #(.INIT(8'h96)) lut_n2356 (.I0(n2344), .I1(n2347), .I2(n2348), .O(n2356));
  LUT3 #(.INIT(8'hE8)) lut_n2357 (.I0(n2352), .I1(n2355), .I2(n2356), .O(n2357));
  LUT3 #(.INIT(8'h96)) lut_n2358 (.I0(n2331), .I1(n2339), .I2(n2340), .O(n2358));
  LUT3 #(.INIT(8'h8E)) lut_n2359 (.I0(n2349), .I1(n2357), .I2(n2358), .O(n2359));
  LUT3 #(.INIT(8'h96)) lut_n2360 (.I0(n2303), .I1(n2321), .I2(n2322), .O(n2360));
  LUT3 #(.INIT(8'hE8)) lut_n2361 (.I0(n2341), .I1(n2359), .I2(n2360), .O(n2361));
  LUT3 #(.INIT(8'h96)) lut_n2362 (.I0(n2245), .I1(n2283), .I2(n2284), .O(n2362));
  LUT3 #(.INIT(8'hE8)) lut_n2363 (.I0(n2323), .I1(n2361), .I2(n2362), .O(n2363));
  LUT3 #(.INIT(8'h96)) lut_n2364 (.I0(n2127), .I1(n2205), .I2(n2206), .O(n2364));
  LUT3 #(.INIT(8'hE8)) lut_n2365 (.I0(n2285), .I1(n2363), .I2(n2364), .O(n2365));
  LUT3 #(.INIT(8'h96)) lut_n2366 (.I0(n1887), .I1(n2045), .I2(n2046), .O(n2366));
  LUT3 #(.INIT(8'hE8)) lut_n2367 (.I0(n2207), .I1(n2365), .I2(n2366), .O(n2367));
  LUT3 #(.INIT(8'h96)) lut_n2368 (.I0(x642), .I1(x643), .I2(x644), .O(n2368));
  LUT5 #(.INIT(32'h96696996)) lut_n2369 (.I0(x633), .I1(x634), .I2(x635), .I3(n2353), .I4(n2354), .O(n2369));
  LUT5 #(.INIT(32'hFF969600)) lut_n2370 (.I0(x639), .I1(x640), .I2(x641), .I3(n2368), .I4(n2369), .O(n2370));
  LUT3 #(.INIT(8'h96)) lut_n2371 (.I0(x648), .I1(x649), .I2(x650), .O(n2371));
  LUT5 #(.INIT(32'h96696996)) lut_n2372 (.I0(x639), .I1(x640), .I2(x641), .I3(n2368), .I4(n2369), .O(n2372));
  LUT5 #(.INIT(32'hFF969600)) lut_n2373 (.I0(x645), .I1(x646), .I2(x647), .I3(n2371), .I4(n2372), .O(n2373));
  LUT3 #(.INIT(8'h96)) lut_n2374 (.I0(n2352), .I1(n2355), .I2(n2356), .O(n2374));
  LUT3 #(.INIT(8'hE8)) lut_n2375 (.I0(n2370), .I1(n2373), .I2(n2374), .O(n2375));
  LUT3 #(.INIT(8'h96)) lut_n2376 (.I0(x654), .I1(x655), .I2(x656), .O(n2376));
  LUT5 #(.INIT(32'h96696996)) lut_n2377 (.I0(x645), .I1(x646), .I2(x647), .I3(n2371), .I4(n2372), .O(n2377));
  LUT5 #(.INIT(32'hFF969600)) lut_n2378 (.I0(x651), .I1(x652), .I2(x653), .I3(n2376), .I4(n2377), .O(n2378));
  LUT3 #(.INIT(8'h96)) lut_n2379 (.I0(x660), .I1(x661), .I2(x662), .O(n2379));
  LUT5 #(.INIT(32'h96696996)) lut_n2380 (.I0(x651), .I1(x652), .I2(x653), .I3(n2376), .I4(n2377), .O(n2380));
  LUT5 #(.INIT(32'hFF969600)) lut_n2381 (.I0(x657), .I1(x658), .I2(x659), .I3(n2379), .I4(n2380), .O(n2381));
  LUT3 #(.INIT(8'h96)) lut_n2382 (.I0(n2370), .I1(n2373), .I2(n2374), .O(n2382));
  LUT3 #(.INIT(8'hE8)) lut_n2383 (.I0(n2378), .I1(n2381), .I2(n2382), .O(n2383));
  LUT3 #(.INIT(8'h96)) lut_n2384 (.I0(n2349), .I1(n2357), .I2(n2358), .O(n2384));
  LUT3 #(.INIT(8'h8E)) lut_n2385 (.I0(n2375), .I1(n2383), .I2(n2384), .O(n2385));
  LUT3 #(.INIT(8'h96)) lut_n2386 (.I0(x666), .I1(x667), .I2(x668), .O(n2386));
  LUT5 #(.INIT(32'h96696996)) lut_n2387 (.I0(x657), .I1(x658), .I2(x659), .I3(n2379), .I4(n2380), .O(n2387));
  LUT5 #(.INIT(32'hFF969600)) lut_n2388 (.I0(x663), .I1(x664), .I2(x665), .I3(n2386), .I4(n2387), .O(n2388));
  LUT3 #(.INIT(8'h96)) lut_n2389 (.I0(x672), .I1(x673), .I2(x674), .O(n2389));
  LUT5 #(.INIT(32'h96696996)) lut_n2390 (.I0(x663), .I1(x664), .I2(x665), .I3(n2386), .I4(n2387), .O(n2390));
  LUT5 #(.INIT(32'hFF969600)) lut_n2391 (.I0(x669), .I1(x670), .I2(x671), .I3(n2389), .I4(n2390), .O(n2391));
  LUT3 #(.INIT(8'h96)) lut_n2392 (.I0(n2378), .I1(n2381), .I2(n2382), .O(n2392));
  LUT3 #(.INIT(8'hE8)) lut_n2393 (.I0(n2388), .I1(n2391), .I2(n2392), .O(n2393));
  LUT3 #(.INIT(8'h96)) lut_n2394 (.I0(x678), .I1(x679), .I2(x680), .O(n2394));
  LUT5 #(.INIT(32'h96696996)) lut_n2395 (.I0(x669), .I1(x670), .I2(x671), .I3(n2389), .I4(n2390), .O(n2395));
  LUT5 #(.INIT(32'hFF969600)) lut_n2396 (.I0(x675), .I1(x676), .I2(x677), .I3(n2394), .I4(n2395), .O(n2396));
  LUT3 #(.INIT(8'h96)) lut_n2397 (.I0(x684), .I1(x685), .I2(x686), .O(n2397));
  LUT5 #(.INIT(32'h96696996)) lut_n2398 (.I0(x675), .I1(x676), .I2(x677), .I3(n2394), .I4(n2395), .O(n2398));
  LUT5 #(.INIT(32'hFF969600)) lut_n2399 (.I0(x681), .I1(x682), .I2(x683), .I3(n2397), .I4(n2398), .O(n2399));
  LUT3 #(.INIT(8'h96)) lut_n2400 (.I0(n2388), .I1(n2391), .I2(n2392), .O(n2400));
  LUT3 #(.INIT(8'hE8)) lut_n2401 (.I0(n2396), .I1(n2399), .I2(n2400), .O(n2401));
  LUT3 #(.INIT(8'h96)) lut_n2402 (.I0(n2375), .I1(n2383), .I2(n2384), .O(n2402));
  LUT3 #(.INIT(8'h8E)) lut_n2403 (.I0(n2393), .I1(n2401), .I2(n2402), .O(n2403));
  LUT3 #(.INIT(8'h96)) lut_n2404 (.I0(n2341), .I1(n2359), .I2(n2360), .O(n2404));
  LUT3 #(.INIT(8'hE8)) lut_n2405 (.I0(n2385), .I1(n2403), .I2(n2404), .O(n2405));
  LUT3 #(.INIT(8'h96)) lut_n2406 (.I0(x690), .I1(x691), .I2(x692), .O(n2406));
  LUT5 #(.INIT(32'h96696996)) lut_n2407 (.I0(x681), .I1(x682), .I2(x683), .I3(n2397), .I4(n2398), .O(n2407));
  LUT5 #(.INIT(32'hFF969600)) lut_n2408 (.I0(x687), .I1(x688), .I2(x689), .I3(n2406), .I4(n2407), .O(n2408));
  LUT3 #(.INIT(8'h96)) lut_n2409 (.I0(x696), .I1(x697), .I2(x698), .O(n2409));
  LUT5 #(.INIT(32'h96696996)) lut_n2410 (.I0(x687), .I1(x688), .I2(x689), .I3(n2406), .I4(n2407), .O(n2410));
  LUT5 #(.INIT(32'hFF969600)) lut_n2411 (.I0(x693), .I1(x694), .I2(x695), .I3(n2409), .I4(n2410), .O(n2411));
  LUT3 #(.INIT(8'h96)) lut_n2412 (.I0(n2396), .I1(n2399), .I2(n2400), .O(n2412));
  LUT3 #(.INIT(8'hE8)) lut_n2413 (.I0(n2408), .I1(n2411), .I2(n2412), .O(n2413));
  LUT3 #(.INIT(8'h96)) lut_n2414 (.I0(x702), .I1(x703), .I2(x704), .O(n2414));
  LUT5 #(.INIT(32'h96696996)) lut_n2415 (.I0(x693), .I1(x694), .I2(x695), .I3(n2409), .I4(n2410), .O(n2415));
  LUT5 #(.INIT(32'hFF969600)) lut_n2416 (.I0(x699), .I1(x700), .I2(x701), .I3(n2414), .I4(n2415), .O(n2416));
  LUT3 #(.INIT(8'h96)) lut_n2417 (.I0(x708), .I1(x709), .I2(x710), .O(n2417));
  LUT5 #(.INIT(32'h96696996)) lut_n2418 (.I0(x699), .I1(x700), .I2(x701), .I3(n2414), .I4(n2415), .O(n2418));
  LUT5 #(.INIT(32'hFF969600)) lut_n2419 (.I0(x705), .I1(x706), .I2(x707), .I3(n2417), .I4(n2418), .O(n2419));
  LUT3 #(.INIT(8'h96)) lut_n2420 (.I0(n2408), .I1(n2411), .I2(n2412), .O(n2420));
  LUT3 #(.INIT(8'hE8)) lut_n2421 (.I0(n2416), .I1(n2419), .I2(n2420), .O(n2421));
  LUT3 #(.INIT(8'h96)) lut_n2422 (.I0(n2393), .I1(n2401), .I2(n2402), .O(n2422));
  LUT3 #(.INIT(8'h8E)) lut_n2423 (.I0(n2413), .I1(n2421), .I2(n2422), .O(n2423));
  LUT3 #(.INIT(8'h96)) lut_n2424 (.I0(x714), .I1(x715), .I2(x716), .O(n2424));
  LUT5 #(.INIT(32'h96696996)) lut_n2425 (.I0(x705), .I1(x706), .I2(x707), .I3(n2417), .I4(n2418), .O(n2425));
  LUT5 #(.INIT(32'hFF969600)) lut_n2426 (.I0(x711), .I1(x712), .I2(x713), .I3(n2424), .I4(n2425), .O(n2426));
  LUT3 #(.INIT(8'h96)) lut_n2427 (.I0(x720), .I1(x721), .I2(x722), .O(n2427));
  LUT5 #(.INIT(32'h96696996)) lut_n2428 (.I0(x711), .I1(x712), .I2(x713), .I3(n2424), .I4(n2425), .O(n2428));
  LUT5 #(.INIT(32'hFF969600)) lut_n2429 (.I0(x717), .I1(x718), .I2(x719), .I3(n2427), .I4(n2428), .O(n2429));
  LUT3 #(.INIT(8'h96)) lut_n2430 (.I0(n2416), .I1(n2419), .I2(n2420), .O(n2430));
  LUT3 #(.INIT(8'hE8)) lut_n2431 (.I0(n2426), .I1(n2429), .I2(n2430), .O(n2431));
  LUT3 #(.INIT(8'h96)) lut_n2432 (.I0(x726), .I1(x727), .I2(x728), .O(n2432));
  LUT5 #(.INIT(32'h96696996)) lut_n2433 (.I0(x717), .I1(x718), .I2(x719), .I3(n2427), .I4(n2428), .O(n2433));
  LUT5 #(.INIT(32'hFF969600)) lut_n2434 (.I0(x723), .I1(x724), .I2(x725), .I3(n2432), .I4(n2433), .O(n2434));
  LUT3 #(.INIT(8'h96)) lut_n2435 (.I0(x732), .I1(x733), .I2(x734), .O(n2435));
  LUT5 #(.INIT(32'h96696996)) lut_n2436 (.I0(x723), .I1(x724), .I2(x725), .I3(n2432), .I4(n2433), .O(n2436));
  LUT5 #(.INIT(32'hFF969600)) lut_n2437 (.I0(x729), .I1(x730), .I2(x731), .I3(n2435), .I4(n2436), .O(n2437));
  LUT3 #(.INIT(8'h96)) lut_n2438 (.I0(n2426), .I1(n2429), .I2(n2430), .O(n2438));
  LUT3 #(.INIT(8'hE8)) lut_n2439 (.I0(n2434), .I1(n2437), .I2(n2438), .O(n2439));
  LUT3 #(.INIT(8'h96)) lut_n2440 (.I0(n2413), .I1(n2421), .I2(n2422), .O(n2440));
  LUT3 #(.INIT(8'h8E)) lut_n2441 (.I0(n2431), .I1(n2439), .I2(n2440), .O(n2441));
  LUT3 #(.INIT(8'h96)) lut_n2442 (.I0(n2385), .I1(n2403), .I2(n2404), .O(n2442));
  LUT3 #(.INIT(8'hE8)) lut_n2443 (.I0(n2423), .I1(n2441), .I2(n2442), .O(n2443));
  LUT3 #(.INIT(8'h96)) lut_n2444 (.I0(n2323), .I1(n2361), .I2(n2362), .O(n2444));
  LUT3 #(.INIT(8'hE8)) lut_n2445 (.I0(n2405), .I1(n2443), .I2(n2444), .O(n2445));
  LUT3 #(.INIT(8'h96)) lut_n2446 (.I0(x738), .I1(x739), .I2(x740), .O(n2446));
  LUT5 #(.INIT(32'h96696996)) lut_n2447 (.I0(x729), .I1(x730), .I2(x731), .I3(n2435), .I4(n2436), .O(n2447));
  LUT5 #(.INIT(32'hFF969600)) lut_n2448 (.I0(x735), .I1(x736), .I2(x737), .I3(n2446), .I4(n2447), .O(n2448));
  LUT3 #(.INIT(8'h96)) lut_n2449 (.I0(x744), .I1(x745), .I2(x746), .O(n2449));
  LUT5 #(.INIT(32'h96696996)) lut_n2450 (.I0(x735), .I1(x736), .I2(x737), .I3(n2446), .I4(n2447), .O(n2450));
  LUT5 #(.INIT(32'hFF969600)) lut_n2451 (.I0(x741), .I1(x742), .I2(x743), .I3(n2449), .I4(n2450), .O(n2451));
  LUT3 #(.INIT(8'h96)) lut_n2452 (.I0(n2434), .I1(n2437), .I2(n2438), .O(n2452));
  LUT3 #(.INIT(8'hE8)) lut_n2453 (.I0(n2448), .I1(n2451), .I2(n2452), .O(n2453));
  LUT3 #(.INIT(8'h96)) lut_n2454 (.I0(x750), .I1(x751), .I2(x752), .O(n2454));
  LUT5 #(.INIT(32'h96696996)) lut_n2455 (.I0(x741), .I1(x742), .I2(x743), .I3(n2449), .I4(n2450), .O(n2455));
  LUT5 #(.INIT(32'hFF969600)) lut_n2456 (.I0(x747), .I1(x748), .I2(x749), .I3(n2454), .I4(n2455), .O(n2456));
  LUT3 #(.INIT(8'h96)) lut_n2457 (.I0(x756), .I1(x757), .I2(x758), .O(n2457));
  LUT5 #(.INIT(32'h96696996)) lut_n2458 (.I0(x747), .I1(x748), .I2(x749), .I3(n2454), .I4(n2455), .O(n2458));
  LUT5 #(.INIT(32'hFF969600)) lut_n2459 (.I0(x753), .I1(x754), .I2(x755), .I3(n2457), .I4(n2458), .O(n2459));
  LUT3 #(.INIT(8'h96)) lut_n2460 (.I0(n2448), .I1(n2451), .I2(n2452), .O(n2460));
  LUT3 #(.INIT(8'hE8)) lut_n2461 (.I0(n2456), .I1(n2459), .I2(n2460), .O(n2461));
  LUT3 #(.INIT(8'h96)) lut_n2462 (.I0(n2431), .I1(n2439), .I2(n2440), .O(n2462));
  LUT3 #(.INIT(8'h8E)) lut_n2463 (.I0(n2453), .I1(n2461), .I2(n2462), .O(n2463));
  LUT3 #(.INIT(8'h96)) lut_n2464 (.I0(x762), .I1(x763), .I2(x764), .O(n2464));
  LUT5 #(.INIT(32'h96696996)) lut_n2465 (.I0(x753), .I1(x754), .I2(x755), .I3(n2457), .I4(n2458), .O(n2465));
  LUT5 #(.INIT(32'hFF969600)) lut_n2466 (.I0(x759), .I1(x760), .I2(x761), .I3(n2464), .I4(n2465), .O(n2466));
  LUT3 #(.INIT(8'h96)) lut_n2467 (.I0(x768), .I1(x769), .I2(x770), .O(n2467));
  LUT5 #(.INIT(32'h96696996)) lut_n2468 (.I0(x759), .I1(x760), .I2(x761), .I3(n2464), .I4(n2465), .O(n2468));
  LUT5 #(.INIT(32'hFF969600)) lut_n2469 (.I0(x765), .I1(x766), .I2(x767), .I3(n2467), .I4(n2468), .O(n2469));
  LUT3 #(.INIT(8'h96)) lut_n2470 (.I0(n2456), .I1(n2459), .I2(n2460), .O(n2470));
  LUT3 #(.INIT(8'hE8)) lut_n2471 (.I0(n2466), .I1(n2469), .I2(n2470), .O(n2471));
  LUT3 #(.INIT(8'h96)) lut_n2472 (.I0(x774), .I1(x775), .I2(x776), .O(n2472));
  LUT5 #(.INIT(32'h96696996)) lut_n2473 (.I0(x765), .I1(x766), .I2(x767), .I3(n2467), .I4(n2468), .O(n2473));
  LUT5 #(.INIT(32'hFF969600)) lut_n2474 (.I0(x771), .I1(x772), .I2(x773), .I3(n2472), .I4(n2473), .O(n2474));
  LUT3 #(.INIT(8'h96)) lut_n2475 (.I0(x780), .I1(x781), .I2(x782), .O(n2475));
  LUT5 #(.INIT(32'h96696996)) lut_n2476 (.I0(x771), .I1(x772), .I2(x773), .I3(n2472), .I4(n2473), .O(n2476));
  LUT5 #(.INIT(32'hFF969600)) lut_n2477 (.I0(x777), .I1(x778), .I2(x779), .I3(n2475), .I4(n2476), .O(n2477));
  LUT3 #(.INIT(8'h96)) lut_n2478 (.I0(n2466), .I1(n2469), .I2(n2470), .O(n2478));
  LUT3 #(.INIT(8'hE8)) lut_n2479 (.I0(n2474), .I1(n2477), .I2(n2478), .O(n2479));
  LUT3 #(.INIT(8'h96)) lut_n2480 (.I0(n2453), .I1(n2461), .I2(n2462), .O(n2480));
  LUT3 #(.INIT(8'h8E)) lut_n2481 (.I0(n2471), .I1(n2479), .I2(n2480), .O(n2481));
  LUT3 #(.INIT(8'h96)) lut_n2482 (.I0(n2423), .I1(n2441), .I2(n2442), .O(n2482));
  LUT3 #(.INIT(8'hE8)) lut_n2483 (.I0(n2463), .I1(n2481), .I2(n2482), .O(n2483));
  LUT3 #(.INIT(8'h96)) lut_n2484 (.I0(x786), .I1(x787), .I2(x788), .O(n2484));
  LUT5 #(.INIT(32'h96696996)) lut_n2485 (.I0(x777), .I1(x778), .I2(x779), .I3(n2475), .I4(n2476), .O(n2485));
  LUT5 #(.INIT(32'hFF969600)) lut_n2486 (.I0(x783), .I1(x784), .I2(x785), .I3(n2484), .I4(n2485), .O(n2486));
  LUT3 #(.INIT(8'h96)) lut_n2487 (.I0(x792), .I1(x793), .I2(x794), .O(n2487));
  LUT5 #(.INIT(32'h96696996)) lut_n2488 (.I0(x783), .I1(x784), .I2(x785), .I3(n2484), .I4(n2485), .O(n2488));
  LUT5 #(.INIT(32'hFF969600)) lut_n2489 (.I0(x789), .I1(x790), .I2(x791), .I3(n2487), .I4(n2488), .O(n2489));
  LUT3 #(.INIT(8'h96)) lut_n2490 (.I0(n2474), .I1(n2477), .I2(n2478), .O(n2490));
  LUT3 #(.INIT(8'hE8)) lut_n2491 (.I0(n2486), .I1(n2489), .I2(n2490), .O(n2491));
  LUT3 #(.INIT(8'h96)) lut_n2492 (.I0(x798), .I1(x799), .I2(x800), .O(n2492));
  LUT5 #(.INIT(32'h96696996)) lut_n2493 (.I0(x789), .I1(x790), .I2(x791), .I3(n2487), .I4(n2488), .O(n2493));
  LUT5 #(.INIT(32'hFF969600)) lut_n2494 (.I0(x795), .I1(x796), .I2(x797), .I3(n2492), .I4(n2493), .O(n2494));
  LUT3 #(.INIT(8'h96)) lut_n2495 (.I0(x804), .I1(x805), .I2(x806), .O(n2495));
  LUT5 #(.INIT(32'h96696996)) lut_n2496 (.I0(x795), .I1(x796), .I2(x797), .I3(n2492), .I4(n2493), .O(n2496));
  LUT5 #(.INIT(32'hFF969600)) lut_n2497 (.I0(x801), .I1(x802), .I2(x803), .I3(n2495), .I4(n2496), .O(n2497));
  LUT3 #(.INIT(8'h96)) lut_n2498 (.I0(n2486), .I1(n2489), .I2(n2490), .O(n2498));
  LUT3 #(.INIT(8'hE8)) lut_n2499 (.I0(n2494), .I1(n2497), .I2(n2498), .O(n2499));
  LUT3 #(.INIT(8'h96)) lut_n2500 (.I0(n2471), .I1(n2479), .I2(n2480), .O(n2500));
  LUT3 #(.INIT(8'h8E)) lut_n2501 (.I0(n2491), .I1(n2499), .I2(n2500), .O(n2501));
  LUT3 #(.INIT(8'h96)) lut_n2502 (.I0(x810), .I1(x811), .I2(x812), .O(n2502));
  LUT5 #(.INIT(32'h96696996)) lut_n2503 (.I0(x801), .I1(x802), .I2(x803), .I3(n2495), .I4(n2496), .O(n2503));
  LUT5 #(.INIT(32'hFF969600)) lut_n2504 (.I0(x807), .I1(x808), .I2(x809), .I3(n2502), .I4(n2503), .O(n2504));
  LUT3 #(.INIT(8'h96)) lut_n2505 (.I0(x816), .I1(x817), .I2(x818), .O(n2505));
  LUT5 #(.INIT(32'h96696996)) lut_n2506 (.I0(x807), .I1(x808), .I2(x809), .I3(n2502), .I4(n2503), .O(n2506));
  LUT5 #(.INIT(32'hFF969600)) lut_n2507 (.I0(x813), .I1(x814), .I2(x815), .I3(n2505), .I4(n2506), .O(n2507));
  LUT3 #(.INIT(8'h96)) lut_n2508 (.I0(n2494), .I1(n2497), .I2(n2498), .O(n2508));
  LUT3 #(.INIT(8'hE8)) lut_n2509 (.I0(n2504), .I1(n2507), .I2(n2508), .O(n2509));
  LUT3 #(.INIT(8'h96)) lut_n2510 (.I0(x822), .I1(x823), .I2(x824), .O(n2510));
  LUT5 #(.INIT(32'h96696996)) lut_n2511 (.I0(x813), .I1(x814), .I2(x815), .I3(n2505), .I4(n2506), .O(n2511));
  LUT5 #(.INIT(32'hFF969600)) lut_n2512 (.I0(x819), .I1(x820), .I2(x821), .I3(n2510), .I4(n2511), .O(n2512));
  LUT3 #(.INIT(8'h96)) lut_n2513 (.I0(x828), .I1(x829), .I2(x830), .O(n2513));
  LUT5 #(.INIT(32'h96696996)) lut_n2514 (.I0(x819), .I1(x820), .I2(x821), .I3(n2510), .I4(n2511), .O(n2514));
  LUT5 #(.INIT(32'hFF969600)) lut_n2515 (.I0(x825), .I1(x826), .I2(x827), .I3(n2513), .I4(n2514), .O(n2515));
  LUT3 #(.INIT(8'h96)) lut_n2516 (.I0(n2504), .I1(n2507), .I2(n2508), .O(n2516));
  LUT3 #(.INIT(8'hE8)) lut_n2517 (.I0(n2512), .I1(n2515), .I2(n2516), .O(n2517));
  LUT3 #(.INIT(8'h96)) lut_n2518 (.I0(n2491), .I1(n2499), .I2(n2500), .O(n2518));
  LUT3 #(.INIT(8'h8E)) lut_n2519 (.I0(n2509), .I1(n2517), .I2(n2518), .O(n2519));
  LUT3 #(.INIT(8'h96)) lut_n2520 (.I0(n2463), .I1(n2481), .I2(n2482), .O(n2520));
  LUT3 #(.INIT(8'hE8)) lut_n2521 (.I0(n2501), .I1(n2519), .I2(n2520), .O(n2521));
  LUT3 #(.INIT(8'h96)) lut_n2522 (.I0(n2405), .I1(n2443), .I2(n2444), .O(n2522));
  LUT3 #(.INIT(8'hE8)) lut_n2523 (.I0(n2483), .I1(n2521), .I2(n2522), .O(n2523));
  LUT3 #(.INIT(8'h96)) lut_n2524 (.I0(n2285), .I1(n2363), .I2(n2364), .O(n2524));
  LUT3 #(.INIT(8'h96)) lut_n2525 (.I0(x834), .I1(x835), .I2(x836), .O(n2525));
  LUT5 #(.INIT(32'h96696996)) lut_n2526 (.I0(x825), .I1(x826), .I2(x827), .I3(n2513), .I4(n2514), .O(n2526));
  LUT5 #(.INIT(32'hFF969600)) lut_n2527 (.I0(x831), .I1(x832), .I2(x833), .I3(n2525), .I4(n2526), .O(n2527));
  LUT3 #(.INIT(8'h96)) lut_n2528 (.I0(x840), .I1(x841), .I2(x842), .O(n2528));
  LUT5 #(.INIT(32'h96696996)) lut_n2529 (.I0(x831), .I1(x832), .I2(x833), .I3(n2525), .I4(n2526), .O(n2529));
  LUT5 #(.INIT(32'hFF969600)) lut_n2530 (.I0(x837), .I1(x838), .I2(x839), .I3(n2528), .I4(n2529), .O(n2530));
  LUT3 #(.INIT(8'h96)) lut_n2531 (.I0(n2512), .I1(n2515), .I2(n2516), .O(n2531));
  LUT3 #(.INIT(8'hE8)) lut_n2532 (.I0(n2527), .I1(n2530), .I2(n2531), .O(n2532));
  LUT3 #(.INIT(8'h96)) lut_n2533 (.I0(x846), .I1(x847), .I2(x848), .O(n2533));
  LUT5 #(.INIT(32'h96696996)) lut_n2534 (.I0(x837), .I1(x838), .I2(x839), .I3(n2528), .I4(n2529), .O(n2534));
  LUT5 #(.INIT(32'hFF969600)) lut_n2535 (.I0(x843), .I1(x844), .I2(x845), .I3(n2533), .I4(n2534), .O(n2535));
  LUT3 #(.INIT(8'h96)) lut_n2536 (.I0(x852), .I1(x853), .I2(x854), .O(n2536));
  LUT5 #(.INIT(32'h96696996)) lut_n2537 (.I0(x843), .I1(x844), .I2(x845), .I3(n2533), .I4(n2534), .O(n2537));
  LUT5 #(.INIT(32'hFF969600)) lut_n2538 (.I0(x849), .I1(x850), .I2(x851), .I3(n2536), .I4(n2537), .O(n2538));
  LUT3 #(.INIT(8'h96)) lut_n2539 (.I0(n2527), .I1(n2530), .I2(n2531), .O(n2539));
  LUT3 #(.INIT(8'hE8)) lut_n2540 (.I0(n2535), .I1(n2538), .I2(n2539), .O(n2540));
  LUT3 #(.INIT(8'h96)) lut_n2541 (.I0(n2509), .I1(n2517), .I2(n2518), .O(n2541));
  LUT3 #(.INIT(8'h8E)) lut_n2542 (.I0(n2532), .I1(n2540), .I2(n2541), .O(n2542));
  LUT3 #(.INIT(8'h96)) lut_n2543 (.I0(x858), .I1(x859), .I2(x860), .O(n2543));
  LUT5 #(.INIT(32'h96696996)) lut_n2544 (.I0(x849), .I1(x850), .I2(x851), .I3(n2536), .I4(n2537), .O(n2544));
  LUT5 #(.INIT(32'hFF969600)) lut_n2545 (.I0(x855), .I1(x856), .I2(x857), .I3(n2543), .I4(n2544), .O(n2545));
  LUT3 #(.INIT(8'h96)) lut_n2546 (.I0(x864), .I1(x865), .I2(x866), .O(n2546));
  LUT5 #(.INIT(32'h96696996)) lut_n2547 (.I0(x855), .I1(x856), .I2(x857), .I3(n2543), .I4(n2544), .O(n2547));
  LUT5 #(.INIT(32'hFF969600)) lut_n2548 (.I0(x861), .I1(x862), .I2(x863), .I3(n2546), .I4(n2547), .O(n2548));
  LUT3 #(.INIT(8'h96)) lut_n2549 (.I0(n2535), .I1(n2538), .I2(n2539), .O(n2549));
  LUT3 #(.INIT(8'hE8)) lut_n2550 (.I0(n2545), .I1(n2548), .I2(n2549), .O(n2550));
  LUT3 #(.INIT(8'h96)) lut_n2551 (.I0(x870), .I1(x871), .I2(x872), .O(n2551));
  LUT5 #(.INIT(32'h96696996)) lut_n2552 (.I0(x861), .I1(x862), .I2(x863), .I3(n2546), .I4(n2547), .O(n2552));
  LUT5 #(.INIT(32'hFF969600)) lut_n2553 (.I0(x867), .I1(x868), .I2(x869), .I3(n2551), .I4(n2552), .O(n2553));
  LUT3 #(.INIT(8'h96)) lut_n2554 (.I0(x876), .I1(x877), .I2(x878), .O(n2554));
  LUT5 #(.INIT(32'h96696996)) lut_n2555 (.I0(x867), .I1(x868), .I2(x869), .I3(n2551), .I4(n2552), .O(n2555));
  LUT5 #(.INIT(32'hFF969600)) lut_n2556 (.I0(x873), .I1(x874), .I2(x875), .I3(n2554), .I4(n2555), .O(n2556));
  LUT3 #(.INIT(8'h96)) lut_n2557 (.I0(n2545), .I1(n2548), .I2(n2549), .O(n2557));
  LUT3 #(.INIT(8'hE8)) lut_n2558 (.I0(n2553), .I1(n2556), .I2(n2557), .O(n2558));
  LUT3 #(.INIT(8'h96)) lut_n2559 (.I0(n2532), .I1(n2540), .I2(n2541), .O(n2559));
  LUT3 #(.INIT(8'h8E)) lut_n2560 (.I0(n2550), .I1(n2558), .I2(n2559), .O(n2560));
  LUT3 #(.INIT(8'h96)) lut_n2561 (.I0(n2501), .I1(n2519), .I2(n2520), .O(n2561));
  LUT3 #(.INIT(8'hE8)) lut_n2562 (.I0(n2542), .I1(n2560), .I2(n2561), .O(n2562));
  LUT3 #(.INIT(8'h96)) lut_n2563 (.I0(x882), .I1(x883), .I2(x884), .O(n2563));
  LUT5 #(.INIT(32'h96696996)) lut_n2564 (.I0(x873), .I1(x874), .I2(x875), .I3(n2554), .I4(n2555), .O(n2564));
  LUT5 #(.INIT(32'hFF969600)) lut_n2565 (.I0(x879), .I1(x880), .I2(x881), .I3(n2563), .I4(n2564), .O(n2565));
  LUT3 #(.INIT(8'h96)) lut_n2566 (.I0(x888), .I1(x889), .I2(x890), .O(n2566));
  LUT5 #(.INIT(32'h96696996)) lut_n2567 (.I0(x879), .I1(x880), .I2(x881), .I3(n2563), .I4(n2564), .O(n2567));
  LUT5 #(.INIT(32'hFF969600)) lut_n2568 (.I0(x885), .I1(x886), .I2(x887), .I3(n2566), .I4(n2567), .O(n2568));
  LUT3 #(.INIT(8'h96)) lut_n2569 (.I0(n2553), .I1(n2556), .I2(n2557), .O(n2569));
  LUT3 #(.INIT(8'hE8)) lut_n2570 (.I0(n2565), .I1(n2568), .I2(n2569), .O(n2570));
  LUT3 #(.INIT(8'h96)) lut_n2571 (.I0(x894), .I1(x895), .I2(x896), .O(n2571));
  LUT5 #(.INIT(32'h96696996)) lut_n2572 (.I0(x885), .I1(x886), .I2(x887), .I3(n2566), .I4(n2567), .O(n2572));
  LUT5 #(.INIT(32'hFF969600)) lut_n2573 (.I0(x891), .I1(x892), .I2(x893), .I3(n2571), .I4(n2572), .O(n2573));
  LUT3 #(.INIT(8'h96)) lut_n2574 (.I0(x900), .I1(x901), .I2(x902), .O(n2574));
  LUT5 #(.INIT(32'h96696996)) lut_n2575 (.I0(x891), .I1(x892), .I2(x893), .I3(n2571), .I4(n2572), .O(n2575));
  LUT5 #(.INIT(32'hFF969600)) lut_n2576 (.I0(x897), .I1(x898), .I2(x899), .I3(n2574), .I4(n2575), .O(n2576));
  LUT3 #(.INIT(8'h96)) lut_n2577 (.I0(n2565), .I1(n2568), .I2(n2569), .O(n2577));
  LUT3 #(.INIT(8'hE8)) lut_n2578 (.I0(n2573), .I1(n2576), .I2(n2577), .O(n2578));
  LUT3 #(.INIT(8'h96)) lut_n2579 (.I0(n2550), .I1(n2558), .I2(n2559), .O(n2579));
  LUT3 #(.INIT(8'h8E)) lut_n2580 (.I0(n2570), .I1(n2578), .I2(n2579), .O(n2580));
  LUT3 #(.INIT(8'h96)) lut_n2581 (.I0(x906), .I1(x907), .I2(x908), .O(n2581));
  LUT5 #(.INIT(32'h96696996)) lut_n2582 (.I0(x897), .I1(x898), .I2(x899), .I3(n2574), .I4(n2575), .O(n2582));
  LUT5 #(.INIT(32'hFF969600)) lut_n2583 (.I0(x903), .I1(x904), .I2(x905), .I3(n2581), .I4(n2582), .O(n2583));
  LUT3 #(.INIT(8'h96)) lut_n2584 (.I0(x912), .I1(x913), .I2(x914), .O(n2584));
  LUT5 #(.INIT(32'h96696996)) lut_n2585 (.I0(x903), .I1(x904), .I2(x905), .I3(n2581), .I4(n2582), .O(n2585));
  LUT5 #(.INIT(32'hFF969600)) lut_n2586 (.I0(x909), .I1(x910), .I2(x911), .I3(n2584), .I4(n2585), .O(n2586));
  LUT3 #(.INIT(8'h96)) lut_n2587 (.I0(n2573), .I1(n2576), .I2(n2577), .O(n2587));
  LUT3 #(.INIT(8'hE8)) lut_n2588 (.I0(n2583), .I1(n2586), .I2(n2587), .O(n2588));
  LUT3 #(.INIT(8'h96)) lut_n2589 (.I0(x918), .I1(x919), .I2(x920), .O(n2589));
  LUT5 #(.INIT(32'h96696996)) lut_n2590 (.I0(x909), .I1(x910), .I2(x911), .I3(n2584), .I4(n2585), .O(n2590));
  LUT5 #(.INIT(32'hFF969600)) lut_n2591 (.I0(x915), .I1(x916), .I2(x917), .I3(n2589), .I4(n2590), .O(n2591));
  LUT3 #(.INIT(8'h96)) lut_n2592 (.I0(x924), .I1(x925), .I2(x926), .O(n2592));
  LUT5 #(.INIT(32'h96696996)) lut_n2593 (.I0(x915), .I1(x916), .I2(x917), .I3(n2589), .I4(n2590), .O(n2593));
  LUT5 #(.INIT(32'hFF969600)) lut_n2594 (.I0(x921), .I1(x922), .I2(x923), .I3(n2592), .I4(n2593), .O(n2594));
  LUT3 #(.INIT(8'h96)) lut_n2595 (.I0(n2583), .I1(n2586), .I2(n2587), .O(n2595));
  LUT3 #(.INIT(8'hE8)) lut_n2596 (.I0(n2591), .I1(n2594), .I2(n2595), .O(n2596));
  LUT3 #(.INIT(8'h96)) lut_n2597 (.I0(n2570), .I1(n2578), .I2(n2579), .O(n2597));
  LUT3 #(.INIT(8'h8E)) lut_n2598 (.I0(n2588), .I1(n2596), .I2(n2597), .O(n2598));
  LUT3 #(.INIT(8'h96)) lut_n2599 (.I0(n2542), .I1(n2560), .I2(n2561), .O(n2599));
  LUT3 #(.INIT(8'hE8)) lut_n2600 (.I0(n2580), .I1(n2598), .I2(n2599), .O(n2600));
  LUT3 #(.INIT(8'h96)) lut_n2601 (.I0(n2483), .I1(n2521), .I2(n2522), .O(n2601));
  LUT3 #(.INIT(8'hE8)) lut_n2602 (.I0(n2562), .I1(n2600), .I2(n2601), .O(n2602));
  LUT3 #(.INIT(8'h96)) lut_n2603 (.I0(x930), .I1(x931), .I2(x932), .O(n2603));
  LUT5 #(.INIT(32'h96696996)) lut_n2604 (.I0(x921), .I1(x922), .I2(x923), .I3(n2592), .I4(n2593), .O(n2604));
  LUT5 #(.INIT(32'hFF969600)) lut_n2605 (.I0(x927), .I1(x928), .I2(x929), .I3(n2603), .I4(n2604), .O(n2605));
  LUT3 #(.INIT(8'h96)) lut_n2606 (.I0(x936), .I1(x937), .I2(x938), .O(n2606));
  LUT5 #(.INIT(32'h96696996)) lut_n2607 (.I0(x927), .I1(x928), .I2(x929), .I3(n2603), .I4(n2604), .O(n2607));
  LUT5 #(.INIT(32'hFF969600)) lut_n2608 (.I0(x933), .I1(x934), .I2(x935), .I3(n2606), .I4(n2607), .O(n2608));
  LUT3 #(.INIT(8'h96)) lut_n2609 (.I0(n2591), .I1(n2594), .I2(n2595), .O(n2609));
  LUT3 #(.INIT(8'hE8)) lut_n2610 (.I0(n2605), .I1(n2608), .I2(n2609), .O(n2610));
  LUT3 #(.INIT(8'h96)) lut_n2611 (.I0(x942), .I1(x943), .I2(x944), .O(n2611));
  LUT5 #(.INIT(32'h96696996)) lut_n2612 (.I0(x933), .I1(x934), .I2(x935), .I3(n2606), .I4(n2607), .O(n2612));
  LUT5 #(.INIT(32'hFF969600)) lut_n2613 (.I0(x939), .I1(x940), .I2(x941), .I3(n2611), .I4(n2612), .O(n2613));
  LUT3 #(.INIT(8'h96)) lut_n2614 (.I0(x948), .I1(x949), .I2(x950), .O(n2614));
  LUT5 #(.INIT(32'h96696996)) lut_n2615 (.I0(x939), .I1(x940), .I2(x941), .I3(n2611), .I4(n2612), .O(n2615));
  LUT5 #(.INIT(32'hFF969600)) lut_n2616 (.I0(x945), .I1(x946), .I2(x947), .I3(n2614), .I4(n2615), .O(n2616));
  LUT3 #(.INIT(8'h96)) lut_n2617 (.I0(n2605), .I1(n2608), .I2(n2609), .O(n2617));
  LUT3 #(.INIT(8'hE8)) lut_n2618 (.I0(n2613), .I1(n2616), .I2(n2617), .O(n2618));
  LUT3 #(.INIT(8'h96)) lut_n2619 (.I0(n2588), .I1(n2596), .I2(n2597), .O(n2619));
  LUT3 #(.INIT(8'h8E)) lut_n2620 (.I0(n2610), .I1(n2618), .I2(n2619), .O(n2620));
  LUT3 #(.INIT(8'h96)) lut_n2621 (.I0(x954), .I1(x955), .I2(x956), .O(n2621));
  LUT5 #(.INIT(32'h96696996)) lut_n2622 (.I0(x945), .I1(x946), .I2(x947), .I3(n2614), .I4(n2615), .O(n2622));
  LUT5 #(.INIT(32'hFF969600)) lut_n2623 (.I0(x951), .I1(x952), .I2(x953), .I3(n2621), .I4(n2622), .O(n2623));
  LUT3 #(.INIT(8'h96)) lut_n2624 (.I0(x960), .I1(x961), .I2(x962), .O(n2624));
  LUT5 #(.INIT(32'h96696996)) lut_n2625 (.I0(x951), .I1(x952), .I2(x953), .I3(n2621), .I4(n2622), .O(n2625));
  LUT5 #(.INIT(32'hFF969600)) lut_n2626 (.I0(x957), .I1(x958), .I2(x959), .I3(n2624), .I4(n2625), .O(n2626));
  LUT3 #(.INIT(8'h96)) lut_n2627 (.I0(n2613), .I1(n2616), .I2(n2617), .O(n2627));
  LUT3 #(.INIT(8'hE8)) lut_n2628 (.I0(n2623), .I1(n2626), .I2(n2627), .O(n2628));
  LUT3 #(.INIT(8'h96)) lut_n2629 (.I0(x966), .I1(x967), .I2(x968), .O(n2629));
  LUT5 #(.INIT(32'h96696996)) lut_n2630 (.I0(x957), .I1(x958), .I2(x959), .I3(n2624), .I4(n2625), .O(n2630));
  LUT5 #(.INIT(32'hFF969600)) lut_n2631 (.I0(x963), .I1(x964), .I2(x965), .I3(n2629), .I4(n2630), .O(n2631));
  LUT3 #(.INIT(8'h96)) lut_n2632 (.I0(x972), .I1(x973), .I2(x974), .O(n2632));
  LUT5 #(.INIT(32'h96696996)) lut_n2633 (.I0(x963), .I1(x964), .I2(x965), .I3(n2629), .I4(n2630), .O(n2633));
  LUT5 #(.INIT(32'hFF969600)) lut_n2634 (.I0(x969), .I1(x970), .I2(x971), .I3(n2632), .I4(n2633), .O(n2634));
  LUT3 #(.INIT(8'h96)) lut_n2635 (.I0(n2623), .I1(n2626), .I2(n2627), .O(n2635));
  LUT3 #(.INIT(8'hE8)) lut_n2636 (.I0(n2631), .I1(n2634), .I2(n2635), .O(n2636));
  LUT3 #(.INIT(8'h96)) lut_n2637 (.I0(n2610), .I1(n2618), .I2(n2619), .O(n2637));
  LUT3 #(.INIT(8'h8E)) lut_n2638 (.I0(n2628), .I1(n2636), .I2(n2637), .O(n2638));
  LUT3 #(.INIT(8'h96)) lut_n2639 (.I0(n2580), .I1(n2598), .I2(n2599), .O(n2639));
  LUT3 #(.INIT(8'h96)) lut_n2640 (.I0(x978), .I1(x979), .I2(x980), .O(n2640));
  LUT5 #(.INIT(32'h96696996)) lut_n2641 (.I0(x969), .I1(x970), .I2(x971), .I3(n2632), .I4(n2633), .O(n2641));
  LUT5 #(.INIT(32'hFF969600)) lut_n2642 (.I0(x975), .I1(x976), .I2(x977), .I3(n2640), .I4(n2641), .O(n2642));
  LUT3 #(.INIT(8'h96)) lut_n2643 (.I0(x984), .I1(x985), .I2(x986), .O(n2643));
  LUT5 #(.INIT(32'h96696996)) lut_n2644 (.I0(x975), .I1(x976), .I2(x977), .I3(n2640), .I4(n2641), .O(n2644));
  LUT5 #(.INIT(32'hFF969600)) lut_n2645 (.I0(x981), .I1(x982), .I2(x983), .I3(n2643), .I4(n2644), .O(n2645));
  LUT3 #(.INIT(8'h96)) lut_n2646 (.I0(n2631), .I1(n2634), .I2(n2635), .O(n2646));
  LUT3 #(.INIT(8'hE8)) lut_n2647 (.I0(n2642), .I1(n2645), .I2(n2646), .O(n2647));
  LUT3 #(.INIT(8'h96)) lut_n2648 (.I0(x990), .I1(x991), .I2(x992), .O(n2648));
  LUT5 #(.INIT(32'h96696996)) lut_n2649 (.I0(x981), .I1(x982), .I2(x983), .I3(n2643), .I4(n2644), .O(n2649));
  LUT5 #(.INIT(32'hFF969600)) lut_n2650 (.I0(x987), .I1(x988), .I2(x989), .I3(n2648), .I4(n2649), .O(n2650));
  LUT3 #(.INIT(8'h96)) lut_n2651 (.I0(x996), .I1(x997), .I2(x998), .O(n2651));
  LUT5 #(.INIT(32'h96696996)) lut_n2652 (.I0(x987), .I1(x988), .I2(x989), .I3(n2648), .I4(n2649), .O(n2652));
  LUT5 #(.INIT(32'hFF969600)) lut_n2653 (.I0(x993), .I1(x994), .I2(x995), .I3(n2651), .I4(n2652), .O(n2653));
  LUT3 #(.INIT(8'h96)) lut_n2654 (.I0(n2642), .I1(n2645), .I2(n2646), .O(n2654));
  LUT3 #(.INIT(8'hE8)) lut_n2655 (.I0(n2650), .I1(n2653), .I2(n2654), .O(n2655));
  LUT3 #(.INIT(8'h96)) lut_n2656 (.I0(n2628), .I1(n2636), .I2(n2637), .O(n2656));
  LUT3 #(.INIT(8'h8E)) lut_n2657 (.I0(n2647), .I1(n2655), .I2(n2656), .O(n2657));
  LUT3 #(.INIT(8'h96)) lut_n2658 (.I0(x1002), .I1(x1003), .I2(x1004), .O(n2658));
  LUT5 #(.INIT(32'h96696996)) lut_n2659 (.I0(x993), .I1(x994), .I2(x995), .I3(n2651), .I4(n2652), .O(n2659));
  LUT5 #(.INIT(32'hFF969600)) lut_n2660 (.I0(x999), .I1(x1000), .I2(x1001), .I3(n2658), .I4(n2659), .O(n2660));
  LUT3 #(.INIT(8'h96)) lut_n2661 (.I0(x1008), .I1(x1009), .I2(x1010), .O(n2661));
  LUT5 #(.INIT(32'h96696996)) lut_n2662 (.I0(x999), .I1(x1000), .I2(x1001), .I3(n2658), .I4(n2659), .O(n2662));
  LUT5 #(.INIT(32'hFF969600)) lut_n2663 (.I0(x1005), .I1(x1006), .I2(x1007), .I3(n2661), .I4(n2662), .O(n2663));
  LUT3 #(.INIT(8'h96)) lut_n2664 (.I0(n2650), .I1(n2653), .I2(n2654), .O(n2664));
  LUT5 #(.INIT(32'h96696996)) lut_n2665 (.I0(x1005), .I1(x1006), .I2(x1007), .I3(n2661), .I4(n2662), .O(n2665));
  LUT5 #(.INIT(32'hFF969600)) lut_n2666 (.I0(x1011), .I1(x1012), .I2(x1013), .I3(x1014), .I4(n2665), .O(n2666));
  LUT3 #(.INIT(8'h96)) lut_n2667 (.I0(n2647), .I1(n2655), .I2(n2656), .O(n2667));
  LUT5 #(.INIT(32'h8000FEE8)) lut_n2668 (.I0(n2660), .I1(n2663), .I2(n2664), .I3(n2666), .I4(n2667), .O(n2668));
  LUT3 #(.INIT(8'h96)) lut_n2669 (.I0(n2562), .I1(n2600), .I2(n2601), .O(n2669));
  LUT6 #(.INIT(64'hFFFEFEE8E8808000)) lut_n2670 (.I0(n2620), .I1(n2638), .I2(n2639), .I3(n2657), .I4(n2668), .I5(n2669), .O(n2670));
  LUT3 #(.INIT(8'h96)) lut_n2671 (.I0(n2207), .I1(n2365), .I2(n2366), .O(n2671));
  LUT6 #(.INIT(64'hFFFEFEE8E8808000)) lut_n2672 (.I0(n2445), .I1(n2523), .I2(n2524), .I3(n2602), .I4(n2670), .I5(n2671), .O(n2672));
  LUT5 #(.INIT(32'hFF969600)) lut_n2673 (.I0(n1788), .I1(n2047), .I2(n2048), .I3(n2367), .I4(n2672), .O(n2673));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n2674 (.I0(n1314), .I1(n1472), .I2(n1630), .I3(n2049), .I4(n2673), .O(n2674));
  assign y0 = n2674;
endmodule
