module top (x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38, y0);
  input x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, x32, x33, x34, x35, x36, x37, x38;
  output y0;
  wire n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88;
  LUT3 #(.INIT(8'hE8)) lut_n41 (.I0(x0), .I1(x1), .I2(x2), .O(n41));
  LUT3 #(.INIT(8'hE8)) lut_n42 (.I0(x6), .I1(x7), .I2(x8), .O(n42));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n43 (.I0(x3), .I1(x4), .I2(x5), .I3(n41), .I4(n42), .O(n43));
  LUT3 #(.INIT(8'hE8)) lut_n44 (.I0(x12), .I1(x13), .I2(x14), .O(n44));
  LUT5 #(.INIT(32'hE81717E8)) lut_n45 (.I0(x3), .I1(x4), .I2(x5), .I3(n41), .I4(n42), .O(n45));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n46 (.I0(x9), .I1(x10), .I2(x11), .I3(n44), .I4(n45), .O(n46));
  LUT3 #(.INIT(8'hE8)) lut_n47 (.I0(x18), .I1(x19), .I2(x20), .O(n47));
  LUT5 #(.INIT(32'hE81717E8)) lut_n48 (.I0(x9), .I1(x10), .I2(x11), .I3(n44), .I4(n45), .O(n48));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n49 (.I0(x15), .I1(x16), .I2(x17), .I3(n47), .I4(n48), .O(n49));
  LUT3 #(.INIT(8'hE8)) lut_n50 (.I0(n43), .I1(n46), .I2(n49), .O(n50));
  LUT3 #(.INIT(8'hE8)) lut_n51 (.I0(x24), .I1(x25), .I2(x26), .O(n51));
  LUT5 #(.INIT(32'hE81717E8)) lut_n52 (.I0(x15), .I1(x16), .I2(x17), .I3(n47), .I4(n48), .O(n52));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n53 (.I0(x21), .I1(x22), .I2(x23), .I3(n51), .I4(n52), .O(n53));
  LUT3 #(.INIT(8'hE8)) lut_n54 (.I0(x27), .I1(x28), .I2(x29), .O(n54));
  LUT5 #(.INIT(32'hE81717E8)) lut_n55 (.I0(x21), .I1(x22), .I2(x23), .I3(n51), .I4(n52), .O(n55));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n56 (.I0(x30), .I1(x31), .I2(x32), .I3(n54), .I4(n55), .O(n56));
  LUT3 #(.INIT(8'h96)) lut_n57 (.I0(n43), .I1(n46), .I2(n49), .O(n57));
  LUT3 #(.INIT(8'hE8)) lut_n58 (.I0(n53), .I1(n56), .I2(n57), .O(n58));
  LUT3 #(.INIT(8'hE8)) lut_n59 (.I0(x36), .I1(x37), .I2(x38), .O(n59));
  LUT5 #(.INIT(32'hE81717E8)) lut_n60 (.I0(x30), .I1(x31), .I2(x32), .I3(n54), .I4(n55), .O(n60));
  LUT5 #(.INIT(32'hFFE8E800)) lut_n61 (.I0(x33), .I1(x34), .I2(x35), .I3(n59), .I4(n60), .O(n61));
  LUT3 #(.INIT(8'h96)) lut_n62 (.I0(x0), .I1(x1), .I2(x2), .O(n62));
  LUT3 #(.INIT(8'h96)) lut_n63 (.I0(x6), .I1(x7), .I2(x8), .O(n63));
  LUT5 #(.INIT(32'hFF969600)) lut_n64 (.I0(x3), .I1(x4), .I2(x5), .I3(n62), .I4(n63), .O(n64));
  LUT3 #(.INIT(8'h96)) lut_n65 (.I0(x12), .I1(x13), .I2(x14), .O(n65));
  LUT5 #(.INIT(32'h96696996)) lut_n66 (.I0(x3), .I1(x4), .I2(x5), .I3(n62), .I4(n63), .O(n66));
  LUT5 #(.INIT(32'hFF969600)) lut_n67 (.I0(x9), .I1(x10), .I2(x11), .I3(n65), .I4(n66), .O(n67));
  LUT5 #(.INIT(32'hE81717E8)) lut_n68 (.I0(x33), .I1(x34), .I2(x35), .I3(n59), .I4(n60), .O(n68));
  LUT3 #(.INIT(8'hE8)) lut_n69 (.I0(n64), .I1(n67), .I2(n68), .O(n69));
  LUT3 #(.INIT(8'h96)) lut_n70 (.I0(n53), .I1(n56), .I2(n57), .O(n70));
  LUT3 #(.INIT(8'hE8)) lut_n71 (.I0(n61), .I1(n69), .I2(n70), .O(n71));
  LUT3 #(.INIT(8'h96)) lut_n72 (.I0(x18), .I1(x19), .I2(x20), .O(n72));
  LUT5 #(.INIT(32'h96696996)) lut_n73 (.I0(x9), .I1(x10), .I2(x11), .I3(n65), .I4(n66), .O(n73));
  LUT5 #(.INIT(32'hFF969600)) lut_n74 (.I0(x15), .I1(x16), .I2(x17), .I3(n72), .I4(n73), .O(n74));
  LUT3 #(.INIT(8'h96)) lut_n75 (.I0(x24), .I1(x25), .I2(x26), .O(n75));
  LUT5 #(.INIT(32'h96696996)) lut_n76 (.I0(x15), .I1(x16), .I2(x17), .I3(n72), .I4(n73), .O(n76));
  LUT5 #(.INIT(32'hFF969600)) lut_n77 (.I0(x21), .I1(x22), .I2(x23), .I3(n75), .I4(n76), .O(n77));
  LUT3 #(.INIT(8'h96)) lut_n78 (.I0(n64), .I1(n67), .I2(n68), .O(n78));
  LUT3 #(.INIT(8'hE8)) lut_n79 (.I0(n74), .I1(n77), .I2(n78), .O(n79));
  LUT3 #(.INIT(8'h96)) lut_n80 (.I0(x30), .I1(x31), .I2(x32), .O(n80));
  LUT3 #(.INIT(8'h96)) lut_n81 (.I0(x27), .I1(x28), .I2(x29), .O(n81));
  LUT5 #(.INIT(32'h96696996)) lut_n82 (.I0(x21), .I1(x22), .I2(x23), .I3(n75), .I4(n76), .O(n82));
  LUT3 #(.INIT(8'h96)) lut_n83 (.I0(x33), .I1(x34), .I2(x35), .O(n83));
  LUT3 #(.INIT(8'h96)) lut_n84 (.I0(x36), .I1(x37), .I2(x38), .O(n84));
  LUT3 #(.INIT(8'h96)) lut_n85 (.I0(n74), .I1(n77), .I2(n78), .O(n85));
  LUT6 #(.INIT(64'hFFFEFEE8E8808000)) lut_n86 (.I0(n80), .I1(n81), .I2(n82), .I3(n83), .I4(n84), .I5(n85), .O(n86));
  LUT3 #(.INIT(8'h96)) lut_n87 (.I0(n61), .I1(n69), .I2(n70), .O(n87));
  LUT6 #(.INIT(64'hFEE8E8E8E8E8E880)) lut_n88 (.I0(n50), .I1(n58), .I2(n71), .I3(n79), .I4(n86), .I5(n87), .O(n88));
  assign y0 = n88;
endmodule
