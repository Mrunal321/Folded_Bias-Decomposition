`timescale 1ns/1ps
`default_nettype none

module tb_top;
  // 511-bit input vector
  reg  [510:0] x = 511'b0;
  wire       y0;
  reg  [63:0] idx;

  // DUT instantiation
  top dut (
    .x0(x[0]), .x1(x[1]), .x2(x[2]), .x3(x[3]), .x4(x[4]), .x5(x[5]), .x6(x[6]), .x7(x[7]), .x8(x[8]), .x9(x[9]), .x10(x[10]), .x11(x[11]), .x12(x[12]), .x13(x[13]), .x14(x[14]), .x15(x[15]), .x16(x[16]), .x17(x[17]), .x18(x[18]), .x19(x[19]), .x20(x[20]), .x21(x[21]), .x22(x[22]), .x23(x[23]), .x24(x[24]), .x25(x[25]), .x26(x[26]), .x27(x[27]), .x28(x[28]), .x29(x[29]), .x30(x[30]), .x31(x[31]), .x32(x[32]), .x33(x[33]), .x34(x[34]), .x35(x[35]), .x36(x[36]), .x37(x[37]), .x38(x[38]), .x39(x[39]), .x40(x[40]), .x41(x[41]), .x42(x[42]), .x43(x[43]), .x44(x[44]), .x45(x[45]), .x46(x[46]), .x47(x[47]), .x48(x[48]), .x49(x[49]), .x50(x[50]), .x51(x[51]), .x52(x[52]), .x53(x[53]), .x54(x[54]), .x55(x[55]), .x56(x[56]), .x57(x[57]), .x58(x[58]), .x59(x[59]), .x60(x[60]), .x61(x[61]), .x62(x[62]), .x63(x[63]), .x64(x[64]), .x65(x[65]), .x66(x[66]), .x67(x[67]), .x68(x[68]), .x69(x[69]), .x70(x[70]), .x71(x[71]), .x72(x[72]), .x73(x[73]), .x74(x[74]), .x75(x[75]), .x76(x[76]), .x77(x[77]), .x78(x[78]), .x79(x[79]), .x80(x[80]), .x81(x[81]), .x82(x[82]), .x83(x[83]), .x84(x[84]), .x85(x[85]), .x86(x[86]), .x87(x[87]), .x88(x[88]), .x89(x[89]), .x90(x[90]), .x91(x[91]), .x92(x[92]), .x93(x[93]), .x94(x[94]), .x95(x[95]), .x96(x[96]), .x97(x[97]), .x98(x[98]), .x99(x[99]), .x100(x[100]), .x101(x[101]), .x102(x[102]), .x103(x[103]), .x104(x[104]), .x105(x[105]), .x106(x[106]), .x107(x[107]), .x108(x[108]), .x109(x[109]), .x110(x[110]), .x111(x[111]), .x112(x[112]), .x113(x[113]), .x114(x[114]), .x115(x[115]), .x116(x[116]), .x117(x[117]), .x118(x[118]), .x119(x[119]), .x120(x[120]), .x121(x[121]), .x122(x[122]), .x123(x[123]), .x124(x[124]), .x125(x[125]), .x126(x[126]), .x127(x[127]), .x128(x[128]), .x129(x[129]), .x130(x[130]), .x131(x[131]), .x132(x[132]), .x133(x[133]), .x134(x[134]), .x135(x[135]), .x136(x[136]), .x137(x[137]), .x138(x[138]), .x139(x[139]), .x140(x[140]), .x141(x[141]), .x142(x[142]), .x143(x[143]), .x144(x[144]), .x145(x[145]), .x146(x[146]), .x147(x[147]), .x148(x[148]), .x149(x[149]), .x150(x[150]), .x151(x[151]), .x152(x[152]), .x153(x[153]), .x154(x[154]), .x155(x[155]), .x156(x[156]), .x157(x[157]), .x158(x[158]), .x159(x[159]), .x160(x[160]), .x161(x[161]), .x162(x[162]), .x163(x[163]), .x164(x[164]), .x165(x[165]), .x166(x[166]), .x167(x[167]), .x168(x[168]), .x169(x[169]), .x170(x[170]), .x171(x[171]), .x172(x[172]), .x173(x[173]), .x174(x[174]), .x175(x[175]), .x176(x[176]), .x177(x[177]), .x178(x[178]), .x179(x[179]), .x180(x[180]), .x181(x[181]), .x182(x[182]), .x183(x[183]), .x184(x[184]), .x185(x[185]), .x186(x[186]), .x187(x[187]), .x188(x[188]), .x189(x[189]), .x190(x[190]), .x191(x[191]), .x192(x[192]), .x193(x[193]), .x194(x[194]), .x195(x[195]), .x196(x[196]), .x197(x[197]), .x198(x[198]), .x199(x[199]), .x200(x[200]), .x201(x[201]), .x202(x[202]), .x203(x[203]), .x204(x[204]), .x205(x[205]), .x206(x[206]), .x207(x[207]), .x208(x[208]), .x209(x[209]), .x210(x[210]), .x211(x[211]), .x212(x[212]), .x213(x[213]), .x214(x[214]), .x215(x[215]), .x216(x[216]), .x217(x[217]), .x218(x[218]), .x219(x[219]), .x220(x[220]), .x221(x[221]), .x222(x[222]), .x223(x[223]), .x224(x[224]), .x225(x[225]), .x226(x[226]), .x227(x[227]), .x228(x[228]), .x229(x[229]), .x230(x[230]), .x231(x[231]), .x232(x[232]), .x233(x[233]), .x234(x[234]), .x235(x[235]), .x236(x[236]), .x237(x[237]), .x238(x[238]), .x239(x[239]), .x240(x[240]), .x241(x[241]), .x242(x[242]), .x243(x[243]), .x244(x[244]), .x245(x[245]), .x246(x[246]), .x247(x[247]), .x248(x[248]), .x249(x[249]), .x250(x[250]), .x251(x[251]), .x252(x[252]), .x253(x[253]), .x254(x[254]), .x255(x[255]), .x256(x[256]), .x257(x[257]), .x258(x[258]), .x259(x[259]), .x260(x[260]), .x261(x[261]), .x262(x[262]), .x263(x[263]), .x264(x[264]), .x265(x[265]), .x266(x[266]), .x267(x[267]), .x268(x[268]), .x269(x[269]), .x270(x[270]), .x271(x[271]), .x272(x[272]), .x273(x[273]), .x274(x[274]), .x275(x[275]), .x276(x[276]), .x277(x[277]), .x278(x[278]), .x279(x[279]), .x280(x[280]), .x281(x[281]), .x282(x[282]), .x283(x[283]), .x284(x[284]), .x285(x[285]), .x286(x[286]), .x287(x[287]), .x288(x[288]), .x289(x[289]), .x290(x[290]), .x291(x[291]), .x292(x[292]), .x293(x[293]), .x294(x[294]), .x295(x[295]), .x296(x[296]), .x297(x[297]), .x298(x[298]), .x299(x[299]), .x300(x[300]), .x301(x[301]), .x302(x[302]), .x303(x[303]), .x304(x[304]), .x305(x[305]), .x306(x[306]), .x307(x[307]), .x308(x[308]), .x309(x[309]), .x310(x[310]), .x311(x[311]), .x312(x[312]), .x313(x[313]), .x314(x[314]), .x315(x[315]), .x316(x[316]), .x317(x[317]), .x318(x[318]), .x319(x[319]), .x320(x[320]), .x321(x[321]), .x322(x[322]), .x323(x[323]), .x324(x[324]), .x325(x[325]), .x326(x[326]), .x327(x[327]), .x328(x[328]), .x329(x[329]), .x330(x[330]), .x331(x[331]), .x332(x[332]), .x333(x[333]), .x334(x[334]), .x335(x[335]), .x336(x[336]), .x337(x[337]), .x338(x[338]), .x339(x[339]), .x340(x[340]), .x341(x[341]), .x342(x[342]), .x343(x[343]), .x344(x[344]), .x345(x[345]), .x346(x[346]), .x347(x[347]), .x348(x[348]), .x349(x[349]), .x350(x[350]), .x351(x[351]), .x352(x[352]), .x353(x[353]), .x354(x[354]), .x355(x[355]), .x356(x[356]), .x357(x[357]), .x358(x[358]), .x359(x[359]), .x360(x[360]), .x361(x[361]), .x362(x[362]), .x363(x[363]), .x364(x[364]), .x365(x[365]), .x366(x[366]), .x367(x[367]), .x368(x[368]), .x369(x[369]), .x370(x[370]), .x371(x[371]), .x372(x[372]), .x373(x[373]), .x374(x[374]), .x375(x[375]), .x376(x[376]), .x377(x[377]), .x378(x[378]), .x379(x[379]), .x380(x[380]), .x381(x[381]), .x382(x[382]), .x383(x[383]), .x384(x[384]), .x385(x[385]), .x386(x[386]), .x387(x[387]), .x388(x[388]), .x389(x[389]), .x390(x[390]), .x391(x[391]), .x392(x[392]), .x393(x[393]), .x394(x[394]), .x395(x[395]), .x396(x[396]), .x397(x[397]), .x398(x[398]), .x399(x[399]), .x400(x[400]), .x401(x[401]), .x402(x[402]), .x403(x[403]), .x404(x[404]), .x405(x[405]), .x406(x[406]), .x407(x[407]), .x408(x[408]), .x409(x[409]), .x410(x[410]), .x411(x[411]), .x412(x[412]), .x413(x[413]), .x414(x[414]), .x415(x[415]), .x416(x[416]), .x417(x[417]), .x418(x[418]), .x419(x[419]), .x420(x[420]), .x421(x[421]), .x422(x[422]), .x423(x[423]), .x424(x[424]), .x425(x[425]), .x426(x[426]), .x427(x[427]), .x428(x[428]), .x429(x[429]), .x430(x[430]), .x431(x[431]), .x432(x[432]), .x433(x[433]), .x434(x[434]), .x435(x[435]), .x436(x[436]), .x437(x[437]), .x438(x[438]), .x439(x[439]), .x440(x[440]), .x441(x[441]), .x442(x[442]), .x443(x[443]), .x444(x[444]), .x445(x[445]), .x446(x[446]), .x447(x[447]), .x448(x[448]), .x449(x[449]), .x450(x[450]), .x451(x[451]), .x452(x[452]), .x453(x[453]), .x454(x[454]), .x455(x[455]), .x456(x[456]), .x457(x[457]), .x458(x[458]), .x459(x[459]), .x460(x[460]), .x461(x[461]), .x462(x[462]), .x463(x[463]), .x464(x[464]), .x465(x[465]), .x466(x[466]), .x467(x[467]), .x468(x[468]), .x469(x[469]), .x470(x[470]), .x471(x[471]), .x472(x[472]), .x473(x[473]), .x474(x[474]), .x475(x[475]), .x476(x[476]), .x477(x[477]), .x478(x[478]), .x479(x[479]), .x480(x[480]), .x481(x[481]), .x482(x[482]), .x483(x[483]), .x484(x[484]), .x485(x[485]), .x486(x[486]), .x487(x[487]), .x488(x[488]), .x489(x[489]), .x490(x[490]), .x491(x[491]), .x492(x[492]), .x493(x[493]), .x494(x[494]), .x495(x[495]), .x496(x[496]), .x497(x[497]), .x498(x[498]), .x499(x[499]), .x500(x[500]), .x501(x[501]), .x502(x[502]), .x503(x[503]), .x504(x[504]), .x505(x[505]), .x506(x[506]), .x507(x[507]), .x508(x[508]), .x509(x[509]), .x510(x[510]),
    .y0(y0)
  );

  // Optional reference function (majority reference for sanity check)
  function [8:0] popcount(input [510:0] v);
    integer i; reg [8:0] c;
    begin
      c = 0;
      for (i = 0; i < 511; i = i + 1)
        c = c + v[i];
      popcount = c;
    end
  endfunction

  // Reference majority: at least 256 ones
  wire y_ref = (popcount(x) >= 256);

  localparam [63:0] TOTAL_VECTORS = 64'd6703903964971298549787012499102923063739682910296196688861780721860882015036773488400937149083451713845015929093243025426876941405973284973216824503042048;

  initial begin
    $display("Time | x510 x509 x508 x507 x506 x505 x504 x503 x502 x501 x500 x499 x498 x497 x496 x495 x494 x493 x492 x491 x490 x489 x488 x487 x486 x485 x484 x483 x482 x481 x480 x479 x478 x477 x476 x475 x474 x473 x472 x471 x470 x469 x468 x467 x466 x465 x464 x463 x462 x461 x460 x459 x458 x457 x456 x455 x454 x453 x452 x451 x450 x449 x448 x447 x446 x445 x444 x443 x442 x441 x440 x439 x438 x437 x436 x435 x434 x433 x432 x431 x430 x429 x428 x427 x426 x425 x424 x423 x422 x421 x420 x419 x418 x417 x416 x415 x414 x413 x412 x411 x410 x409 x408 x407 x406 x405 x404 x403 x402 x401 x400 x399 x398 x397 x396 x395 x394 x393 x392 x391 x390 x389 x388 x387 x386 x385 x384 x383 x382 x381 x380 x379 x378 x377 x376 x375 x374 x373 x372 x371 x370 x369 x368 x367 x366 x365 x364 x363 x362 x361 x360 x359 x358 x357 x356 x355 x354 x353 x352 x351 x350 x349 x348 x347 x346 x345 x344 x343 x342 x341 x340 x339 x338 x337 x336 x335 x334 x333 x332 x331 x330 x329 x328 x327 x326 x325 x324 x323 x322 x321 x320 x319 x318 x317 x316 x315 x314 x313 x312 x311 x310 x309 x308 x307 x306 x305 x304 x303 x302 x301 x300 x299 x298 x297 x296 x295 x294 x293 x292 x291 x290 x289 x288 x287 x286 x285 x284 x283 x282 x281 x280 x279 x278 x277 x276 x275 x274 x273 x272 x271 x270 x269 x268 x267 x266 x265 x264 x263 x262 x261 x260 x259 x258 x257 x256 x255 x254 x253 x252 x251 x250 x249 x248 x247 x246 x245 x244 x243 x242 x241 x240 x239 x238 x237 x236 x235 x234 x233 x232 x231 x230 x229 x228 x227 x226 x225 x224 x223 x222 x221 x220 x219 x218 x217 x216 x215 x214 x213 x212 x211 x210 x209 x208 x207 x206 x205 x204 x203 x202 x201 x200 x199 x198 x197 x196 x195 x194 x193 x192 x191 x190 x189 x188 x187 x186 x185 x184 x183 x182 x181 x180 x179 x178 x177 x176 x175 x174 x173 x172 x171 x170 x169 x168 x167 x166 x165 x164 x163 x162 x161 x160 x159 x158 x157 x156 x155 x154 x153 x152 x151 x150 x149 x148 x147 x146 x145 x144 x143 x142 x141 x140 x139 x138 x137 x136 x135 x134 x133 x132 x131 x130 x129 x128 x127 x126 x125 x124 x123 x122 x121 x120 x119 x118 x117 x116 x115 x114 x113 x112 x111 x110 x109 x108 x107 x106 x105 x104 x103 x102 x101 x100 x99 x98 x97 x96 x95 x94 x93 x92 x91 x90 x89 x88 x87 x86 x85 x84 x83 x82 x81 x80 x79 x78 x77 x76 x75 x74 x73 x72 x71 x70 x69 x68 x67 x66 x65 x64 x63 x62 x61 x60 x59 x58 x57 x56 x55 x54 x53 x52 x51 x50 x49 x48 x47 x46 x45 x44 x43 x42 x41 x40 x39 x38 x37 x36 x35 x34 x33 x32 x31 x30 x29 x28 x27 x26 x25 x24 x23 x22 x21 x20 x19 x18 x17 x16 x15 x14 x13 x12 x11 x10 x9 x8 x7 x6 x5 x4 x3 x2 x1 x0 | y0 (DUT) y_ref (Maj511)");
    $display("-----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------");
    // Loop through all 6703903964971298549787012499102923063739682910296196688861780721860882015036773488400937149083451713845015929093243025426876941405973284973216824503042048 combinations
    for (idx = 0; idx < TOTAL_VECTORS; idx = idx + 1) begin
      x = idx[510:0];
      #10 $display("%4t |  %b  |   %b       %b",
                   $time, x, y0, y_ref);
    end
    #10 $finish;
  end

  // Optional mismatch check
  always #1 if (^x !== 1'bx && y0 !== y_ref)
    $display("Mismatch at t=%0t x=%b HW=%0d y0=%0b ref=%0b",
             $time, x, popcount(x), y0, y_ref);

endmodule

`default_nettype wire
